VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.970 524.520 2008.290 524.580 ;
        RECT 2777.090 524.520 2777.410 524.580 ;
        RECT 2007.970 524.380 2777.410 524.520 ;
        RECT 2007.970 524.320 2008.290 524.380 ;
        RECT 2777.090 524.320 2777.410 524.380 ;
        RECT 2777.090 89.660 2777.410 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2777.090 89.520 2899.310 89.660 ;
        RECT 2777.090 89.460 2777.410 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2008.000 524.320 2008.260 524.580 ;
        RECT 2777.120 524.320 2777.380 524.580 ;
        RECT 2777.120 89.460 2777.380 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2007.990 527.835 2008.270 528.205 ;
        RECT 2008.060 524.610 2008.200 527.835 ;
        RECT 2008.000 524.290 2008.260 524.610 ;
        RECT 2777.120 524.290 2777.380 524.610 ;
        RECT 2777.180 89.750 2777.320 524.290 ;
        RECT 2777.120 89.430 2777.380 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2007.990 527.880 2008.270 528.160 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 1997.465 528.170 2001.465 528.320 ;
        RECT 2007.965 528.170 2008.295 528.185 ;
        RECT 1997.465 527.870 2008.295 528.170 ;
        RECT 1997.465 527.720 2001.465 527.870 ;
        RECT 2007.965 527.855 2008.295 527.870 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2770.190 2429.200 2770.510 2429.260 ;
        RECT 2899.450 2429.200 2899.770 2429.260 ;
        RECT 2770.190 2429.060 2899.770 2429.200 ;
        RECT 2770.190 2429.000 2770.510 2429.060 ;
        RECT 2899.450 2429.000 2899.770 2429.060 ;
        RECT 2007.970 1600.620 2008.290 1600.680 ;
        RECT 2770.190 1600.620 2770.510 1600.680 ;
        RECT 2007.970 1600.480 2770.510 1600.620 ;
        RECT 2007.970 1600.420 2008.290 1600.480 ;
        RECT 2770.190 1600.420 2770.510 1600.480 ;
      LAYER via ;
        RECT 2770.220 2429.000 2770.480 2429.260 ;
        RECT 2899.480 2429.000 2899.740 2429.260 ;
        RECT 2008.000 1600.420 2008.260 1600.680 ;
        RECT 2770.220 1600.420 2770.480 1600.680 ;
      LAYER met2 ;
        RECT 2899.470 2433.875 2899.750 2434.245 ;
        RECT 2899.540 2429.290 2899.680 2433.875 ;
        RECT 2770.220 2428.970 2770.480 2429.290 ;
        RECT 2899.480 2428.970 2899.740 2429.290 ;
        RECT 2770.280 1600.710 2770.420 2428.970 ;
        RECT 2008.000 1600.390 2008.260 1600.710 ;
        RECT 2770.220 1600.390 2770.480 1600.710 ;
        RECT 2008.060 1595.805 2008.200 1600.390 ;
        RECT 2007.990 1595.435 2008.270 1595.805 ;
      LAYER via2 ;
        RECT 2899.470 2433.920 2899.750 2434.200 ;
        RECT 2007.990 1595.480 2008.270 1595.760 ;
      LAYER met3 ;
        RECT 2899.445 2434.210 2899.775 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2899.445 2433.910 2924.800 2434.210 ;
        RECT 2899.445 2433.895 2899.775 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 1997.465 1595.770 2001.465 1595.920 ;
        RECT 2007.965 1595.770 2008.295 1595.785 ;
        RECT 1997.465 1595.470 2008.295 1595.770 ;
        RECT 1997.465 1595.320 2001.465 1595.470 ;
        RECT 2007.965 1595.455 2008.295 1595.470 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.970 1704.320 2008.290 1704.380 ;
        RECT 2894.390 1704.320 2894.710 1704.380 ;
        RECT 2007.970 1704.180 2894.710 1704.320 ;
        RECT 2007.970 1704.120 2008.290 1704.180 ;
        RECT 2894.390 1704.120 2894.710 1704.180 ;
      LAYER via ;
        RECT 2008.000 1704.120 2008.260 1704.380 ;
        RECT 2894.420 1704.120 2894.680 1704.380 ;
      LAYER met2 ;
        RECT 2894.410 2669.155 2894.690 2669.525 ;
        RECT 2894.480 1704.410 2894.620 2669.155 ;
        RECT 2008.000 1704.090 2008.260 1704.410 ;
        RECT 2894.420 1704.090 2894.680 1704.410 ;
        RECT 2008.060 1702.565 2008.200 1704.090 ;
        RECT 2007.990 1702.195 2008.270 1702.565 ;
      LAYER via2 ;
        RECT 2894.410 2669.200 2894.690 2669.480 ;
        RECT 2007.990 1702.240 2008.270 1702.520 ;
      LAYER met3 ;
        RECT 2894.385 2669.490 2894.715 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2894.385 2669.190 2924.800 2669.490 ;
        RECT 2894.385 2669.175 2894.715 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 1997.465 1702.530 2001.465 1702.680 ;
        RECT 2007.965 1702.530 2008.295 1702.545 ;
        RECT 1997.465 1702.230 2008.295 1702.530 ;
        RECT 1997.465 1702.080 2001.465 1702.230 ;
        RECT 2007.965 1702.215 2008.295 1702.230 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2777.090 2898.400 2777.410 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2777.090 2898.260 2901.150 2898.400 ;
        RECT 2777.090 2898.200 2777.410 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2007.970 1814.480 2008.290 1814.540 ;
        RECT 2777.090 1814.480 2777.410 1814.540 ;
        RECT 2007.970 1814.340 2777.410 1814.480 ;
        RECT 2007.970 1814.280 2008.290 1814.340 ;
        RECT 2777.090 1814.280 2777.410 1814.340 ;
      LAYER via ;
        RECT 2777.120 2898.200 2777.380 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2008.000 1814.280 2008.260 1814.540 ;
        RECT 2777.120 1814.280 2777.380 1814.540 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2777.120 2898.170 2777.380 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2777.180 1814.570 2777.320 2898.170 ;
        RECT 2008.000 1814.250 2008.260 1814.570 ;
        RECT 2777.120 1814.250 2777.380 1814.570 ;
        RECT 2008.060 1809.325 2008.200 1814.250 ;
        RECT 2007.990 1808.955 2008.270 1809.325 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2007.990 1809.000 2008.270 1809.280 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 1997.465 1809.290 2001.465 1809.440 ;
        RECT 2007.965 1809.290 2008.295 1809.305 ;
        RECT 1997.465 1808.990 2008.295 1809.290 ;
        RECT 1997.465 1808.840 2001.465 1808.990 ;
        RECT 2007.965 1808.975 2008.295 1808.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2783.990 3133.000 2784.310 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2783.990 3132.860 2901.150 3133.000 ;
        RECT 2783.990 3132.800 2784.310 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2007.970 1918.180 2008.290 1918.240 ;
        RECT 2783.990 1918.180 2784.310 1918.240 ;
        RECT 2007.970 1918.040 2784.310 1918.180 ;
        RECT 2007.970 1917.980 2008.290 1918.040 ;
        RECT 2783.990 1917.980 2784.310 1918.040 ;
      LAYER via ;
        RECT 2784.020 3132.800 2784.280 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2008.000 1917.980 2008.260 1918.240 ;
        RECT 2784.020 1917.980 2784.280 1918.240 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2784.020 3132.770 2784.280 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2784.080 1918.270 2784.220 3132.770 ;
        RECT 2008.000 1917.950 2008.260 1918.270 ;
        RECT 2784.020 1917.950 2784.280 1918.270 ;
        RECT 2008.060 1916.085 2008.200 1917.950 ;
        RECT 2007.990 1915.715 2008.270 1916.085 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2007.990 1915.760 2008.270 1916.040 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 1997.465 1916.050 2001.465 1916.200 ;
        RECT 2007.965 1916.050 2008.295 1916.065 ;
        RECT 1997.465 1915.750 2008.295 1916.050 ;
        RECT 1997.465 1915.600 2001.465 1915.750 ;
        RECT 2007.965 1915.735 2008.295 1915.750 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2790.890 3367.600 2791.210 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2790.890 3367.460 2901.150 3367.600 ;
        RECT 2790.890 3367.400 2791.210 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2007.970 2028.340 2008.290 2028.400 ;
        RECT 2790.890 2028.340 2791.210 2028.400 ;
        RECT 2007.970 2028.200 2791.210 2028.340 ;
        RECT 2007.970 2028.140 2008.290 2028.200 ;
        RECT 2790.890 2028.140 2791.210 2028.200 ;
      LAYER via ;
        RECT 2790.920 3367.400 2791.180 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2008.000 2028.140 2008.260 2028.400 ;
        RECT 2790.920 2028.140 2791.180 2028.400 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2790.920 3367.370 2791.180 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2790.980 2028.430 2791.120 3367.370 ;
        RECT 2008.000 2028.110 2008.260 2028.430 ;
        RECT 2790.920 2028.110 2791.180 2028.430 ;
        RECT 2008.060 2022.845 2008.200 2028.110 ;
        RECT 2007.990 2022.475 2008.270 2022.845 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2007.990 2022.520 2008.270 2022.800 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 1997.465 2022.810 2001.465 2022.960 ;
        RECT 2007.965 2022.810 2008.295 2022.825 ;
        RECT 1997.465 2022.510 2008.295 2022.810 ;
        RECT 1997.465 2022.360 2001.465 2022.510 ;
        RECT 2007.965 2022.495 2008.295 2022.510 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3415.555 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
        RECT 2795.105 2753.065 2795.275 2801.175 ;
        RECT 2795.565 2428.705 2795.735 2463.215 ;
        RECT 2795.565 2331.805 2795.735 2366.655 ;
        RECT 2795.565 2138.685 2795.735 2173.535 ;
      LAYER mcon ;
        RECT 2796.485 3415.385 2796.655 3415.555 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
        RECT 2795.105 2801.005 2795.275 2801.175 ;
        RECT 2795.565 2463.045 2795.735 2463.215 ;
        RECT 2795.565 2366.485 2795.735 2366.655 ;
        RECT 2795.565 2173.365 2795.735 2173.535 ;
      LAYER met1 ;
        RECT 2794.570 3422.340 2794.890 3422.400 ;
        RECT 2798.250 3422.340 2798.570 3422.400 ;
        RECT 2794.570 3422.200 2798.570 3422.340 ;
        RECT 2794.570 3422.140 2794.890 3422.200 ;
        RECT 2798.250 3422.140 2798.570 3422.200 ;
        RECT 2794.570 3415.540 2794.890 3415.600 ;
        RECT 2796.425 3415.540 2796.715 3415.585 ;
        RECT 2794.570 3415.400 2796.715 3415.540 ;
        RECT 2794.570 3415.340 2794.890 3415.400 ;
        RECT 2796.425 3415.355 2796.715 3415.400 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2795.030 2801.160 2795.350 2801.220 ;
        RECT 2794.835 2801.020 2795.350 2801.160 ;
        RECT 2795.030 2800.960 2795.350 2801.020 ;
        RECT 2795.045 2753.220 2795.335 2753.265 ;
        RECT 2795.950 2753.220 2796.270 2753.280 ;
        RECT 2795.045 2753.080 2796.270 2753.220 ;
        RECT 2795.045 2753.035 2795.335 2753.080 ;
        RECT 2795.950 2753.020 2796.270 2753.080 ;
        RECT 2795.030 2718.200 2795.350 2718.260 ;
        RECT 2795.950 2718.200 2796.270 2718.260 ;
        RECT 2795.030 2718.060 2796.270 2718.200 ;
        RECT 2795.030 2718.000 2795.350 2718.060 ;
        RECT 2795.950 2718.000 2796.270 2718.060 ;
        RECT 2795.030 2670.260 2795.350 2670.320 ;
        RECT 2795.950 2670.260 2796.270 2670.320 ;
        RECT 2795.030 2670.120 2796.270 2670.260 ;
        RECT 2795.030 2670.060 2795.350 2670.120 ;
        RECT 2795.950 2670.060 2796.270 2670.120 ;
        RECT 2795.950 2622.120 2796.270 2622.380 ;
        RECT 2796.040 2621.980 2796.180 2622.120 ;
        RECT 2796.410 2621.980 2796.730 2622.040 ;
        RECT 2796.040 2621.840 2796.730 2621.980 ;
        RECT 2796.410 2621.780 2796.730 2621.840 ;
        RECT 2795.490 2560.100 2795.810 2560.160 ;
        RECT 2796.870 2560.100 2797.190 2560.160 ;
        RECT 2795.490 2559.960 2797.190 2560.100 ;
        RECT 2795.490 2559.900 2795.810 2559.960 ;
        RECT 2796.870 2559.900 2797.190 2559.960 ;
        RECT 2795.950 2511.820 2796.270 2511.880 ;
        RECT 2796.870 2511.820 2797.190 2511.880 ;
        RECT 2795.950 2511.680 2797.190 2511.820 ;
        RECT 2795.950 2511.620 2796.270 2511.680 ;
        RECT 2796.870 2511.620 2797.190 2511.680 ;
        RECT 2795.490 2463.200 2795.810 2463.260 ;
        RECT 2795.295 2463.060 2795.810 2463.200 ;
        RECT 2795.490 2463.000 2795.810 2463.060 ;
        RECT 2795.490 2428.860 2795.810 2428.920 ;
        RECT 2795.295 2428.720 2795.810 2428.860 ;
        RECT 2795.490 2428.660 2795.810 2428.720 ;
        RECT 2795.030 2380.580 2795.350 2380.640 ;
        RECT 2795.950 2380.580 2796.270 2380.640 ;
        RECT 2795.030 2380.440 2796.270 2380.580 ;
        RECT 2795.030 2380.380 2795.350 2380.440 ;
        RECT 2795.950 2380.380 2796.270 2380.440 ;
        RECT 2795.490 2366.640 2795.810 2366.700 ;
        RECT 2795.295 2366.500 2795.810 2366.640 ;
        RECT 2795.490 2366.440 2795.810 2366.500 ;
        RECT 2795.490 2331.960 2795.810 2332.020 ;
        RECT 2795.295 2331.820 2795.810 2331.960 ;
        RECT 2795.490 2331.760 2795.810 2331.820 ;
        RECT 2794.570 2235.540 2794.890 2235.800 ;
        RECT 2794.660 2235.400 2794.800 2235.540 ;
        RECT 2795.030 2235.400 2795.350 2235.460 ;
        RECT 2794.660 2235.260 2795.350 2235.400 ;
        RECT 2795.030 2235.200 2795.350 2235.260 ;
        RECT 2795.490 2173.520 2795.810 2173.580 ;
        RECT 2795.295 2173.380 2795.810 2173.520 ;
        RECT 2795.490 2173.320 2795.810 2173.380 ;
        RECT 2795.490 2138.840 2795.810 2138.900 ;
        RECT 2795.295 2138.700 2795.810 2138.840 ;
        RECT 2795.490 2138.640 2795.810 2138.700 ;
        RECT 1971.630 2121.840 1971.950 2121.900 ;
        RECT 2795.950 2121.840 2796.270 2121.900 ;
        RECT 1971.630 2121.700 2796.270 2121.840 ;
        RECT 1971.630 2121.640 1971.950 2121.700 ;
        RECT 2795.950 2121.640 2796.270 2121.700 ;
      LAYER via ;
        RECT 2794.600 3422.140 2794.860 3422.400 ;
        RECT 2798.280 3422.140 2798.540 3422.400 ;
        RECT 2794.600 3415.340 2794.860 3415.600 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2795.060 2800.960 2795.320 2801.220 ;
        RECT 2795.980 2753.020 2796.240 2753.280 ;
        RECT 2795.060 2718.000 2795.320 2718.260 ;
        RECT 2795.980 2718.000 2796.240 2718.260 ;
        RECT 2795.060 2670.060 2795.320 2670.320 ;
        RECT 2795.980 2670.060 2796.240 2670.320 ;
        RECT 2795.980 2622.120 2796.240 2622.380 ;
        RECT 2796.440 2621.780 2796.700 2622.040 ;
        RECT 2795.520 2559.900 2795.780 2560.160 ;
        RECT 2796.900 2559.900 2797.160 2560.160 ;
        RECT 2795.980 2511.620 2796.240 2511.880 ;
        RECT 2796.900 2511.620 2797.160 2511.880 ;
        RECT 2795.520 2463.000 2795.780 2463.260 ;
        RECT 2795.520 2428.660 2795.780 2428.920 ;
        RECT 2795.060 2380.380 2795.320 2380.640 ;
        RECT 2795.980 2380.380 2796.240 2380.640 ;
        RECT 2795.520 2366.440 2795.780 2366.700 ;
        RECT 2795.520 2331.760 2795.780 2332.020 ;
        RECT 2794.600 2235.540 2794.860 2235.800 ;
        RECT 2795.060 2235.200 2795.320 2235.460 ;
        RECT 2795.520 2173.320 2795.780 2173.580 ;
        RECT 2795.520 2138.640 2795.780 2138.900 ;
        RECT 1971.660 2121.640 1971.920 2121.900 ;
        RECT 2795.980 2121.640 2796.240 2121.900 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.430 2798.480 3517.600 ;
        RECT 2794.600 3422.110 2794.860 3422.430 ;
        RECT 2798.280 3422.110 2798.540 3422.430 ;
        RECT 2794.660 3415.630 2794.800 3422.110 ;
        RECT 2794.600 3415.310 2794.860 3415.630 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.250 2795.260 2814.870 ;
        RECT 2795.060 2800.930 2795.320 2801.250 ;
        RECT 2795.980 2752.990 2796.240 2753.310 ;
        RECT 2796.040 2718.290 2796.180 2752.990 ;
        RECT 2795.060 2717.970 2795.320 2718.290 ;
        RECT 2795.980 2717.970 2796.240 2718.290 ;
        RECT 2795.120 2670.350 2795.260 2717.970 ;
        RECT 2795.060 2670.030 2795.320 2670.350 ;
        RECT 2795.980 2670.030 2796.240 2670.350 ;
        RECT 2796.040 2622.410 2796.180 2670.030 ;
        RECT 2795.980 2622.090 2796.240 2622.410 ;
        RECT 2796.440 2621.750 2796.700 2622.070 ;
        RECT 2796.500 2608.325 2796.640 2621.750 ;
        RECT 2795.510 2607.955 2795.790 2608.325 ;
        RECT 2796.430 2607.955 2796.710 2608.325 ;
        RECT 2795.580 2560.190 2795.720 2607.955 ;
        RECT 2795.520 2559.870 2795.780 2560.190 ;
        RECT 2796.900 2559.870 2797.160 2560.190 ;
        RECT 2796.960 2511.910 2797.100 2559.870 ;
        RECT 2795.980 2511.765 2796.240 2511.910 ;
        RECT 2794.590 2511.395 2794.870 2511.765 ;
        RECT 2795.970 2511.395 2796.250 2511.765 ;
        RECT 2796.900 2511.590 2797.160 2511.910 ;
        RECT 2794.660 2463.485 2794.800 2511.395 ;
        RECT 2794.590 2463.115 2794.870 2463.485 ;
        RECT 2795.510 2463.115 2795.790 2463.485 ;
        RECT 2795.520 2462.970 2795.780 2463.115 ;
        RECT 2795.520 2428.630 2795.780 2428.950 ;
        RECT 2795.580 2415.090 2795.720 2428.630 ;
        RECT 2795.580 2414.950 2796.180 2415.090 ;
        RECT 2796.040 2380.670 2796.180 2414.950 ;
        RECT 2795.060 2380.410 2795.320 2380.670 ;
        RECT 2795.060 2380.350 2795.720 2380.410 ;
        RECT 2795.980 2380.350 2796.240 2380.670 ;
        RECT 2795.120 2380.270 2795.720 2380.350 ;
        RECT 2795.580 2366.730 2795.720 2380.270 ;
        RECT 2795.520 2366.410 2795.780 2366.730 ;
        RECT 2795.520 2331.730 2795.780 2332.050 ;
        RECT 2795.580 2318.530 2795.720 2331.730 ;
        RECT 2795.580 2318.390 2796.180 2318.530 ;
        RECT 2796.040 2270.365 2796.180 2318.390 ;
        RECT 2794.590 2269.995 2794.870 2270.365 ;
        RECT 2795.970 2269.995 2796.250 2270.365 ;
        RECT 2794.660 2235.830 2794.800 2269.995 ;
        RECT 2794.600 2235.510 2794.860 2235.830 ;
        RECT 2795.060 2235.170 2795.320 2235.490 ;
        RECT 2795.120 2187.290 2795.260 2235.170 ;
        RECT 2795.120 2187.150 2795.720 2187.290 ;
        RECT 2795.580 2173.610 2795.720 2187.150 ;
        RECT 2795.520 2173.290 2795.780 2173.610 ;
        RECT 2795.520 2138.610 2795.780 2138.930 ;
        RECT 2795.580 2125.410 2795.720 2138.610 ;
        RECT 2795.580 2125.270 2796.180 2125.410 ;
        RECT 2796.040 2121.930 2796.180 2125.270 ;
        RECT 1971.660 2121.610 1971.920 2121.930 ;
        RECT 2795.980 2121.610 2796.240 2121.930 ;
        RECT 1971.720 2112.185 1971.860 2121.610 ;
        RECT 1971.720 2111.740 1972.070 2112.185 ;
        RECT 1971.790 2108.185 1972.070 2111.740 ;
      LAYER via2 ;
        RECT 2795.510 2608.000 2795.790 2608.280 ;
        RECT 2796.430 2608.000 2796.710 2608.280 ;
        RECT 2794.590 2511.440 2794.870 2511.720 ;
        RECT 2795.970 2511.440 2796.250 2511.720 ;
        RECT 2794.590 2463.160 2794.870 2463.440 ;
        RECT 2795.510 2463.160 2795.790 2463.440 ;
        RECT 2794.590 2270.040 2794.870 2270.320 ;
        RECT 2795.970 2270.040 2796.250 2270.320 ;
      LAYER met3 ;
        RECT 2795.485 2608.290 2795.815 2608.305 ;
        RECT 2796.405 2608.290 2796.735 2608.305 ;
        RECT 2795.485 2607.990 2796.735 2608.290 ;
        RECT 2795.485 2607.975 2795.815 2607.990 ;
        RECT 2796.405 2607.975 2796.735 2607.990 ;
        RECT 2794.565 2511.730 2794.895 2511.745 ;
        RECT 2795.945 2511.730 2796.275 2511.745 ;
        RECT 2794.565 2511.430 2796.275 2511.730 ;
        RECT 2794.565 2511.415 2794.895 2511.430 ;
        RECT 2795.945 2511.415 2796.275 2511.430 ;
        RECT 2794.565 2463.450 2794.895 2463.465 ;
        RECT 2795.485 2463.450 2795.815 2463.465 ;
        RECT 2794.565 2463.150 2795.815 2463.450 ;
        RECT 2794.565 2463.135 2794.895 2463.150 ;
        RECT 2795.485 2463.135 2795.815 2463.150 ;
        RECT 2794.565 2270.330 2794.895 2270.345 ;
        RECT 2795.945 2270.330 2796.275 2270.345 ;
        RECT 2794.565 2270.030 2796.275 2270.330 ;
        RECT 2794.565 2270.015 2794.895 2270.030 ;
        RECT 2795.945 2270.015 2796.275 2270.030 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 2898.245 2470.515 2946.355 ;
        RECT 2470.805 2815.285 2470.975 2849.455 ;
      LAYER mcon ;
        RECT 2470.345 2946.185 2470.515 2946.355 ;
        RECT 2470.805 2849.285 2470.975 2849.455 ;
      LAYER met1 ;
        RECT 2470.270 3464.160 2470.590 3464.220 ;
        RECT 2474.410 3464.160 2474.730 3464.220 ;
        RECT 2470.270 3464.020 2474.730 3464.160 ;
        RECT 2470.270 3463.960 2470.590 3464.020 ;
        RECT 2474.410 3463.960 2474.730 3464.020 ;
        RECT 2470.270 3367.600 2470.590 3367.660 ;
        RECT 2471.190 3367.600 2471.510 3367.660 ;
        RECT 2470.270 3367.460 2471.510 3367.600 ;
        RECT 2470.270 3367.400 2470.590 3367.460 ;
        RECT 2471.190 3367.400 2471.510 3367.460 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2470.285 2946.340 2470.575 2946.385 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2470.285 2946.200 2471.050 2946.340 ;
        RECT 2470.285 2946.155 2470.575 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2470.270 2898.400 2470.590 2898.460 ;
        RECT 2470.075 2898.260 2470.590 2898.400 ;
        RECT 2470.270 2898.200 2470.590 2898.260 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2470.535 2849.300 2471.050 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2470.745 2815.440 2471.035 2815.485 ;
        RECT 2471.650 2815.440 2471.970 2815.500 ;
        RECT 2470.745 2815.300 2471.970 2815.440 ;
        RECT 2470.745 2815.255 2471.035 2815.300 ;
        RECT 2471.650 2815.240 2471.970 2815.300 ;
        RECT 2470.730 2753.220 2471.050 2753.280 ;
        RECT 2472.110 2753.220 2472.430 2753.280 ;
        RECT 2470.730 2753.080 2472.430 2753.220 ;
        RECT 2470.730 2753.020 2471.050 2753.080 ;
        RECT 2472.110 2753.020 2472.430 2753.080 ;
        RECT 2472.110 2719.220 2472.430 2719.280 ;
        RECT 2471.740 2719.080 2472.430 2719.220 ;
        RECT 2471.740 2718.600 2471.880 2719.080 ;
        RECT 2472.110 2719.020 2472.430 2719.080 ;
        RECT 2471.650 2718.340 2471.970 2718.600 ;
        RECT 2470.730 2656.660 2471.050 2656.720 ;
        RECT 2472.110 2656.660 2472.430 2656.720 ;
        RECT 2470.730 2656.520 2472.430 2656.660 ;
        RECT 2470.730 2656.460 2471.050 2656.520 ;
        RECT 2472.110 2656.460 2472.430 2656.520 ;
        RECT 2472.110 2622.660 2472.430 2622.720 ;
        RECT 2471.740 2622.520 2472.430 2622.660 ;
        RECT 2471.740 2622.040 2471.880 2622.520 ;
        RECT 2472.110 2622.460 2472.430 2622.520 ;
        RECT 2471.650 2621.780 2471.970 2622.040 ;
        RECT 2470.730 2560.100 2471.050 2560.160 ;
        RECT 2472.110 2560.100 2472.430 2560.160 ;
        RECT 2470.730 2559.960 2472.430 2560.100 ;
        RECT 2470.730 2559.900 2471.050 2559.960 ;
        RECT 2472.110 2559.900 2472.430 2559.960 ;
        RECT 2471.190 2511.820 2471.510 2511.880 ;
        RECT 2472.110 2511.820 2472.430 2511.880 ;
        RECT 2471.190 2511.680 2472.430 2511.820 ;
        RECT 2471.190 2511.620 2471.510 2511.680 ;
        RECT 2472.110 2511.620 2472.430 2511.680 ;
        RECT 2470.270 2401.320 2470.590 2401.380 ;
        RECT 2471.190 2401.320 2471.510 2401.380 ;
        RECT 2470.270 2401.180 2471.510 2401.320 ;
        RECT 2470.270 2401.120 2470.590 2401.180 ;
        RECT 2471.190 2401.120 2471.510 2401.180 ;
        RECT 2470.270 2304.760 2470.590 2304.820 ;
        RECT 2471.190 2304.760 2471.510 2304.820 ;
        RECT 2470.270 2304.620 2471.510 2304.760 ;
        RECT 2470.270 2304.560 2470.590 2304.620 ;
        RECT 2471.190 2304.560 2471.510 2304.620 ;
        RECT 2470.270 2208.200 2470.590 2208.260 ;
        RECT 2471.190 2208.200 2471.510 2208.260 ;
        RECT 2470.270 2208.060 2471.510 2208.200 ;
        RECT 2470.270 2208.000 2470.590 2208.060 ;
        RECT 2471.190 2208.000 2471.510 2208.060 ;
        RECT 1794.990 2122.860 1795.310 2122.920 ;
        RECT 2471.190 2122.860 2471.510 2122.920 ;
        RECT 1794.990 2122.720 2471.510 2122.860 ;
        RECT 1794.990 2122.660 1795.310 2122.720 ;
        RECT 2471.190 2122.660 2471.510 2122.720 ;
      LAYER via ;
        RECT 2470.300 3463.960 2470.560 3464.220 ;
        RECT 2474.440 3463.960 2474.700 3464.220 ;
        RECT 2470.300 3367.400 2470.560 3367.660 ;
        RECT 2471.220 3367.400 2471.480 3367.660 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2470.300 2898.200 2470.560 2898.460 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 2470.760 2753.020 2471.020 2753.280 ;
        RECT 2472.140 2753.020 2472.400 2753.280 ;
        RECT 2472.140 2719.020 2472.400 2719.280 ;
        RECT 2471.680 2718.340 2471.940 2718.600 ;
        RECT 2470.760 2656.460 2471.020 2656.720 ;
        RECT 2472.140 2656.460 2472.400 2656.720 ;
        RECT 2472.140 2622.460 2472.400 2622.720 ;
        RECT 2471.680 2621.780 2471.940 2622.040 ;
        RECT 2470.760 2559.900 2471.020 2560.160 ;
        RECT 2472.140 2559.900 2472.400 2560.160 ;
        RECT 2471.220 2511.620 2471.480 2511.880 ;
        RECT 2472.140 2511.620 2472.400 2511.880 ;
        RECT 2470.300 2401.120 2470.560 2401.380 ;
        RECT 2471.220 2401.120 2471.480 2401.380 ;
        RECT 2470.300 2304.560 2470.560 2304.820 ;
        RECT 2471.220 2304.560 2471.480 2304.820 ;
        RECT 2470.300 2208.000 2470.560 2208.260 ;
        RECT 2471.220 2208.000 2471.480 2208.260 ;
        RECT 1795.020 2122.660 1795.280 2122.920 ;
        RECT 2471.220 2122.660 2471.480 2122.920 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3464.250 2474.640 3517.230 ;
        RECT 2470.300 3463.930 2470.560 3464.250 ;
        RECT 2474.440 3463.930 2474.700 3464.250 ;
        RECT 2470.360 3415.370 2470.500 3463.930 ;
        RECT 2470.360 3415.230 2471.420 3415.370 ;
        RECT 2471.280 3367.690 2471.420 3415.230 ;
        RECT 2470.300 3367.370 2470.560 3367.690 ;
        RECT 2471.220 3367.370 2471.480 3367.690 ;
        RECT 2470.360 3318.810 2470.500 3367.370 ;
        RECT 2470.360 3318.670 2471.420 3318.810 ;
        RECT 2471.280 3270.790 2471.420 3318.670 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2470.300 2898.170 2470.560 2898.490 ;
        RECT 2470.360 2863.210 2470.500 2898.170 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.445 2471.880 2815.210 ;
        RECT 2470.750 2801.075 2471.030 2801.445 ;
        RECT 2471.670 2801.075 2471.950 2801.445 ;
        RECT 2470.820 2753.310 2470.960 2801.075 ;
        RECT 2470.760 2752.990 2471.020 2753.310 ;
        RECT 2472.140 2752.990 2472.400 2753.310 ;
        RECT 2472.200 2719.310 2472.340 2752.990 ;
        RECT 2472.140 2718.990 2472.400 2719.310 ;
        RECT 2471.680 2718.310 2471.940 2718.630 ;
        RECT 2471.740 2704.885 2471.880 2718.310 ;
        RECT 2470.750 2704.515 2471.030 2704.885 ;
        RECT 2471.670 2704.515 2471.950 2704.885 ;
        RECT 2470.820 2656.750 2470.960 2704.515 ;
        RECT 2470.760 2656.430 2471.020 2656.750 ;
        RECT 2472.140 2656.430 2472.400 2656.750 ;
        RECT 2472.200 2622.750 2472.340 2656.430 ;
        RECT 2472.140 2622.430 2472.400 2622.750 ;
        RECT 2471.680 2621.750 2471.940 2622.070 ;
        RECT 2471.740 2608.325 2471.880 2621.750 ;
        RECT 2470.750 2607.955 2471.030 2608.325 ;
        RECT 2471.670 2607.955 2471.950 2608.325 ;
        RECT 2470.820 2560.190 2470.960 2607.955 ;
        RECT 2470.760 2559.870 2471.020 2560.190 ;
        RECT 2472.140 2559.870 2472.400 2560.190 ;
        RECT 2472.200 2511.910 2472.340 2559.870 ;
        RECT 2471.220 2511.765 2471.480 2511.910 ;
        RECT 2469.830 2511.395 2470.110 2511.765 ;
        RECT 2471.210 2511.395 2471.490 2511.765 ;
        RECT 2472.140 2511.590 2472.400 2511.910 ;
        RECT 2469.900 2463.485 2470.040 2511.395 ;
        RECT 2469.830 2463.115 2470.110 2463.485 ;
        RECT 2470.750 2463.115 2471.030 2463.485 ;
        RECT 2470.820 2449.770 2470.960 2463.115 ;
        RECT 2470.820 2449.630 2471.420 2449.770 ;
        RECT 2471.280 2401.410 2471.420 2449.630 ;
        RECT 2470.300 2401.090 2470.560 2401.410 ;
        RECT 2471.220 2401.090 2471.480 2401.410 ;
        RECT 2470.360 2400.810 2470.500 2401.090 ;
        RECT 2470.360 2400.670 2470.960 2400.810 ;
        RECT 2470.820 2353.210 2470.960 2400.670 ;
        RECT 2470.820 2353.070 2471.420 2353.210 ;
        RECT 2471.280 2304.850 2471.420 2353.070 ;
        RECT 2470.300 2304.530 2470.560 2304.850 ;
        RECT 2471.220 2304.530 2471.480 2304.850 ;
        RECT 2470.360 2304.250 2470.500 2304.530 ;
        RECT 2470.360 2304.110 2470.960 2304.250 ;
        RECT 2470.820 2256.650 2470.960 2304.110 ;
        RECT 2470.820 2256.510 2471.420 2256.650 ;
        RECT 2471.280 2208.290 2471.420 2256.510 ;
        RECT 2470.300 2207.970 2470.560 2208.290 ;
        RECT 2471.220 2207.970 2471.480 2208.290 ;
        RECT 2470.360 2207.690 2470.500 2207.970 ;
        RECT 2470.360 2207.550 2470.960 2207.690 ;
        RECT 2470.820 2160.090 2470.960 2207.550 ;
        RECT 2470.820 2159.950 2471.420 2160.090 ;
        RECT 2471.280 2122.950 2471.420 2159.950 ;
        RECT 1795.020 2122.630 1795.280 2122.950 ;
        RECT 2471.220 2122.630 2471.480 2122.950 ;
        RECT 1795.080 2112.185 1795.220 2122.630 ;
        RECT 1795.080 2111.740 1795.430 2112.185 ;
        RECT 1795.150 2108.185 1795.430 2111.740 ;
      LAYER via2 ;
        RECT 2470.750 2801.120 2471.030 2801.400 ;
        RECT 2471.670 2801.120 2471.950 2801.400 ;
        RECT 2470.750 2704.560 2471.030 2704.840 ;
        RECT 2471.670 2704.560 2471.950 2704.840 ;
        RECT 2470.750 2608.000 2471.030 2608.280 ;
        RECT 2471.670 2608.000 2471.950 2608.280 ;
        RECT 2469.830 2511.440 2470.110 2511.720 ;
        RECT 2471.210 2511.440 2471.490 2511.720 ;
        RECT 2469.830 2463.160 2470.110 2463.440 ;
        RECT 2470.750 2463.160 2471.030 2463.440 ;
      LAYER met3 ;
        RECT 2470.725 2801.410 2471.055 2801.425 ;
        RECT 2471.645 2801.410 2471.975 2801.425 ;
        RECT 2470.725 2801.110 2471.975 2801.410 ;
        RECT 2470.725 2801.095 2471.055 2801.110 ;
        RECT 2471.645 2801.095 2471.975 2801.110 ;
        RECT 2470.725 2704.850 2471.055 2704.865 ;
        RECT 2471.645 2704.850 2471.975 2704.865 ;
        RECT 2470.725 2704.550 2471.975 2704.850 ;
        RECT 2470.725 2704.535 2471.055 2704.550 ;
        RECT 2471.645 2704.535 2471.975 2704.550 ;
        RECT 2470.725 2608.290 2471.055 2608.305 ;
        RECT 2471.645 2608.290 2471.975 2608.305 ;
        RECT 2470.725 2607.990 2471.975 2608.290 ;
        RECT 2470.725 2607.975 2471.055 2607.990 ;
        RECT 2471.645 2607.975 2471.975 2607.990 ;
        RECT 2469.805 2511.730 2470.135 2511.745 ;
        RECT 2471.185 2511.730 2471.515 2511.745 ;
        RECT 2469.805 2511.430 2471.515 2511.730 ;
        RECT 2469.805 2511.415 2470.135 2511.430 ;
        RECT 2471.185 2511.415 2471.515 2511.430 ;
        RECT 2469.805 2463.450 2470.135 2463.465 ;
        RECT 2470.725 2463.450 2471.055 2463.465 ;
        RECT 2469.805 2463.150 2471.055 2463.450 ;
        RECT 2469.805 2463.135 2470.135 2463.150 ;
        RECT 2470.725 2463.135 2471.055 2463.150 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3415.555 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
        RECT 2146.505 2753.065 2146.675 2801.175 ;
        RECT 2146.965 2428.705 2147.135 2463.215 ;
        RECT 2146.965 2331.805 2147.135 2366.655 ;
        RECT 2146.965 2138.685 2147.135 2173.535 ;
      LAYER mcon ;
        RECT 2147.885 3415.385 2148.055 3415.555 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
        RECT 2146.505 2801.005 2146.675 2801.175 ;
        RECT 2146.965 2463.045 2147.135 2463.215 ;
        RECT 2146.965 2366.485 2147.135 2366.655 ;
        RECT 2146.965 2173.365 2147.135 2173.535 ;
      LAYER met1 ;
        RECT 2145.970 3422.340 2146.290 3422.400 ;
        RECT 2149.190 3422.340 2149.510 3422.400 ;
        RECT 2145.970 3422.200 2149.510 3422.340 ;
        RECT 2145.970 3422.140 2146.290 3422.200 ;
        RECT 2149.190 3422.140 2149.510 3422.200 ;
        RECT 2145.970 3415.540 2146.290 3415.600 ;
        RECT 2147.825 3415.540 2148.115 3415.585 ;
        RECT 2145.970 3415.400 2148.115 3415.540 ;
        RECT 2145.970 3415.340 2146.290 3415.400 ;
        RECT 2147.825 3415.355 2148.115 3415.400 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2146.235 2801.020 2146.750 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2146.445 2753.220 2146.735 2753.265 ;
        RECT 2147.350 2753.220 2147.670 2753.280 ;
        RECT 2146.445 2753.080 2147.670 2753.220 ;
        RECT 2146.445 2753.035 2146.735 2753.080 ;
        RECT 2147.350 2753.020 2147.670 2753.080 ;
        RECT 2146.430 2718.200 2146.750 2718.260 ;
        RECT 2147.350 2718.200 2147.670 2718.260 ;
        RECT 2146.430 2718.060 2147.670 2718.200 ;
        RECT 2146.430 2718.000 2146.750 2718.060 ;
        RECT 2147.350 2718.000 2147.670 2718.060 ;
        RECT 2146.430 2670.260 2146.750 2670.320 ;
        RECT 2147.350 2670.260 2147.670 2670.320 ;
        RECT 2146.430 2670.120 2147.670 2670.260 ;
        RECT 2146.430 2670.060 2146.750 2670.120 ;
        RECT 2147.350 2670.060 2147.670 2670.120 ;
        RECT 2147.350 2622.120 2147.670 2622.380 ;
        RECT 2147.440 2621.980 2147.580 2622.120 ;
        RECT 2147.810 2621.980 2148.130 2622.040 ;
        RECT 2147.440 2621.840 2148.130 2621.980 ;
        RECT 2147.810 2621.780 2148.130 2621.840 ;
        RECT 2146.890 2560.100 2147.210 2560.160 ;
        RECT 2148.270 2560.100 2148.590 2560.160 ;
        RECT 2146.890 2559.960 2148.590 2560.100 ;
        RECT 2146.890 2559.900 2147.210 2559.960 ;
        RECT 2148.270 2559.900 2148.590 2559.960 ;
        RECT 2147.350 2511.820 2147.670 2511.880 ;
        RECT 2148.270 2511.820 2148.590 2511.880 ;
        RECT 2147.350 2511.680 2148.590 2511.820 ;
        RECT 2147.350 2511.620 2147.670 2511.680 ;
        RECT 2148.270 2511.620 2148.590 2511.680 ;
        RECT 2146.890 2463.200 2147.210 2463.260 ;
        RECT 2146.695 2463.060 2147.210 2463.200 ;
        RECT 2146.890 2463.000 2147.210 2463.060 ;
        RECT 2146.890 2428.860 2147.210 2428.920 ;
        RECT 2146.695 2428.720 2147.210 2428.860 ;
        RECT 2146.890 2428.660 2147.210 2428.720 ;
        RECT 2146.430 2380.580 2146.750 2380.640 ;
        RECT 2147.350 2380.580 2147.670 2380.640 ;
        RECT 2146.430 2380.440 2147.670 2380.580 ;
        RECT 2146.430 2380.380 2146.750 2380.440 ;
        RECT 2147.350 2380.380 2147.670 2380.440 ;
        RECT 2146.890 2366.640 2147.210 2366.700 ;
        RECT 2146.695 2366.500 2147.210 2366.640 ;
        RECT 2146.890 2366.440 2147.210 2366.500 ;
        RECT 2146.890 2331.960 2147.210 2332.020 ;
        RECT 2146.695 2331.820 2147.210 2331.960 ;
        RECT 2146.890 2331.760 2147.210 2331.820 ;
        RECT 2145.970 2235.540 2146.290 2235.800 ;
        RECT 2146.060 2235.400 2146.200 2235.540 ;
        RECT 2146.430 2235.400 2146.750 2235.460 ;
        RECT 2146.060 2235.260 2146.750 2235.400 ;
        RECT 2146.430 2235.200 2146.750 2235.260 ;
        RECT 2146.890 2173.520 2147.210 2173.580 ;
        RECT 2146.695 2173.380 2147.210 2173.520 ;
        RECT 2146.890 2173.320 2147.210 2173.380 ;
        RECT 2146.890 2138.840 2147.210 2138.900 ;
        RECT 2146.695 2138.700 2147.210 2138.840 ;
        RECT 2146.890 2138.640 2147.210 2138.700 ;
        RECT 1617.890 2123.880 1618.210 2123.940 ;
        RECT 2147.350 2123.880 2147.670 2123.940 ;
        RECT 1617.890 2123.740 2147.670 2123.880 ;
        RECT 1617.890 2123.680 1618.210 2123.740 ;
        RECT 2147.350 2123.680 2147.670 2123.740 ;
      LAYER via ;
        RECT 2146.000 3422.140 2146.260 3422.400 ;
        RECT 2149.220 3422.140 2149.480 3422.400 ;
        RECT 2146.000 3415.340 2146.260 3415.600 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2753.020 2147.640 2753.280 ;
        RECT 2146.460 2718.000 2146.720 2718.260 ;
        RECT 2147.380 2718.000 2147.640 2718.260 ;
        RECT 2146.460 2670.060 2146.720 2670.320 ;
        RECT 2147.380 2670.060 2147.640 2670.320 ;
        RECT 2147.380 2622.120 2147.640 2622.380 ;
        RECT 2147.840 2621.780 2148.100 2622.040 ;
        RECT 2146.920 2559.900 2147.180 2560.160 ;
        RECT 2148.300 2559.900 2148.560 2560.160 ;
        RECT 2147.380 2511.620 2147.640 2511.880 ;
        RECT 2148.300 2511.620 2148.560 2511.880 ;
        RECT 2146.920 2463.000 2147.180 2463.260 ;
        RECT 2146.920 2428.660 2147.180 2428.920 ;
        RECT 2146.460 2380.380 2146.720 2380.640 ;
        RECT 2147.380 2380.380 2147.640 2380.640 ;
        RECT 2146.920 2366.440 2147.180 2366.700 ;
        RECT 2146.920 2331.760 2147.180 2332.020 ;
        RECT 2146.000 2235.540 2146.260 2235.800 ;
        RECT 2146.460 2235.200 2146.720 2235.460 ;
        RECT 2146.920 2173.320 2147.180 2173.580 ;
        RECT 2146.920 2138.640 2147.180 2138.900 ;
        RECT 1617.920 2123.680 1618.180 2123.940 ;
        RECT 2147.380 2123.680 2147.640 2123.940 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3422.430 2149.420 3517.600 ;
        RECT 2146.000 3422.110 2146.260 3422.430 ;
        RECT 2149.220 3422.110 2149.480 3422.430 ;
        RECT 2146.060 3415.630 2146.200 3422.110 ;
        RECT 2146.000 3415.310 2146.260 3415.630 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.250 2146.660 2814.870 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2752.990 2147.640 2753.310 ;
        RECT 2147.440 2718.290 2147.580 2752.990 ;
        RECT 2146.460 2717.970 2146.720 2718.290 ;
        RECT 2147.380 2717.970 2147.640 2718.290 ;
        RECT 2146.520 2670.350 2146.660 2717.970 ;
        RECT 2146.460 2670.030 2146.720 2670.350 ;
        RECT 2147.380 2670.030 2147.640 2670.350 ;
        RECT 2147.440 2622.410 2147.580 2670.030 ;
        RECT 2147.380 2622.090 2147.640 2622.410 ;
        RECT 2147.840 2621.750 2148.100 2622.070 ;
        RECT 2147.900 2608.325 2148.040 2621.750 ;
        RECT 2146.910 2607.955 2147.190 2608.325 ;
        RECT 2147.830 2607.955 2148.110 2608.325 ;
        RECT 2146.980 2560.190 2147.120 2607.955 ;
        RECT 2146.920 2559.870 2147.180 2560.190 ;
        RECT 2148.300 2559.870 2148.560 2560.190 ;
        RECT 2148.360 2511.910 2148.500 2559.870 ;
        RECT 2147.380 2511.765 2147.640 2511.910 ;
        RECT 2145.990 2511.395 2146.270 2511.765 ;
        RECT 2147.370 2511.395 2147.650 2511.765 ;
        RECT 2148.300 2511.590 2148.560 2511.910 ;
        RECT 2146.060 2463.485 2146.200 2511.395 ;
        RECT 2145.990 2463.115 2146.270 2463.485 ;
        RECT 2146.910 2463.115 2147.190 2463.485 ;
        RECT 2146.920 2462.970 2147.180 2463.115 ;
        RECT 2146.920 2428.630 2147.180 2428.950 ;
        RECT 2146.980 2415.090 2147.120 2428.630 ;
        RECT 2146.980 2414.950 2147.580 2415.090 ;
        RECT 2147.440 2380.670 2147.580 2414.950 ;
        RECT 2146.460 2380.410 2146.720 2380.670 ;
        RECT 2146.460 2380.350 2147.120 2380.410 ;
        RECT 2147.380 2380.350 2147.640 2380.670 ;
        RECT 2146.520 2380.270 2147.120 2380.350 ;
        RECT 2146.980 2366.730 2147.120 2380.270 ;
        RECT 2146.920 2366.410 2147.180 2366.730 ;
        RECT 2146.920 2331.730 2147.180 2332.050 ;
        RECT 2146.980 2318.530 2147.120 2331.730 ;
        RECT 2146.980 2318.390 2147.580 2318.530 ;
        RECT 2147.440 2270.365 2147.580 2318.390 ;
        RECT 2145.990 2269.995 2146.270 2270.365 ;
        RECT 2147.370 2269.995 2147.650 2270.365 ;
        RECT 2146.060 2235.830 2146.200 2269.995 ;
        RECT 2146.000 2235.510 2146.260 2235.830 ;
        RECT 2146.460 2235.170 2146.720 2235.490 ;
        RECT 2146.520 2187.290 2146.660 2235.170 ;
        RECT 2146.520 2187.150 2147.120 2187.290 ;
        RECT 2146.980 2173.610 2147.120 2187.150 ;
        RECT 2146.920 2173.290 2147.180 2173.610 ;
        RECT 2146.920 2138.610 2147.180 2138.930 ;
        RECT 2146.980 2125.410 2147.120 2138.610 ;
        RECT 2146.980 2125.270 2147.580 2125.410 ;
        RECT 2147.440 2123.970 2147.580 2125.270 ;
        RECT 1617.920 2123.650 1618.180 2123.970 ;
        RECT 2147.380 2123.650 2147.640 2123.970 ;
        RECT 1617.980 2112.185 1618.120 2123.650 ;
        RECT 1617.980 2111.740 1618.330 2112.185 ;
        RECT 1618.050 2108.185 1618.330 2111.740 ;
      LAYER via2 ;
        RECT 2146.910 2608.000 2147.190 2608.280 ;
        RECT 2147.830 2608.000 2148.110 2608.280 ;
        RECT 2145.990 2511.440 2146.270 2511.720 ;
        RECT 2147.370 2511.440 2147.650 2511.720 ;
        RECT 2145.990 2463.160 2146.270 2463.440 ;
        RECT 2146.910 2463.160 2147.190 2463.440 ;
        RECT 2145.990 2270.040 2146.270 2270.320 ;
        RECT 2147.370 2270.040 2147.650 2270.320 ;
      LAYER met3 ;
        RECT 2146.885 2608.290 2147.215 2608.305 ;
        RECT 2147.805 2608.290 2148.135 2608.305 ;
        RECT 2146.885 2607.990 2148.135 2608.290 ;
        RECT 2146.885 2607.975 2147.215 2607.990 ;
        RECT 2147.805 2607.975 2148.135 2607.990 ;
        RECT 2145.965 2511.730 2146.295 2511.745 ;
        RECT 2147.345 2511.730 2147.675 2511.745 ;
        RECT 2145.965 2511.430 2147.675 2511.730 ;
        RECT 2145.965 2511.415 2146.295 2511.430 ;
        RECT 2147.345 2511.415 2147.675 2511.430 ;
        RECT 2145.965 2463.450 2146.295 2463.465 ;
        RECT 2146.885 2463.450 2147.215 2463.465 ;
        RECT 2145.965 2463.150 2147.215 2463.450 ;
        RECT 2145.965 2463.135 2146.295 2463.150 ;
        RECT 2146.885 2463.135 2147.215 2463.150 ;
        RECT 2145.965 2270.330 2146.295 2270.345 ;
        RECT 2147.345 2270.330 2147.675 2270.345 ;
        RECT 2145.965 2270.030 2147.675 2270.330 ;
        RECT 2145.965 2270.015 2146.295 2270.030 ;
        RECT 2147.345 2270.015 2147.675 2270.030 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 2898.245 1821.915 2946.355 ;
        RECT 1822.205 2815.285 1822.375 2849.455 ;
      LAYER mcon ;
        RECT 1821.745 2946.185 1821.915 2946.355 ;
        RECT 1822.205 2849.285 1822.375 2849.455 ;
      LAYER met1 ;
        RECT 1821.670 3464.160 1821.990 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1821.670 3464.020 1825.670 3464.160 ;
        RECT 1821.670 3463.960 1821.990 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1821.670 3367.600 1821.990 3367.660 ;
        RECT 1822.590 3367.600 1822.910 3367.660 ;
        RECT 1821.670 3367.460 1822.910 3367.600 ;
        RECT 1821.670 3367.400 1821.990 3367.460 ;
        RECT 1822.590 3367.400 1822.910 3367.460 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1821.685 2946.340 1821.975 2946.385 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1821.685 2946.200 1822.450 2946.340 ;
        RECT 1821.685 2946.155 1821.975 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1821.670 2898.400 1821.990 2898.460 ;
        RECT 1821.475 2898.260 1821.990 2898.400 ;
        RECT 1821.670 2898.200 1821.990 2898.260 ;
        RECT 1822.130 2849.440 1822.450 2849.500 ;
        RECT 1821.935 2849.300 1822.450 2849.440 ;
        RECT 1822.130 2849.240 1822.450 2849.300 ;
        RECT 1822.145 2815.440 1822.435 2815.485 ;
        RECT 1823.050 2815.440 1823.370 2815.500 ;
        RECT 1822.145 2815.300 1823.370 2815.440 ;
        RECT 1822.145 2815.255 1822.435 2815.300 ;
        RECT 1823.050 2815.240 1823.370 2815.300 ;
        RECT 1822.130 2753.220 1822.450 2753.280 ;
        RECT 1823.510 2753.220 1823.830 2753.280 ;
        RECT 1822.130 2753.080 1823.830 2753.220 ;
        RECT 1822.130 2753.020 1822.450 2753.080 ;
        RECT 1823.510 2753.020 1823.830 2753.080 ;
        RECT 1823.510 2719.220 1823.830 2719.280 ;
        RECT 1823.140 2719.080 1823.830 2719.220 ;
        RECT 1823.140 2718.600 1823.280 2719.080 ;
        RECT 1823.510 2719.020 1823.830 2719.080 ;
        RECT 1823.050 2718.340 1823.370 2718.600 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1823.510 2622.660 1823.830 2622.720 ;
        RECT 1823.140 2622.520 1823.830 2622.660 ;
        RECT 1823.140 2622.040 1823.280 2622.520 ;
        RECT 1823.510 2622.460 1823.830 2622.520 ;
        RECT 1823.050 2621.780 1823.370 2622.040 ;
        RECT 1822.130 2560.100 1822.450 2560.160 ;
        RECT 1823.510 2560.100 1823.830 2560.160 ;
        RECT 1822.130 2559.960 1823.830 2560.100 ;
        RECT 1822.130 2559.900 1822.450 2559.960 ;
        RECT 1823.510 2559.900 1823.830 2559.960 ;
        RECT 1822.590 2511.820 1822.910 2511.880 ;
        RECT 1823.510 2511.820 1823.830 2511.880 ;
        RECT 1822.590 2511.680 1823.830 2511.820 ;
        RECT 1822.590 2511.620 1822.910 2511.680 ;
        RECT 1823.510 2511.620 1823.830 2511.680 ;
        RECT 1821.670 2401.320 1821.990 2401.380 ;
        RECT 1822.590 2401.320 1822.910 2401.380 ;
        RECT 1821.670 2401.180 1822.910 2401.320 ;
        RECT 1821.670 2401.120 1821.990 2401.180 ;
        RECT 1822.590 2401.120 1822.910 2401.180 ;
        RECT 1821.670 2304.760 1821.990 2304.820 ;
        RECT 1822.590 2304.760 1822.910 2304.820 ;
        RECT 1821.670 2304.620 1822.910 2304.760 ;
        RECT 1821.670 2304.560 1821.990 2304.620 ;
        RECT 1822.590 2304.560 1822.910 2304.620 ;
        RECT 1821.670 2208.200 1821.990 2208.260 ;
        RECT 1822.590 2208.200 1822.910 2208.260 ;
        RECT 1821.670 2208.060 1822.910 2208.200 ;
        RECT 1821.670 2208.000 1821.990 2208.060 ;
        RECT 1822.590 2208.000 1822.910 2208.060 ;
        RECT 1441.250 2121.840 1441.570 2121.900 ;
        RECT 1822.590 2121.840 1822.910 2121.900 ;
        RECT 1441.250 2121.700 1822.910 2121.840 ;
        RECT 1441.250 2121.640 1441.570 2121.700 ;
        RECT 1822.590 2121.640 1822.910 2121.700 ;
      LAYER via ;
        RECT 1821.700 3463.960 1821.960 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1821.700 3367.400 1821.960 3367.660 ;
        RECT 1822.620 3367.400 1822.880 3367.660 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1821.700 2898.200 1821.960 2898.460 ;
        RECT 1822.160 2849.240 1822.420 2849.500 ;
        RECT 1823.080 2815.240 1823.340 2815.500 ;
        RECT 1822.160 2753.020 1822.420 2753.280 ;
        RECT 1823.540 2753.020 1823.800 2753.280 ;
        RECT 1823.540 2719.020 1823.800 2719.280 ;
        RECT 1823.080 2718.340 1823.340 2718.600 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1823.540 2622.460 1823.800 2622.720 ;
        RECT 1823.080 2621.780 1823.340 2622.040 ;
        RECT 1822.160 2559.900 1822.420 2560.160 ;
        RECT 1823.540 2559.900 1823.800 2560.160 ;
        RECT 1822.620 2511.620 1822.880 2511.880 ;
        RECT 1823.540 2511.620 1823.800 2511.880 ;
        RECT 1821.700 2401.120 1821.960 2401.380 ;
        RECT 1822.620 2401.120 1822.880 2401.380 ;
        RECT 1821.700 2304.560 1821.960 2304.820 ;
        RECT 1822.620 2304.560 1822.880 2304.820 ;
        RECT 1821.700 2208.000 1821.960 2208.260 ;
        RECT 1822.620 2208.000 1822.880 2208.260 ;
        RECT 1441.280 2121.640 1441.540 2121.900 ;
        RECT 1822.620 2121.640 1822.880 2121.900 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1821.700 3463.930 1821.960 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1821.760 3415.370 1821.900 3463.930 ;
        RECT 1821.760 3415.230 1822.820 3415.370 ;
        RECT 1822.680 3367.690 1822.820 3415.230 ;
        RECT 1821.700 3367.370 1821.960 3367.690 ;
        RECT 1822.620 3367.370 1822.880 3367.690 ;
        RECT 1821.760 3318.810 1821.900 3367.370 ;
        RECT 1821.760 3318.670 1822.820 3318.810 ;
        RECT 1822.680 3270.790 1822.820 3318.670 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1821.700 2898.170 1821.960 2898.490 ;
        RECT 1821.760 2863.210 1821.900 2898.170 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2849.530 1822.360 2863.070 ;
        RECT 1822.160 2849.210 1822.420 2849.530 ;
        RECT 1823.080 2815.210 1823.340 2815.530 ;
        RECT 1823.140 2801.445 1823.280 2815.210 ;
        RECT 1822.150 2801.075 1822.430 2801.445 ;
        RECT 1823.070 2801.075 1823.350 2801.445 ;
        RECT 1822.220 2753.310 1822.360 2801.075 ;
        RECT 1822.160 2752.990 1822.420 2753.310 ;
        RECT 1823.540 2752.990 1823.800 2753.310 ;
        RECT 1823.600 2719.310 1823.740 2752.990 ;
        RECT 1823.540 2718.990 1823.800 2719.310 ;
        RECT 1823.080 2718.310 1823.340 2718.630 ;
        RECT 1823.140 2704.885 1823.280 2718.310 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2622.750 1823.740 2656.430 ;
        RECT 1823.540 2622.430 1823.800 2622.750 ;
        RECT 1823.080 2621.750 1823.340 2622.070 ;
        RECT 1823.140 2608.325 1823.280 2621.750 ;
        RECT 1822.150 2607.955 1822.430 2608.325 ;
        RECT 1823.070 2607.955 1823.350 2608.325 ;
        RECT 1822.220 2560.190 1822.360 2607.955 ;
        RECT 1822.160 2559.870 1822.420 2560.190 ;
        RECT 1823.540 2559.870 1823.800 2560.190 ;
        RECT 1823.600 2511.910 1823.740 2559.870 ;
        RECT 1822.620 2511.765 1822.880 2511.910 ;
        RECT 1821.230 2511.395 1821.510 2511.765 ;
        RECT 1822.610 2511.395 1822.890 2511.765 ;
        RECT 1823.540 2511.590 1823.800 2511.910 ;
        RECT 1821.300 2463.485 1821.440 2511.395 ;
        RECT 1821.230 2463.115 1821.510 2463.485 ;
        RECT 1822.150 2463.115 1822.430 2463.485 ;
        RECT 1822.220 2449.770 1822.360 2463.115 ;
        RECT 1822.220 2449.630 1822.820 2449.770 ;
        RECT 1822.680 2401.410 1822.820 2449.630 ;
        RECT 1821.700 2401.090 1821.960 2401.410 ;
        RECT 1822.620 2401.090 1822.880 2401.410 ;
        RECT 1821.760 2400.810 1821.900 2401.090 ;
        RECT 1821.760 2400.670 1822.360 2400.810 ;
        RECT 1822.220 2353.210 1822.360 2400.670 ;
        RECT 1822.220 2353.070 1822.820 2353.210 ;
        RECT 1822.680 2304.850 1822.820 2353.070 ;
        RECT 1821.700 2304.530 1821.960 2304.850 ;
        RECT 1822.620 2304.530 1822.880 2304.850 ;
        RECT 1821.760 2304.250 1821.900 2304.530 ;
        RECT 1821.760 2304.110 1822.360 2304.250 ;
        RECT 1822.220 2256.650 1822.360 2304.110 ;
        RECT 1822.220 2256.510 1822.820 2256.650 ;
        RECT 1822.680 2208.290 1822.820 2256.510 ;
        RECT 1821.700 2207.970 1821.960 2208.290 ;
        RECT 1822.620 2207.970 1822.880 2208.290 ;
        RECT 1821.760 2207.690 1821.900 2207.970 ;
        RECT 1821.760 2207.550 1822.360 2207.690 ;
        RECT 1822.220 2160.090 1822.360 2207.550 ;
        RECT 1822.220 2159.950 1822.820 2160.090 ;
        RECT 1822.680 2121.930 1822.820 2159.950 ;
        RECT 1441.280 2121.610 1441.540 2121.930 ;
        RECT 1822.620 2121.610 1822.880 2121.930 ;
        RECT 1441.340 2112.185 1441.480 2121.610 ;
        RECT 1441.340 2111.740 1441.690 2112.185 ;
        RECT 1441.410 2108.185 1441.690 2111.740 ;
      LAYER via2 ;
        RECT 1822.150 2801.120 1822.430 2801.400 ;
        RECT 1823.070 2801.120 1823.350 2801.400 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
        RECT 1822.150 2608.000 1822.430 2608.280 ;
        RECT 1823.070 2608.000 1823.350 2608.280 ;
        RECT 1821.230 2511.440 1821.510 2511.720 ;
        RECT 1822.610 2511.440 1822.890 2511.720 ;
        RECT 1821.230 2463.160 1821.510 2463.440 ;
        RECT 1822.150 2463.160 1822.430 2463.440 ;
      LAYER met3 ;
        RECT 1822.125 2801.410 1822.455 2801.425 ;
        RECT 1823.045 2801.410 1823.375 2801.425 ;
        RECT 1822.125 2801.110 1823.375 2801.410 ;
        RECT 1822.125 2801.095 1822.455 2801.110 ;
        RECT 1823.045 2801.095 1823.375 2801.110 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
        RECT 1822.125 2608.290 1822.455 2608.305 ;
        RECT 1823.045 2608.290 1823.375 2608.305 ;
        RECT 1822.125 2607.990 1823.375 2608.290 ;
        RECT 1822.125 2607.975 1822.455 2607.990 ;
        RECT 1823.045 2607.975 1823.375 2607.990 ;
        RECT 1821.205 2511.730 1821.535 2511.745 ;
        RECT 1822.585 2511.730 1822.915 2511.745 ;
        RECT 1821.205 2511.430 1822.915 2511.730 ;
        RECT 1821.205 2511.415 1821.535 2511.430 ;
        RECT 1822.585 2511.415 1822.915 2511.430 ;
        RECT 1821.205 2463.450 1821.535 2463.465 ;
        RECT 1822.125 2463.450 1822.455 2463.465 ;
        RECT 1821.205 2463.150 1822.455 2463.450 ;
        RECT 1821.205 2463.135 1821.535 2463.150 ;
        RECT 1822.125 2463.135 1822.455 2463.150 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3415.555 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1499.285 2946.525 1499.455 2994.635 ;
        RECT 1498.365 2428.705 1498.535 2463.215 ;
        RECT 1498.365 2331.805 1498.535 2366.655 ;
        RECT 1497.905 2235.245 1498.075 2269.755 ;
        RECT 1498.365 2138.685 1498.535 2173.535 ;
      LAYER mcon ;
        RECT 1499.285 3415.385 1499.455 3415.555 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1499.285 2994.465 1499.455 2994.635 ;
        RECT 1498.365 2463.045 1498.535 2463.215 ;
        RECT 1498.365 2366.485 1498.535 2366.655 ;
        RECT 1497.905 2269.585 1498.075 2269.755 ;
        RECT 1498.365 2173.365 1498.535 2173.535 ;
      LAYER met1 ;
        RECT 1497.370 3422.340 1497.690 3422.400 ;
        RECT 1500.590 3422.340 1500.910 3422.400 ;
        RECT 1497.370 3422.200 1500.910 3422.340 ;
        RECT 1497.370 3422.140 1497.690 3422.200 ;
        RECT 1500.590 3422.140 1500.910 3422.200 ;
        RECT 1497.370 3415.540 1497.690 3415.600 ;
        RECT 1499.225 3415.540 1499.515 3415.585 ;
        RECT 1497.370 3415.400 1499.515 3415.540 ;
        RECT 1497.370 3415.340 1497.690 3415.400 ;
        RECT 1499.225 3415.355 1499.515 3415.400 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1499.015 2994.480 1499.530 2994.620 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.225 2946.680 1499.515 2946.725 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1499.225 2946.540 1499.990 2946.680 ;
        RECT 1499.225 2946.495 1499.515 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.370 2753.220 1497.690 2753.280 ;
        RECT 1498.750 2753.220 1499.070 2753.280 ;
        RECT 1497.370 2753.080 1499.070 2753.220 ;
        RECT 1497.370 2753.020 1497.690 2753.080 ;
        RECT 1498.750 2753.020 1499.070 2753.080 ;
        RECT 1497.370 2718.680 1497.690 2718.940 ;
        RECT 1497.460 2718.200 1497.600 2718.680 ;
        RECT 1497.830 2718.200 1498.150 2718.260 ;
        RECT 1497.460 2718.060 1498.150 2718.200 ;
        RECT 1497.830 2718.000 1498.150 2718.060 ;
        RECT 1497.830 2670.260 1498.150 2670.320 ;
        RECT 1498.750 2670.260 1499.070 2670.320 ;
        RECT 1497.830 2670.120 1499.070 2670.260 ;
        RECT 1497.830 2670.060 1498.150 2670.120 ;
        RECT 1498.750 2670.060 1499.070 2670.120 ;
        RECT 1498.750 2622.120 1499.070 2622.380 ;
        RECT 1498.840 2621.980 1498.980 2622.120 ;
        RECT 1499.210 2621.980 1499.530 2622.040 ;
        RECT 1498.840 2621.840 1499.530 2621.980 ;
        RECT 1499.210 2621.780 1499.530 2621.840 ;
        RECT 1498.290 2560.100 1498.610 2560.160 ;
        RECT 1499.670 2560.100 1499.990 2560.160 ;
        RECT 1498.290 2559.960 1499.990 2560.100 ;
        RECT 1498.290 2559.900 1498.610 2559.960 ;
        RECT 1499.670 2559.900 1499.990 2559.960 ;
        RECT 1498.750 2511.820 1499.070 2511.880 ;
        RECT 1499.670 2511.820 1499.990 2511.880 ;
        RECT 1498.750 2511.680 1499.990 2511.820 ;
        RECT 1498.750 2511.620 1499.070 2511.680 ;
        RECT 1499.670 2511.620 1499.990 2511.680 ;
        RECT 1498.290 2463.200 1498.610 2463.260 ;
        RECT 1498.095 2463.060 1498.610 2463.200 ;
        RECT 1498.290 2463.000 1498.610 2463.060 ;
        RECT 1498.290 2428.860 1498.610 2428.920 ;
        RECT 1498.095 2428.720 1498.610 2428.860 ;
        RECT 1498.290 2428.660 1498.610 2428.720 ;
        RECT 1497.830 2380.580 1498.150 2380.640 ;
        RECT 1498.750 2380.580 1499.070 2380.640 ;
        RECT 1497.830 2380.440 1499.070 2380.580 ;
        RECT 1497.830 2380.380 1498.150 2380.440 ;
        RECT 1498.750 2380.380 1499.070 2380.440 ;
        RECT 1498.290 2366.640 1498.610 2366.700 ;
        RECT 1498.095 2366.500 1498.610 2366.640 ;
        RECT 1498.290 2366.440 1498.610 2366.500 ;
        RECT 1498.290 2331.960 1498.610 2332.020 ;
        RECT 1498.095 2331.820 1498.610 2331.960 ;
        RECT 1498.290 2331.760 1498.610 2331.820 ;
        RECT 1497.830 2269.740 1498.150 2269.800 ;
        RECT 1497.635 2269.600 1498.150 2269.740 ;
        RECT 1497.830 2269.540 1498.150 2269.600 ;
        RECT 1497.830 2235.400 1498.150 2235.460 ;
        RECT 1497.635 2235.260 1498.150 2235.400 ;
        RECT 1497.830 2235.200 1498.150 2235.260 ;
        RECT 1498.290 2173.520 1498.610 2173.580 ;
        RECT 1498.095 2173.380 1498.610 2173.520 ;
        RECT 1498.290 2173.320 1498.610 2173.380 ;
        RECT 1498.290 2138.840 1498.610 2138.900 ;
        RECT 1498.095 2138.700 1498.610 2138.840 ;
        RECT 1498.290 2138.640 1498.610 2138.700 ;
        RECT 1264.610 2122.860 1264.930 2122.920 ;
        RECT 1498.750 2122.860 1499.070 2122.920 ;
        RECT 1264.610 2122.720 1499.070 2122.860 ;
        RECT 1264.610 2122.660 1264.930 2122.720 ;
        RECT 1498.750 2122.660 1499.070 2122.720 ;
      LAYER via ;
        RECT 1497.400 3422.140 1497.660 3422.400 ;
        RECT 1500.620 3422.140 1500.880 3422.400 ;
        RECT 1497.400 3415.340 1497.660 3415.600 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.400 2753.020 1497.660 2753.280 ;
        RECT 1498.780 2753.020 1499.040 2753.280 ;
        RECT 1497.400 2718.680 1497.660 2718.940 ;
        RECT 1497.860 2718.000 1498.120 2718.260 ;
        RECT 1497.860 2670.060 1498.120 2670.320 ;
        RECT 1498.780 2670.060 1499.040 2670.320 ;
        RECT 1498.780 2622.120 1499.040 2622.380 ;
        RECT 1499.240 2621.780 1499.500 2622.040 ;
        RECT 1498.320 2559.900 1498.580 2560.160 ;
        RECT 1499.700 2559.900 1499.960 2560.160 ;
        RECT 1498.780 2511.620 1499.040 2511.880 ;
        RECT 1499.700 2511.620 1499.960 2511.880 ;
        RECT 1498.320 2463.000 1498.580 2463.260 ;
        RECT 1498.320 2428.660 1498.580 2428.920 ;
        RECT 1497.860 2380.380 1498.120 2380.640 ;
        RECT 1498.780 2380.380 1499.040 2380.640 ;
        RECT 1498.320 2366.440 1498.580 2366.700 ;
        RECT 1498.320 2331.760 1498.580 2332.020 ;
        RECT 1497.860 2269.540 1498.120 2269.800 ;
        RECT 1497.860 2235.200 1498.120 2235.460 ;
        RECT 1498.320 2173.320 1498.580 2173.580 ;
        RECT 1498.320 2138.640 1498.580 2138.900 ;
        RECT 1264.640 2122.660 1264.900 2122.920 ;
        RECT 1498.780 2122.660 1499.040 2122.920 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3422.430 1500.820 3517.600 ;
        RECT 1497.400 3422.110 1497.660 3422.430 ;
        RECT 1500.620 3422.110 1500.880 3422.430 ;
        RECT 1497.460 3415.630 1497.600 3422.110 ;
        RECT 1497.400 3415.310 1497.660 3415.630 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.725 1498.520 2863.070 ;
        RECT 1498.310 2849.355 1498.590 2849.725 ;
        RECT 1497.850 2801.755 1498.130 2802.125 ;
        RECT 1497.920 2801.445 1498.060 2801.755 ;
        RECT 1497.850 2801.075 1498.130 2801.445 ;
        RECT 1498.770 2801.075 1499.050 2801.445 ;
        RECT 1498.840 2753.310 1498.980 2801.075 ;
        RECT 1497.400 2752.990 1497.660 2753.310 ;
        RECT 1498.780 2752.990 1499.040 2753.310 ;
        RECT 1497.460 2718.970 1497.600 2752.990 ;
        RECT 1497.400 2718.650 1497.660 2718.970 ;
        RECT 1497.860 2717.970 1498.120 2718.290 ;
        RECT 1497.920 2670.350 1498.060 2717.970 ;
        RECT 1497.860 2670.030 1498.120 2670.350 ;
        RECT 1498.780 2670.030 1499.040 2670.350 ;
        RECT 1498.840 2622.410 1498.980 2670.030 ;
        RECT 1498.780 2622.090 1499.040 2622.410 ;
        RECT 1499.240 2621.750 1499.500 2622.070 ;
        RECT 1499.300 2608.325 1499.440 2621.750 ;
        RECT 1498.310 2607.955 1498.590 2608.325 ;
        RECT 1499.230 2607.955 1499.510 2608.325 ;
        RECT 1498.380 2560.190 1498.520 2607.955 ;
        RECT 1498.320 2559.870 1498.580 2560.190 ;
        RECT 1499.700 2559.870 1499.960 2560.190 ;
        RECT 1499.760 2511.910 1499.900 2559.870 ;
        RECT 1498.780 2511.765 1499.040 2511.910 ;
        RECT 1497.390 2511.395 1497.670 2511.765 ;
        RECT 1498.770 2511.395 1499.050 2511.765 ;
        RECT 1499.700 2511.590 1499.960 2511.910 ;
        RECT 1497.460 2463.485 1497.600 2511.395 ;
        RECT 1497.390 2463.115 1497.670 2463.485 ;
        RECT 1498.310 2463.115 1498.590 2463.485 ;
        RECT 1498.320 2462.970 1498.580 2463.115 ;
        RECT 1498.320 2428.630 1498.580 2428.950 ;
        RECT 1498.380 2415.090 1498.520 2428.630 ;
        RECT 1498.380 2414.950 1498.980 2415.090 ;
        RECT 1498.840 2380.670 1498.980 2414.950 ;
        RECT 1497.860 2380.410 1498.120 2380.670 ;
        RECT 1497.860 2380.350 1498.520 2380.410 ;
        RECT 1498.780 2380.350 1499.040 2380.670 ;
        RECT 1497.920 2380.270 1498.520 2380.350 ;
        RECT 1498.380 2366.730 1498.520 2380.270 ;
        RECT 1498.320 2366.410 1498.580 2366.730 ;
        RECT 1498.320 2331.730 1498.580 2332.050 ;
        RECT 1498.380 2318.530 1498.520 2331.730 ;
        RECT 1498.380 2318.390 1498.980 2318.530 ;
        RECT 1498.840 2270.250 1498.980 2318.390 ;
        RECT 1497.920 2270.110 1498.980 2270.250 ;
        RECT 1497.920 2269.830 1498.060 2270.110 ;
        RECT 1497.860 2269.510 1498.120 2269.830 ;
        RECT 1497.860 2235.170 1498.120 2235.490 ;
        RECT 1497.920 2187.290 1498.060 2235.170 ;
        RECT 1497.920 2187.150 1498.520 2187.290 ;
        RECT 1498.380 2173.610 1498.520 2187.150 ;
        RECT 1498.320 2173.290 1498.580 2173.610 ;
        RECT 1498.320 2138.610 1498.580 2138.930 ;
        RECT 1498.380 2125.410 1498.520 2138.610 ;
        RECT 1498.380 2125.270 1498.980 2125.410 ;
        RECT 1498.840 2122.950 1498.980 2125.270 ;
        RECT 1264.640 2122.630 1264.900 2122.950 ;
        RECT 1498.780 2122.630 1499.040 2122.950 ;
        RECT 1264.700 2112.185 1264.840 2122.630 ;
        RECT 1264.700 2111.740 1265.050 2112.185 ;
        RECT 1264.770 2108.185 1265.050 2111.740 ;
      LAYER via2 ;
        RECT 1498.310 2849.400 1498.590 2849.680 ;
        RECT 1497.850 2801.800 1498.130 2802.080 ;
        RECT 1497.850 2801.120 1498.130 2801.400 ;
        RECT 1498.770 2801.120 1499.050 2801.400 ;
        RECT 1498.310 2608.000 1498.590 2608.280 ;
        RECT 1499.230 2608.000 1499.510 2608.280 ;
        RECT 1497.390 2511.440 1497.670 2511.720 ;
        RECT 1498.770 2511.440 1499.050 2511.720 ;
        RECT 1497.390 2463.160 1497.670 2463.440 ;
        RECT 1498.310 2463.160 1498.590 2463.440 ;
      LAYER met3 ;
        RECT 1498.285 2849.700 1498.615 2849.705 ;
        RECT 1498.030 2849.690 1498.615 2849.700 ;
        RECT 1497.830 2849.390 1498.615 2849.690 ;
        RECT 1498.030 2849.380 1498.615 2849.390 ;
        RECT 1498.285 2849.375 1498.615 2849.380 ;
        RECT 1497.825 2802.100 1498.155 2802.105 ;
        RECT 1497.825 2802.090 1498.410 2802.100 ;
        RECT 1497.600 2801.790 1498.410 2802.090 ;
        RECT 1497.825 2801.780 1498.410 2801.790 ;
        RECT 1497.825 2801.775 1498.155 2801.780 ;
        RECT 1497.825 2801.410 1498.155 2801.425 ;
        RECT 1498.745 2801.410 1499.075 2801.425 ;
        RECT 1497.825 2801.110 1499.075 2801.410 ;
        RECT 1497.825 2801.095 1498.155 2801.110 ;
        RECT 1498.745 2801.095 1499.075 2801.110 ;
        RECT 1498.285 2608.290 1498.615 2608.305 ;
        RECT 1499.205 2608.290 1499.535 2608.305 ;
        RECT 1498.285 2607.990 1499.535 2608.290 ;
        RECT 1498.285 2607.975 1498.615 2607.990 ;
        RECT 1499.205 2607.975 1499.535 2607.990 ;
        RECT 1497.365 2511.730 1497.695 2511.745 ;
        RECT 1498.745 2511.730 1499.075 2511.745 ;
        RECT 1497.365 2511.430 1499.075 2511.730 ;
        RECT 1497.365 2511.415 1497.695 2511.430 ;
        RECT 1498.745 2511.415 1499.075 2511.430 ;
        RECT 1497.365 2463.450 1497.695 2463.465 ;
        RECT 1498.285 2463.450 1498.615 2463.465 ;
        RECT 1497.365 2463.150 1498.615 2463.450 ;
        RECT 1497.365 2463.135 1497.695 2463.150 ;
        RECT 1498.285 2463.135 1498.615 2463.150 ;
      LAYER via3 ;
        RECT 1498.060 2849.380 1498.380 2849.700 ;
        RECT 1498.060 2801.780 1498.380 2802.100 ;
      LAYER met4 ;
        RECT 1498.055 2849.375 1498.385 2849.705 ;
        RECT 1498.070 2802.105 1498.370 2849.375 ;
        RECT 1498.055 2801.775 1498.385 2802.105 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.970 628.220 2008.290 628.280 ;
        RECT 2894.390 628.220 2894.710 628.280 ;
        RECT 2007.970 628.080 2894.710 628.220 ;
        RECT 2007.970 628.020 2008.290 628.080 ;
        RECT 2894.390 628.020 2894.710 628.080 ;
      LAYER via ;
        RECT 2008.000 628.020 2008.260 628.280 ;
        RECT 2894.420 628.020 2894.680 628.280 ;
      LAYER met2 ;
        RECT 2007.990 634.595 2008.270 634.965 ;
        RECT 2008.060 628.310 2008.200 634.595 ;
        RECT 2008.000 627.990 2008.260 628.310 ;
        RECT 2894.420 627.990 2894.680 628.310 ;
        RECT 2894.480 322.845 2894.620 627.990 ;
        RECT 2894.410 322.475 2894.690 322.845 ;
      LAYER via2 ;
        RECT 2007.990 634.640 2008.270 634.920 ;
        RECT 2894.410 322.520 2894.690 322.800 ;
      LAYER met3 ;
        RECT 1997.465 634.930 2001.465 635.080 ;
        RECT 2007.965 634.930 2008.295 634.945 ;
        RECT 1997.465 634.630 2008.295 634.930 ;
        RECT 1997.465 634.480 2001.465 634.630 ;
        RECT 2007.965 634.615 2008.295 634.630 ;
        RECT 2894.385 322.810 2894.715 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2894.385 322.510 2924.800 322.810 ;
        RECT 2894.385 322.495 2894.715 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1173.145 2898.245 1173.315 2946.355 ;
        RECT 1173.605 2815.285 1173.775 2849.455 ;
      LAYER mcon ;
        RECT 1173.145 2946.185 1173.315 2946.355 ;
        RECT 1173.605 2849.285 1173.775 2849.455 ;
      LAYER met1 ;
        RECT 1173.070 3464.160 1173.390 3464.220 ;
        RECT 1176.290 3464.160 1176.610 3464.220 ;
        RECT 1173.070 3464.020 1176.610 3464.160 ;
        RECT 1173.070 3463.960 1173.390 3464.020 ;
        RECT 1176.290 3463.960 1176.610 3464.020 ;
        RECT 1173.070 3367.600 1173.390 3367.660 ;
        RECT 1173.990 3367.600 1174.310 3367.660 ;
        RECT 1173.070 3367.460 1174.310 3367.600 ;
        RECT 1173.070 3367.400 1173.390 3367.460 ;
        RECT 1173.990 3367.400 1174.310 3367.460 ;
        RECT 1173.070 3270.700 1173.390 3270.760 ;
        RECT 1173.990 3270.700 1174.310 3270.760 ;
        RECT 1173.070 3270.560 1174.310 3270.700 ;
        RECT 1173.070 3270.500 1173.390 3270.560 ;
        RECT 1173.990 3270.500 1174.310 3270.560 ;
        RECT 1173.070 3174.140 1173.390 3174.200 ;
        RECT 1173.990 3174.140 1174.310 3174.200 ;
        RECT 1173.070 3174.000 1174.310 3174.140 ;
        RECT 1173.070 3173.940 1173.390 3174.000 ;
        RECT 1173.990 3173.940 1174.310 3174.000 ;
        RECT 1173.070 3077.580 1173.390 3077.640 ;
        RECT 1173.990 3077.580 1174.310 3077.640 ;
        RECT 1173.070 3077.440 1174.310 3077.580 ;
        RECT 1173.070 3077.380 1173.390 3077.440 ;
        RECT 1173.990 3077.380 1174.310 3077.440 ;
        RECT 1173.070 2981.020 1173.390 2981.080 ;
        RECT 1173.990 2981.020 1174.310 2981.080 ;
        RECT 1173.070 2980.880 1174.310 2981.020 ;
        RECT 1173.070 2980.820 1173.390 2980.880 ;
        RECT 1173.990 2980.820 1174.310 2980.880 ;
        RECT 1173.085 2946.340 1173.375 2946.385 ;
        RECT 1173.530 2946.340 1173.850 2946.400 ;
        RECT 1173.085 2946.200 1173.850 2946.340 ;
        RECT 1173.085 2946.155 1173.375 2946.200 ;
        RECT 1173.530 2946.140 1173.850 2946.200 ;
        RECT 1173.070 2898.400 1173.390 2898.460 ;
        RECT 1172.875 2898.260 1173.390 2898.400 ;
        RECT 1173.070 2898.200 1173.390 2898.260 ;
        RECT 1173.530 2849.440 1173.850 2849.500 ;
        RECT 1173.335 2849.300 1173.850 2849.440 ;
        RECT 1173.530 2849.240 1173.850 2849.300 ;
        RECT 1173.545 2815.440 1173.835 2815.485 ;
        RECT 1174.450 2815.440 1174.770 2815.500 ;
        RECT 1173.545 2815.300 1174.770 2815.440 ;
        RECT 1173.545 2815.255 1173.835 2815.300 ;
        RECT 1174.450 2815.240 1174.770 2815.300 ;
        RECT 1173.530 2753.220 1173.850 2753.280 ;
        RECT 1174.910 2753.220 1175.230 2753.280 ;
        RECT 1173.530 2753.080 1175.230 2753.220 ;
        RECT 1173.530 2753.020 1173.850 2753.080 ;
        RECT 1174.910 2753.020 1175.230 2753.080 ;
        RECT 1174.910 2719.220 1175.230 2719.280 ;
        RECT 1174.540 2719.080 1175.230 2719.220 ;
        RECT 1174.540 2718.600 1174.680 2719.080 ;
        RECT 1174.910 2719.020 1175.230 2719.080 ;
        RECT 1174.450 2718.340 1174.770 2718.600 ;
        RECT 1173.530 2656.660 1173.850 2656.720 ;
        RECT 1174.910 2656.660 1175.230 2656.720 ;
        RECT 1173.530 2656.520 1175.230 2656.660 ;
        RECT 1173.530 2656.460 1173.850 2656.520 ;
        RECT 1174.910 2656.460 1175.230 2656.520 ;
        RECT 1174.910 2622.660 1175.230 2622.720 ;
        RECT 1174.540 2622.520 1175.230 2622.660 ;
        RECT 1174.540 2622.040 1174.680 2622.520 ;
        RECT 1174.910 2622.460 1175.230 2622.520 ;
        RECT 1174.450 2621.780 1174.770 2622.040 ;
        RECT 1173.530 2560.100 1173.850 2560.160 ;
        RECT 1174.910 2560.100 1175.230 2560.160 ;
        RECT 1173.530 2559.960 1175.230 2560.100 ;
        RECT 1173.530 2559.900 1173.850 2559.960 ;
        RECT 1174.910 2559.900 1175.230 2559.960 ;
        RECT 1173.990 2511.820 1174.310 2511.880 ;
        RECT 1174.910 2511.820 1175.230 2511.880 ;
        RECT 1173.990 2511.680 1175.230 2511.820 ;
        RECT 1173.990 2511.620 1174.310 2511.680 ;
        RECT 1174.910 2511.620 1175.230 2511.680 ;
        RECT 1173.070 2401.320 1173.390 2401.380 ;
        RECT 1173.990 2401.320 1174.310 2401.380 ;
        RECT 1173.070 2401.180 1174.310 2401.320 ;
        RECT 1173.070 2401.120 1173.390 2401.180 ;
        RECT 1173.990 2401.120 1174.310 2401.180 ;
        RECT 1173.070 2304.760 1173.390 2304.820 ;
        RECT 1173.990 2304.760 1174.310 2304.820 ;
        RECT 1173.070 2304.620 1174.310 2304.760 ;
        RECT 1173.070 2304.560 1173.390 2304.620 ;
        RECT 1173.990 2304.560 1174.310 2304.620 ;
        RECT 1173.070 2208.200 1173.390 2208.260 ;
        RECT 1173.990 2208.200 1174.310 2208.260 ;
        RECT 1173.070 2208.060 1174.310 2208.200 ;
        RECT 1173.070 2208.000 1173.390 2208.060 ;
        RECT 1173.990 2208.000 1174.310 2208.060 ;
        RECT 1087.510 2121.840 1087.830 2121.900 ;
        RECT 1173.990 2121.840 1174.310 2121.900 ;
        RECT 1087.510 2121.700 1174.310 2121.840 ;
        RECT 1087.510 2121.640 1087.830 2121.700 ;
        RECT 1173.990 2121.640 1174.310 2121.700 ;
      LAYER via ;
        RECT 1173.100 3463.960 1173.360 3464.220 ;
        RECT 1176.320 3463.960 1176.580 3464.220 ;
        RECT 1173.100 3367.400 1173.360 3367.660 ;
        RECT 1174.020 3367.400 1174.280 3367.660 ;
        RECT 1173.100 3270.500 1173.360 3270.760 ;
        RECT 1174.020 3270.500 1174.280 3270.760 ;
        RECT 1173.100 3173.940 1173.360 3174.200 ;
        RECT 1174.020 3173.940 1174.280 3174.200 ;
        RECT 1173.100 3077.380 1173.360 3077.640 ;
        RECT 1174.020 3077.380 1174.280 3077.640 ;
        RECT 1173.100 2980.820 1173.360 2981.080 ;
        RECT 1174.020 2980.820 1174.280 2981.080 ;
        RECT 1173.560 2946.140 1173.820 2946.400 ;
        RECT 1173.100 2898.200 1173.360 2898.460 ;
        RECT 1173.560 2849.240 1173.820 2849.500 ;
        RECT 1174.480 2815.240 1174.740 2815.500 ;
        RECT 1173.560 2753.020 1173.820 2753.280 ;
        RECT 1174.940 2753.020 1175.200 2753.280 ;
        RECT 1174.940 2719.020 1175.200 2719.280 ;
        RECT 1174.480 2718.340 1174.740 2718.600 ;
        RECT 1173.560 2656.460 1173.820 2656.720 ;
        RECT 1174.940 2656.460 1175.200 2656.720 ;
        RECT 1174.940 2622.460 1175.200 2622.720 ;
        RECT 1174.480 2621.780 1174.740 2622.040 ;
        RECT 1173.560 2559.900 1173.820 2560.160 ;
        RECT 1174.940 2559.900 1175.200 2560.160 ;
        RECT 1174.020 2511.620 1174.280 2511.880 ;
        RECT 1174.940 2511.620 1175.200 2511.880 ;
        RECT 1173.100 2401.120 1173.360 2401.380 ;
        RECT 1174.020 2401.120 1174.280 2401.380 ;
        RECT 1173.100 2304.560 1173.360 2304.820 ;
        RECT 1174.020 2304.560 1174.280 2304.820 ;
        RECT 1173.100 2208.000 1173.360 2208.260 ;
        RECT 1174.020 2208.000 1174.280 2208.260 ;
        RECT 1087.540 2121.640 1087.800 2121.900 ;
        RECT 1174.020 2121.640 1174.280 2121.900 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3517.370 1176.060 3517.600 ;
        RECT 1175.920 3517.230 1176.520 3517.370 ;
        RECT 1176.380 3464.250 1176.520 3517.230 ;
        RECT 1173.100 3463.930 1173.360 3464.250 ;
        RECT 1176.320 3463.930 1176.580 3464.250 ;
        RECT 1173.160 3415.370 1173.300 3463.930 ;
        RECT 1173.160 3415.230 1174.220 3415.370 ;
        RECT 1174.080 3367.690 1174.220 3415.230 ;
        RECT 1173.100 3367.370 1173.360 3367.690 ;
        RECT 1174.020 3367.370 1174.280 3367.690 ;
        RECT 1173.160 3318.810 1173.300 3367.370 ;
        RECT 1173.160 3318.670 1174.220 3318.810 ;
        RECT 1174.080 3270.790 1174.220 3318.670 ;
        RECT 1173.100 3270.470 1173.360 3270.790 ;
        RECT 1174.020 3270.470 1174.280 3270.790 ;
        RECT 1173.160 3222.250 1173.300 3270.470 ;
        RECT 1173.160 3222.110 1174.220 3222.250 ;
        RECT 1174.080 3174.230 1174.220 3222.110 ;
        RECT 1173.100 3173.910 1173.360 3174.230 ;
        RECT 1174.020 3173.910 1174.280 3174.230 ;
        RECT 1173.160 3125.690 1173.300 3173.910 ;
        RECT 1173.160 3125.550 1174.220 3125.690 ;
        RECT 1174.080 3077.670 1174.220 3125.550 ;
        RECT 1173.100 3077.350 1173.360 3077.670 ;
        RECT 1174.020 3077.350 1174.280 3077.670 ;
        RECT 1173.160 3029.130 1173.300 3077.350 ;
        RECT 1173.160 3028.990 1174.220 3029.130 ;
        RECT 1174.080 2981.110 1174.220 3028.990 ;
        RECT 1173.100 2980.850 1173.360 2981.110 ;
        RECT 1173.100 2980.790 1173.760 2980.850 ;
        RECT 1174.020 2980.790 1174.280 2981.110 ;
        RECT 1173.160 2980.710 1173.760 2980.790 ;
        RECT 1173.620 2980.170 1173.760 2980.710 ;
        RECT 1173.620 2980.030 1174.220 2980.170 ;
        RECT 1174.080 2959.770 1174.220 2980.030 ;
        RECT 1173.620 2959.630 1174.220 2959.770 ;
        RECT 1173.620 2946.430 1173.760 2959.630 ;
        RECT 1173.560 2946.110 1173.820 2946.430 ;
        RECT 1173.100 2898.170 1173.360 2898.490 ;
        RECT 1173.160 2863.210 1173.300 2898.170 ;
        RECT 1173.160 2863.070 1173.760 2863.210 ;
        RECT 1173.620 2849.530 1173.760 2863.070 ;
        RECT 1173.560 2849.210 1173.820 2849.530 ;
        RECT 1174.480 2815.210 1174.740 2815.530 ;
        RECT 1174.540 2801.445 1174.680 2815.210 ;
        RECT 1173.550 2801.075 1173.830 2801.445 ;
        RECT 1174.470 2801.075 1174.750 2801.445 ;
        RECT 1173.620 2753.310 1173.760 2801.075 ;
        RECT 1173.560 2752.990 1173.820 2753.310 ;
        RECT 1174.940 2752.990 1175.200 2753.310 ;
        RECT 1175.000 2719.310 1175.140 2752.990 ;
        RECT 1174.940 2718.990 1175.200 2719.310 ;
        RECT 1174.480 2718.310 1174.740 2718.630 ;
        RECT 1174.540 2704.885 1174.680 2718.310 ;
        RECT 1173.550 2704.515 1173.830 2704.885 ;
        RECT 1174.470 2704.515 1174.750 2704.885 ;
        RECT 1173.620 2656.750 1173.760 2704.515 ;
        RECT 1173.560 2656.430 1173.820 2656.750 ;
        RECT 1174.940 2656.430 1175.200 2656.750 ;
        RECT 1175.000 2622.750 1175.140 2656.430 ;
        RECT 1174.940 2622.430 1175.200 2622.750 ;
        RECT 1174.480 2621.750 1174.740 2622.070 ;
        RECT 1174.540 2608.325 1174.680 2621.750 ;
        RECT 1173.550 2607.955 1173.830 2608.325 ;
        RECT 1174.470 2607.955 1174.750 2608.325 ;
        RECT 1173.620 2560.190 1173.760 2607.955 ;
        RECT 1173.560 2559.870 1173.820 2560.190 ;
        RECT 1174.940 2559.870 1175.200 2560.190 ;
        RECT 1175.000 2511.910 1175.140 2559.870 ;
        RECT 1174.020 2511.765 1174.280 2511.910 ;
        RECT 1172.630 2511.395 1172.910 2511.765 ;
        RECT 1174.010 2511.395 1174.290 2511.765 ;
        RECT 1174.940 2511.590 1175.200 2511.910 ;
        RECT 1172.700 2463.485 1172.840 2511.395 ;
        RECT 1172.630 2463.115 1172.910 2463.485 ;
        RECT 1173.550 2463.115 1173.830 2463.485 ;
        RECT 1173.620 2449.770 1173.760 2463.115 ;
        RECT 1173.620 2449.630 1174.220 2449.770 ;
        RECT 1174.080 2401.410 1174.220 2449.630 ;
        RECT 1173.100 2401.090 1173.360 2401.410 ;
        RECT 1174.020 2401.090 1174.280 2401.410 ;
        RECT 1173.160 2400.810 1173.300 2401.090 ;
        RECT 1173.160 2400.670 1173.760 2400.810 ;
        RECT 1173.620 2353.210 1173.760 2400.670 ;
        RECT 1173.620 2353.070 1174.220 2353.210 ;
        RECT 1174.080 2304.850 1174.220 2353.070 ;
        RECT 1173.100 2304.530 1173.360 2304.850 ;
        RECT 1174.020 2304.530 1174.280 2304.850 ;
        RECT 1173.160 2304.250 1173.300 2304.530 ;
        RECT 1173.160 2304.110 1173.760 2304.250 ;
        RECT 1173.620 2256.650 1173.760 2304.110 ;
        RECT 1173.620 2256.510 1174.220 2256.650 ;
        RECT 1174.080 2208.290 1174.220 2256.510 ;
        RECT 1173.100 2207.970 1173.360 2208.290 ;
        RECT 1174.020 2207.970 1174.280 2208.290 ;
        RECT 1173.160 2207.690 1173.300 2207.970 ;
        RECT 1173.160 2207.550 1173.760 2207.690 ;
        RECT 1173.620 2160.090 1173.760 2207.550 ;
        RECT 1173.620 2159.950 1174.220 2160.090 ;
        RECT 1174.080 2121.930 1174.220 2159.950 ;
        RECT 1087.540 2121.610 1087.800 2121.930 ;
        RECT 1174.020 2121.610 1174.280 2121.930 ;
        RECT 1087.600 2112.185 1087.740 2121.610 ;
        RECT 1087.600 2111.740 1087.950 2112.185 ;
        RECT 1087.670 2108.185 1087.950 2111.740 ;
      LAYER via2 ;
        RECT 1173.550 2801.120 1173.830 2801.400 ;
        RECT 1174.470 2801.120 1174.750 2801.400 ;
        RECT 1173.550 2704.560 1173.830 2704.840 ;
        RECT 1174.470 2704.560 1174.750 2704.840 ;
        RECT 1173.550 2608.000 1173.830 2608.280 ;
        RECT 1174.470 2608.000 1174.750 2608.280 ;
        RECT 1172.630 2511.440 1172.910 2511.720 ;
        RECT 1174.010 2511.440 1174.290 2511.720 ;
        RECT 1172.630 2463.160 1172.910 2463.440 ;
        RECT 1173.550 2463.160 1173.830 2463.440 ;
      LAYER met3 ;
        RECT 1173.525 2801.410 1173.855 2801.425 ;
        RECT 1174.445 2801.410 1174.775 2801.425 ;
        RECT 1173.525 2801.110 1174.775 2801.410 ;
        RECT 1173.525 2801.095 1173.855 2801.110 ;
        RECT 1174.445 2801.095 1174.775 2801.110 ;
        RECT 1173.525 2704.850 1173.855 2704.865 ;
        RECT 1174.445 2704.850 1174.775 2704.865 ;
        RECT 1173.525 2704.550 1174.775 2704.850 ;
        RECT 1173.525 2704.535 1173.855 2704.550 ;
        RECT 1174.445 2704.535 1174.775 2704.550 ;
        RECT 1173.525 2608.290 1173.855 2608.305 ;
        RECT 1174.445 2608.290 1174.775 2608.305 ;
        RECT 1173.525 2607.990 1174.775 2608.290 ;
        RECT 1173.525 2607.975 1173.855 2607.990 ;
        RECT 1174.445 2607.975 1174.775 2607.990 ;
        RECT 1172.605 2511.730 1172.935 2511.745 ;
        RECT 1173.985 2511.730 1174.315 2511.745 ;
        RECT 1172.605 2511.430 1174.315 2511.730 ;
        RECT 1172.605 2511.415 1172.935 2511.430 ;
        RECT 1173.985 2511.415 1174.315 2511.430 ;
        RECT 1172.605 2463.450 1172.935 2463.465 ;
        RECT 1173.525 2463.450 1173.855 2463.465 ;
        RECT 1172.605 2463.150 1173.855 2463.450 ;
        RECT 1172.605 2463.135 1172.935 2463.150 ;
        RECT 1173.525 2463.135 1173.855 2463.150 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 2121.840 855.530 2121.900 ;
        RECT 910.870 2121.840 911.190 2121.900 ;
        RECT 855.210 2121.700 911.190 2121.840 ;
        RECT 855.210 2121.640 855.530 2121.700 ;
        RECT 910.870 2121.640 911.190 2121.700 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 2121.640 855.500 2121.900 ;
        RECT 910.900 2121.640 911.160 2121.900 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 2121.930 855.440 3500.990 ;
        RECT 855.240 2121.610 855.500 2121.930 ;
        RECT 910.900 2121.610 911.160 2121.930 ;
        RECT 910.960 2112.185 911.100 2121.610 ;
        RECT 910.960 2111.740 911.310 2112.185 ;
        RECT 911.030 2108.185 911.310 2111.740 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 2122.180 531.230 2122.240 ;
        RECT 733.770 2122.180 734.090 2122.240 ;
        RECT 530.910 2122.040 734.090 2122.180 ;
        RECT 530.910 2121.980 531.230 2122.040 ;
        RECT 733.770 2121.980 734.090 2122.040 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 2121.980 531.200 2122.240 ;
        RECT 733.800 2121.980 734.060 2122.240 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2122.270 531.140 3498.270 ;
        RECT 530.940 2121.950 531.200 2122.270 ;
        RECT 733.800 2121.950 734.060 2122.270 ;
        RECT 733.860 2112.185 734.000 2121.950 ;
        RECT 733.860 2111.740 734.210 2112.185 ;
        RECT 733.930 2108.185 734.210 2111.740 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 2122.520 206.930 2122.580 ;
        RECT 557.130 2122.520 557.450 2122.580 ;
        RECT 206.610 2122.380 557.450 2122.520 ;
        RECT 206.610 2122.320 206.930 2122.380 ;
        RECT 557.130 2122.320 557.450 2122.380 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 2122.320 206.900 2122.580 ;
        RECT 557.160 2122.320 557.420 2122.580 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 2122.610 206.840 3501.670 ;
        RECT 206.640 2122.290 206.900 2122.610 ;
        RECT 557.160 2122.290 557.420 2122.610 ;
        RECT 557.220 2112.185 557.360 2122.290 ;
        RECT 557.220 2111.740 557.570 2112.185 ;
        RECT 557.290 2108.185 557.570 2111.740 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 44.690 3408.740 45.010 3408.800 ;
        RECT 17.550 3408.600 45.010 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 44.690 3408.540 45.010 3408.600 ;
        RECT 44.690 2097.360 45.010 2097.420 ;
        RECT 393.370 2097.360 393.690 2097.420 ;
        RECT 44.690 2097.220 393.690 2097.360 ;
        RECT 44.690 2097.160 45.010 2097.220 ;
        RECT 393.370 2097.160 393.690 2097.220 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 44.720 3408.540 44.980 3408.800 ;
        RECT 44.720 2097.160 44.980 2097.420 ;
        RECT 393.400 2097.160 393.660 2097.420 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 44.720 3408.510 44.980 3408.830 ;
        RECT 44.780 2097.450 44.920 3408.510 ;
        RECT 44.720 2097.130 44.980 2097.450 ;
        RECT 393.400 2097.130 393.660 2097.450 ;
        RECT 393.460 2092.885 393.600 2097.130 ;
        RECT 393.390 2092.515 393.670 2092.885 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 393.390 2092.560 393.670 2092.840 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 393.365 2092.850 393.695 2092.865 ;
        RECT 410.000 2092.850 414.000 2093.000 ;
        RECT 393.365 2092.550 414.000 2092.850 ;
        RECT 393.365 2092.535 393.695 2092.550 ;
        RECT 410.000 2092.400 414.000 2092.550 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 148.190 3119.060 148.510 3119.120 ;
        RECT 16.170 3118.920 148.510 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 148.190 3118.860 148.510 3118.920 ;
        RECT 148.190 1980.060 148.510 1980.120 ;
        RECT 393.370 1980.060 393.690 1980.120 ;
        RECT 148.190 1979.920 393.690 1980.060 ;
        RECT 148.190 1979.860 148.510 1979.920 ;
        RECT 393.370 1979.860 393.690 1979.920 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 148.220 3118.860 148.480 3119.120 ;
        RECT 148.220 1979.860 148.480 1980.120 ;
        RECT 393.400 1979.860 393.660 1980.120 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 148.220 3118.830 148.480 3119.150 ;
        RECT 148.280 1980.150 148.420 3118.830 ;
        RECT 148.220 1979.830 148.480 1980.150 ;
        RECT 393.400 1979.830 393.660 1980.150 ;
        RECT 393.460 1978.645 393.600 1979.830 ;
        RECT 393.390 1978.275 393.670 1978.645 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
        RECT 393.390 1978.320 393.670 1978.600 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
        RECT 393.365 1978.610 393.695 1978.625 ;
        RECT 410.000 1978.610 414.000 1978.760 ;
        RECT 393.365 1978.310 414.000 1978.610 ;
        RECT 393.365 1978.295 393.695 1978.310 ;
        RECT 410.000 1978.160 414.000 1978.310 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2836.180 20.630 2836.240 ;
        RECT 65.390 2836.180 65.710 2836.240 ;
        RECT 20.310 2836.040 65.710 2836.180 ;
        RECT 20.310 2835.980 20.630 2836.040 ;
        RECT 65.390 2835.980 65.710 2836.040 ;
        RECT 65.390 1869.900 65.710 1869.960 ;
        RECT 393.370 1869.900 393.690 1869.960 ;
        RECT 65.390 1869.760 393.690 1869.900 ;
        RECT 65.390 1869.700 65.710 1869.760 ;
        RECT 393.370 1869.700 393.690 1869.760 ;
      LAYER via ;
        RECT 20.340 2835.980 20.600 2836.240 ;
        RECT 65.420 2835.980 65.680 2836.240 ;
        RECT 65.420 1869.700 65.680 1869.960 ;
        RECT 393.400 1869.700 393.660 1869.960 ;
      LAYER met2 ;
        RECT 20.330 2836.435 20.610 2836.805 ;
        RECT 20.400 2836.270 20.540 2836.435 ;
        RECT 20.340 2835.950 20.600 2836.270 ;
        RECT 65.420 2835.950 65.680 2836.270 ;
        RECT 65.480 1869.990 65.620 2835.950 ;
        RECT 65.420 1869.670 65.680 1869.990 ;
        RECT 393.400 1869.670 393.660 1869.990 ;
        RECT 393.460 1864.405 393.600 1869.670 ;
        RECT 393.390 1864.035 393.670 1864.405 ;
      LAYER via2 ;
        RECT 20.330 2836.480 20.610 2836.760 ;
        RECT 393.390 1864.080 393.670 1864.360 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 20.305 2836.770 20.635 2836.785 ;
        RECT -4.800 2836.470 20.635 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 20.305 2836.455 20.635 2836.470 ;
        RECT 393.365 1864.370 393.695 1864.385 ;
        RECT 410.000 1864.370 414.000 1864.520 ;
        RECT 393.365 1864.070 414.000 1864.370 ;
        RECT 393.365 1864.055 393.695 1864.070 ;
        RECT 410.000 1863.920 414.000 1864.070 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 2546.500 19.710 2546.560 ;
        RECT 196.490 2546.500 196.810 2546.560 ;
        RECT 19.390 2546.360 196.810 2546.500 ;
        RECT 19.390 2546.300 19.710 2546.360 ;
        RECT 196.490 2546.300 196.810 2546.360 ;
        RECT 196.490 1752.600 196.810 1752.660 ;
        RECT 393.370 1752.600 393.690 1752.660 ;
        RECT 196.490 1752.460 393.690 1752.600 ;
        RECT 196.490 1752.400 196.810 1752.460 ;
        RECT 393.370 1752.400 393.690 1752.460 ;
      LAYER via ;
        RECT 19.420 2546.300 19.680 2546.560 ;
        RECT 196.520 2546.300 196.780 2546.560 ;
        RECT 196.520 1752.400 196.780 1752.660 ;
        RECT 393.400 1752.400 393.660 1752.660 ;
      LAYER met2 ;
        RECT 19.410 2549.475 19.690 2549.845 ;
        RECT 19.480 2546.590 19.620 2549.475 ;
        RECT 19.420 2546.270 19.680 2546.590 ;
        RECT 196.520 2546.270 196.780 2546.590 ;
        RECT 196.580 1752.690 196.720 2546.270 ;
        RECT 196.520 1752.370 196.780 1752.690 ;
        RECT 393.400 1752.370 393.660 1752.690 ;
        RECT 393.460 1750.165 393.600 1752.370 ;
        RECT 393.390 1749.795 393.670 1750.165 ;
      LAYER via2 ;
        RECT 19.410 2549.520 19.690 2549.800 ;
        RECT 393.390 1749.840 393.670 1750.120 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 19.385 2549.810 19.715 2549.825 ;
        RECT -4.800 2549.510 19.715 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 19.385 2549.495 19.715 2549.510 ;
        RECT 393.365 1750.130 393.695 1750.145 ;
        RECT 410.000 1750.130 414.000 1750.280 ;
        RECT 393.365 1749.830 414.000 1750.130 ;
        RECT 393.365 1749.815 393.695 1749.830 ;
        RECT 410.000 1749.680 414.000 1749.830 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 2256.480 15.570 2256.540 ;
        RECT 30.890 2256.480 31.210 2256.540 ;
        RECT 15.250 2256.340 31.210 2256.480 ;
        RECT 15.250 2256.280 15.570 2256.340 ;
        RECT 30.890 2256.280 31.210 2256.340 ;
        RECT 30.890 1635.300 31.210 1635.360 ;
        RECT 393.370 1635.300 393.690 1635.360 ;
        RECT 30.890 1635.160 393.690 1635.300 ;
        RECT 30.890 1635.100 31.210 1635.160 ;
        RECT 393.370 1635.100 393.690 1635.160 ;
      LAYER via ;
        RECT 15.280 2256.280 15.540 2256.540 ;
        RECT 30.920 2256.280 31.180 2256.540 ;
        RECT 30.920 1635.100 31.180 1635.360 ;
        RECT 393.400 1635.100 393.660 1635.360 ;
      LAYER met2 ;
        RECT 15.270 2261.835 15.550 2262.205 ;
        RECT 15.340 2256.570 15.480 2261.835 ;
        RECT 15.280 2256.250 15.540 2256.570 ;
        RECT 30.920 2256.250 31.180 2256.570 ;
        RECT 30.980 1635.390 31.120 2256.250 ;
        RECT 30.920 1635.070 31.180 1635.390 ;
        RECT 393.400 1635.245 393.660 1635.390 ;
        RECT 393.390 1634.875 393.670 1635.245 ;
      LAYER via2 ;
        RECT 15.270 2261.880 15.550 2262.160 ;
        RECT 393.390 1634.920 393.670 1635.200 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.245 2262.170 15.575 2262.185 ;
        RECT -4.800 2261.870 15.575 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.245 2261.855 15.575 2261.870 ;
        RECT 393.365 1635.210 393.695 1635.225 ;
        RECT 410.000 1635.210 414.000 1635.360 ;
        RECT 393.365 1634.910 414.000 1635.210 ;
        RECT 393.365 1634.895 393.695 1634.910 ;
        RECT 410.000 1634.760 414.000 1634.910 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1973.600 16.030 1973.660 ;
        RECT 106.790 1973.600 107.110 1973.660 ;
        RECT 15.710 1973.460 107.110 1973.600 ;
        RECT 15.710 1973.400 16.030 1973.460 ;
        RECT 106.790 1973.400 107.110 1973.460 ;
        RECT 106.790 1524.800 107.110 1524.860 ;
        RECT 393.370 1524.800 393.690 1524.860 ;
        RECT 106.790 1524.660 393.690 1524.800 ;
        RECT 106.790 1524.600 107.110 1524.660 ;
        RECT 393.370 1524.600 393.690 1524.660 ;
      LAYER via ;
        RECT 15.740 1973.400 16.000 1973.660 ;
        RECT 106.820 1973.400 107.080 1973.660 ;
        RECT 106.820 1524.600 107.080 1524.860 ;
        RECT 393.400 1524.600 393.660 1524.860 ;
      LAYER met2 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
        RECT 15.800 1973.690 15.940 1974.875 ;
        RECT 15.740 1973.370 16.000 1973.690 ;
        RECT 106.820 1973.370 107.080 1973.690 ;
        RECT 106.880 1524.890 107.020 1973.370 ;
        RECT 106.820 1524.570 107.080 1524.890 ;
        RECT 393.400 1524.570 393.660 1524.890 ;
        RECT 393.460 1521.005 393.600 1524.570 ;
        RECT 393.390 1520.635 393.670 1521.005 ;
      LAYER via2 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
        RECT 393.390 1520.680 393.670 1520.960 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
        RECT 393.365 1520.970 393.695 1520.985 ;
        RECT 410.000 1520.970 414.000 1521.120 ;
        RECT 393.365 1520.670 414.000 1520.970 ;
        RECT 393.365 1520.655 393.695 1520.670 ;
        RECT 410.000 1520.520 414.000 1520.670 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2013.030 558.860 2013.350 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2013.030 558.720 2899.310 558.860 ;
        RECT 2013.030 558.660 2013.350 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2013.060 558.660 2013.320 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2013.050 741.355 2013.330 741.725 ;
        RECT 2013.120 558.950 2013.260 741.355 ;
        RECT 2013.060 558.630 2013.320 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2013.050 741.400 2013.330 741.680 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 1997.465 741.690 2001.465 741.840 ;
        RECT 2013.025 741.690 2013.355 741.705 ;
        RECT 1997.465 741.390 2013.355 741.690 ;
        RECT 1997.465 741.240 2001.465 741.390 ;
        RECT 2013.025 741.375 2013.355 741.390 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 1683.920 15.570 1683.980 ;
        RECT 189.590 1683.920 189.910 1683.980 ;
        RECT 15.250 1683.780 189.910 1683.920 ;
        RECT 15.250 1683.720 15.570 1683.780 ;
        RECT 189.590 1683.720 189.910 1683.780 ;
        RECT 189.590 1407.500 189.910 1407.560 ;
        RECT 393.370 1407.500 393.690 1407.560 ;
        RECT 189.590 1407.360 393.690 1407.500 ;
        RECT 189.590 1407.300 189.910 1407.360 ;
        RECT 393.370 1407.300 393.690 1407.360 ;
      LAYER via ;
        RECT 15.280 1683.720 15.540 1683.980 ;
        RECT 189.620 1683.720 189.880 1683.980 ;
        RECT 189.620 1407.300 189.880 1407.560 ;
        RECT 393.400 1407.300 393.660 1407.560 ;
      LAYER met2 ;
        RECT 15.270 1687.235 15.550 1687.605 ;
        RECT 15.340 1684.010 15.480 1687.235 ;
        RECT 15.280 1683.690 15.540 1684.010 ;
        RECT 189.620 1683.690 189.880 1684.010 ;
        RECT 189.680 1407.590 189.820 1683.690 ;
        RECT 189.620 1407.270 189.880 1407.590 ;
        RECT 393.400 1407.270 393.660 1407.590 ;
        RECT 393.460 1406.765 393.600 1407.270 ;
        RECT 393.390 1406.395 393.670 1406.765 ;
      LAYER via2 ;
        RECT 15.270 1687.280 15.550 1687.560 ;
        RECT 393.390 1406.440 393.670 1406.720 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 15.245 1687.570 15.575 1687.585 ;
        RECT -4.800 1687.270 15.575 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 15.245 1687.255 15.575 1687.270 ;
        RECT 393.365 1406.730 393.695 1406.745 ;
        RECT 410.000 1406.730 414.000 1406.880 ;
        RECT 393.365 1406.430 414.000 1406.730 ;
        RECT 393.365 1406.415 393.695 1406.430 ;
        RECT 410.000 1406.280 414.000 1406.430 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1297.000 17.410 1297.060 ;
        RECT 393.370 1297.000 393.690 1297.060 ;
        RECT 17.090 1296.860 393.690 1297.000 ;
        RECT 17.090 1296.800 17.410 1296.860 ;
        RECT 393.370 1296.800 393.690 1296.860 ;
      LAYER via ;
        RECT 17.120 1296.800 17.380 1297.060 ;
        RECT 393.400 1296.800 393.660 1297.060 ;
      LAYER met2 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
        RECT 17.180 1297.090 17.320 1471.675 ;
        RECT 17.120 1296.770 17.380 1297.090 ;
        RECT 393.400 1296.770 393.660 1297.090 ;
        RECT 393.460 1291.845 393.600 1296.770 ;
        RECT 393.390 1291.475 393.670 1291.845 ;
      LAYER via2 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
        RECT 393.390 1291.520 393.670 1291.800 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
        RECT 393.365 1291.810 393.695 1291.825 ;
        RECT 410.000 1291.810 414.000 1291.960 ;
        RECT 393.365 1291.510 414.000 1291.810 ;
        RECT 393.365 1291.495 393.695 1291.510 ;
        RECT 410.000 1291.360 414.000 1291.510 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1179.700 17.410 1179.760 ;
        RECT 393.370 1179.700 393.690 1179.760 ;
        RECT 17.090 1179.560 393.690 1179.700 ;
        RECT 17.090 1179.500 17.410 1179.560 ;
        RECT 393.370 1179.500 393.690 1179.560 ;
      LAYER via ;
        RECT 17.120 1179.500 17.380 1179.760 ;
        RECT 393.400 1179.500 393.660 1179.760 ;
      LAYER met2 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
        RECT 17.180 1179.790 17.320 1256.115 ;
        RECT 17.120 1179.470 17.380 1179.790 ;
        RECT 393.400 1179.470 393.660 1179.790 ;
        RECT 393.460 1177.605 393.600 1179.470 ;
        RECT 393.390 1177.235 393.670 1177.605 ;
      LAYER via2 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
        RECT 393.390 1177.280 393.670 1177.560 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
        RECT 393.365 1177.570 393.695 1177.585 ;
        RECT 410.000 1177.570 414.000 1177.720 ;
        RECT 393.365 1177.270 414.000 1177.570 ;
        RECT 393.365 1177.255 393.695 1177.270 ;
        RECT 410.000 1177.120 414.000 1177.270 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 396.590 1041.660 396.910 1041.720 ;
        RECT 17.090 1041.520 396.910 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 396.590 1041.460 396.910 1041.520 ;
      LAYER via ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 396.620 1041.460 396.880 1041.720 ;
      LAYER met2 ;
        RECT 396.610 1062.995 396.890 1063.365 ;
        RECT 396.680 1041.750 396.820 1062.995 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 396.620 1041.430 396.880 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 396.610 1063.040 396.890 1063.320 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 396.585 1063.330 396.915 1063.345 ;
        RECT 410.000 1063.330 414.000 1063.480 ;
        RECT 396.585 1063.030 414.000 1063.330 ;
        RECT 396.585 1063.015 396.915 1063.030 ;
        RECT 410.000 1062.880 414.000 1063.030 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 396.590 827.800 396.910 827.860 ;
        RECT 17.550 827.660 396.910 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 396.590 827.600 396.910 827.660 ;
      LAYER via ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 396.620 827.600 396.880 827.860 ;
      LAYER met2 ;
        RECT 396.610 948.755 396.890 949.125 ;
        RECT 396.680 827.890 396.820 948.755 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 396.620 827.570 396.880 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 396.610 948.800 396.890 949.080 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT 396.585 949.090 396.915 949.105 ;
        RECT 410.000 949.090 414.000 949.240 ;
        RECT 396.585 948.790 414.000 949.090 ;
        RECT 396.585 948.775 396.915 948.790 ;
        RECT 410.000 948.640 414.000 948.790 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.790 828.140 107.110 828.200 ;
        RECT 393.370 828.140 393.690 828.200 ;
        RECT 106.790 828.000 393.690 828.140 ;
        RECT 106.790 827.940 107.110 828.000 ;
        RECT 393.370 827.940 393.690 828.000 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 106.790 613.940 107.110 614.000 ;
        RECT 17.090 613.800 107.110 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 106.790 613.740 107.110 613.800 ;
      LAYER via ;
        RECT 106.820 827.940 107.080 828.200 ;
        RECT 393.400 827.940 393.660 828.200 ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 106.820 613.740 107.080 614.000 ;
      LAYER met2 ;
        RECT 393.390 833.835 393.670 834.205 ;
        RECT 393.460 828.230 393.600 833.835 ;
        RECT 106.820 827.910 107.080 828.230 ;
        RECT 393.400 827.910 393.660 828.230 ;
        RECT 106.880 614.030 107.020 827.910 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 106.820 613.710 107.080 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 393.390 833.880 393.670 834.160 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 393.365 834.170 393.695 834.185 ;
        RECT 410.000 834.170 414.000 834.320 ;
        RECT 393.365 833.870 414.000 834.170 ;
        RECT 393.365 833.855 393.695 833.870 ;
        RECT 410.000 833.720 414.000 833.870 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 717.980 45.010 718.040 ;
        RECT 393.370 717.980 393.690 718.040 ;
        RECT 44.690 717.840 393.690 717.980 ;
        RECT 44.690 717.780 45.010 717.840 ;
        RECT 393.370 717.780 393.690 717.840 ;
        RECT 17.550 397.360 17.870 397.420 ;
        RECT 44.690 397.360 45.010 397.420 ;
        RECT 17.550 397.220 45.010 397.360 ;
        RECT 17.550 397.160 17.870 397.220 ;
        RECT 44.690 397.160 45.010 397.220 ;
      LAYER via ;
        RECT 44.720 717.780 44.980 718.040 ;
        RECT 393.400 717.780 393.660 718.040 ;
        RECT 17.580 397.160 17.840 397.420 ;
        RECT 44.720 397.160 44.980 397.420 ;
      LAYER met2 ;
        RECT 393.390 719.595 393.670 719.965 ;
        RECT 393.460 718.070 393.600 719.595 ;
        RECT 44.720 717.750 44.980 718.070 ;
        RECT 393.400 717.750 393.660 718.070 ;
        RECT 44.780 397.450 44.920 717.750 ;
        RECT 17.580 397.130 17.840 397.450 ;
        RECT 44.720 397.130 44.980 397.450 ;
        RECT 17.640 394.925 17.780 397.130 ;
        RECT 17.570 394.555 17.850 394.925 ;
      LAYER via2 ;
        RECT 393.390 719.640 393.670 719.920 ;
        RECT 17.570 394.600 17.850 394.880 ;
      LAYER met3 ;
        RECT 393.365 719.930 393.695 719.945 ;
        RECT 410.000 719.930 414.000 720.080 ;
        RECT 393.365 719.630 414.000 719.930 ;
        RECT 393.365 719.615 393.695 719.630 ;
        RECT 410.000 719.480 414.000 719.630 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.545 394.890 17.875 394.905 ;
        RECT -4.800 394.590 17.875 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.545 394.575 17.875 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.790 600.680 107.110 600.740 ;
        RECT 393.370 600.680 393.690 600.740 ;
        RECT 106.790 600.540 393.690 600.680 ;
        RECT 106.790 600.480 107.110 600.540 ;
        RECT 393.370 600.480 393.690 600.540 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 106.790 179.420 107.110 179.480 ;
        RECT 17.090 179.280 107.110 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 106.790 179.220 107.110 179.280 ;
      LAYER via ;
        RECT 106.820 600.480 107.080 600.740 ;
        RECT 393.400 600.480 393.660 600.740 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 106.820 179.220 107.080 179.480 ;
      LAYER met2 ;
        RECT 393.390 605.355 393.670 605.725 ;
        RECT 393.460 600.770 393.600 605.355 ;
        RECT 106.820 600.450 107.080 600.770 ;
        RECT 393.400 600.450 393.660 600.770 ;
        RECT 106.880 179.510 107.020 600.450 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 106.820 179.190 107.080 179.510 ;
      LAYER via2 ;
        RECT 393.390 605.400 393.670 605.680 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 393.365 605.690 393.695 605.705 ;
        RECT 410.000 605.690 414.000 605.840 ;
        RECT 393.365 605.390 414.000 605.690 ;
        RECT 393.365 605.375 393.695 605.390 ;
        RECT 410.000 605.240 414.000 605.390 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2011.190 793.460 2011.510 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2011.190 793.320 2899.310 793.460 ;
        RECT 2011.190 793.260 2011.510 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2011.220 793.260 2011.480 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2011.210 848.115 2011.490 848.485 ;
        RECT 2011.280 793.550 2011.420 848.115 ;
        RECT 2011.220 793.230 2011.480 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2011.210 848.160 2011.490 848.440 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 1997.465 848.450 2001.465 848.600 ;
        RECT 2011.185 848.450 2011.515 848.465 ;
        RECT 1997.465 848.150 2011.515 848.450 ;
        RECT 1997.465 848.000 2001.465 848.150 ;
        RECT 2011.185 848.135 2011.515 848.150 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.970 959.040 2008.290 959.100 ;
        RECT 2901.750 959.040 2902.070 959.100 ;
        RECT 2007.970 958.900 2902.070 959.040 ;
        RECT 2007.970 958.840 2008.290 958.900 ;
        RECT 2901.750 958.840 2902.070 958.900 ;
      LAYER via ;
        RECT 2008.000 958.840 2008.260 959.100 ;
        RECT 2901.780 958.840 2902.040 959.100 ;
      LAYER met2 ;
        RECT 2901.770 1026.275 2902.050 1026.645 ;
        RECT 2901.840 959.130 2901.980 1026.275 ;
        RECT 2008.000 958.810 2008.260 959.130 ;
        RECT 2901.780 958.810 2902.040 959.130 ;
        RECT 2008.060 955.245 2008.200 958.810 ;
        RECT 2007.990 954.875 2008.270 955.245 ;
      LAYER via2 ;
        RECT 2901.770 1026.320 2902.050 1026.600 ;
        RECT 2007.990 954.920 2008.270 955.200 ;
      LAYER met3 ;
        RECT 2901.745 1026.610 2902.075 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2901.745 1026.310 2924.800 1026.610 ;
        RECT 2901.745 1026.295 2902.075 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 1997.465 955.210 2001.465 955.360 ;
        RECT 2007.965 955.210 2008.295 955.225 ;
        RECT 1997.465 954.910 2008.295 955.210 ;
        RECT 1997.465 954.760 2001.465 954.910 ;
        RECT 2007.965 954.895 2008.295 954.910 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.090 1256.200 2018.410 1256.260 ;
        RECT 2900.830 1256.200 2901.150 1256.260 ;
        RECT 2018.090 1256.060 2901.150 1256.200 ;
        RECT 2018.090 1256.000 2018.410 1256.060 ;
        RECT 2900.830 1256.000 2901.150 1256.060 ;
        RECT 2007.970 1062.060 2008.290 1062.120 ;
        RECT 2018.090 1062.060 2018.410 1062.120 ;
        RECT 2007.970 1061.920 2018.410 1062.060 ;
        RECT 2007.970 1061.860 2008.290 1061.920 ;
        RECT 2018.090 1061.860 2018.410 1061.920 ;
      LAYER via ;
        RECT 2018.120 1256.000 2018.380 1256.260 ;
        RECT 2900.860 1256.000 2901.120 1256.260 ;
        RECT 2008.000 1061.860 2008.260 1062.120 ;
        RECT 2018.120 1061.860 2018.380 1062.120 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 1256.290 2901.060 1260.875 ;
        RECT 2018.120 1255.970 2018.380 1256.290 ;
        RECT 2900.860 1255.970 2901.120 1256.290 ;
        RECT 2018.180 1062.150 2018.320 1255.970 ;
        RECT 2008.000 1062.005 2008.260 1062.150 ;
        RECT 2007.990 1061.635 2008.270 1062.005 ;
        RECT 2018.120 1061.830 2018.380 1062.150 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2007.990 1061.680 2008.270 1061.960 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 1997.465 1061.970 2001.465 1062.120 ;
        RECT 2007.965 1061.970 2008.295 1061.985 ;
        RECT 1997.465 1061.670 2008.295 1061.970 ;
        RECT 1997.465 1061.520 2001.465 1061.670 ;
        RECT 2007.965 1061.655 2008.295 1061.670 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.970 1172.900 2008.290 1172.960 ;
        RECT 2894.390 1172.900 2894.710 1172.960 ;
        RECT 2007.970 1172.760 2894.710 1172.900 ;
        RECT 2007.970 1172.700 2008.290 1172.760 ;
        RECT 2894.390 1172.700 2894.710 1172.760 ;
      LAYER via ;
        RECT 2008.000 1172.700 2008.260 1172.960 ;
        RECT 2894.420 1172.700 2894.680 1172.960 ;
      LAYER met2 ;
        RECT 2894.410 1495.475 2894.690 1495.845 ;
        RECT 2894.480 1172.990 2894.620 1495.475 ;
        RECT 2008.000 1172.670 2008.260 1172.990 ;
        RECT 2894.420 1172.670 2894.680 1172.990 ;
        RECT 2008.060 1168.765 2008.200 1172.670 ;
        RECT 2007.990 1168.395 2008.270 1168.765 ;
      LAYER via2 ;
        RECT 2894.410 1495.520 2894.690 1495.800 ;
        RECT 2007.990 1168.440 2008.270 1168.720 ;
      LAYER met3 ;
        RECT 2894.385 1495.810 2894.715 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2894.385 1495.510 2924.800 1495.810 ;
        RECT 2894.385 1495.495 2894.715 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 1997.465 1168.730 2001.465 1168.880 ;
        RECT 2007.965 1168.730 2008.295 1168.745 ;
        RECT 1997.465 1168.430 2008.295 1168.730 ;
        RECT 1997.465 1168.280 2001.465 1168.430 ;
        RECT 2007.965 1168.415 2008.295 1168.430 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.090 1725.400 2018.410 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 2018.090 1725.260 2901.150 1725.400 ;
        RECT 2018.090 1725.200 2018.410 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
        RECT 2007.970 1275.580 2008.290 1275.640 ;
        RECT 2018.090 1275.580 2018.410 1275.640 ;
        RECT 2007.970 1275.440 2018.410 1275.580 ;
        RECT 2007.970 1275.380 2008.290 1275.440 ;
        RECT 2018.090 1275.380 2018.410 1275.440 ;
      LAYER via ;
        RECT 2018.120 1725.200 2018.380 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
        RECT 2008.000 1275.380 2008.260 1275.640 ;
        RECT 2018.120 1275.380 2018.380 1275.640 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 2018.120 1725.170 2018.380 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 2018.180 1275.670 2018.320 1725.170 ;
        RECT 2008.000 1275.525 2008.260 1275.670 ;
        RECT 2007.990 1275.155 2008.270 1275.525 ;
        RECT 2018.120 1275.350 2018.380 1275.670 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2007.990 1275.200 2008.270 1275.480 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 1997.465 1275.490 2001.465 1275.640 ;
        RECT 2007.965 1275.490 2008.295 1275.505 ;
        RECT 1997.465 1275.190 2008.295 1275.490 ;
        RECT 1997.465 1275.040 2001.465 1275.190 ;
        RECT 2007.965 1275.175 2008.295 1275.190 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2038.790 1960.000 2039.110 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2038.790 1959.860 2901.150 1960.000 ;
        RECT 2038.790 1959.800 2039.110 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
        RECT 2007.970 1386.760 2008.290 1386.820 ;
        RECT 2038.790 1386.760 2039.110 1386.820 ;
        RECT 2007.970 1386.620 2039.110 1386.760 ;
        RECT 2007.970 1386.560 2008.290 1386.620 ;
        RECT 2038.790 1386.560 2039.110 1386.620 ;
      LAYER via ;
        RECT 2038.820 1959.800 2039.080 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
        RECT 2008.000 1386.560 2008.260 1386.820 ;
        RECT 2038.820 1386.560 2039.080 1386.820 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2038.820 1959.770 2039.080 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2038.880 1386.850 2039.020 1959.770 ;
        RECT 2008.000 1386.530 2008.260 1386.850 ;
        RECT 2038.820 1386.530 2039.080 1386.850 ;
        RECT 2008.060 1382.285 2008.200 1386.530 ;
        RECT 2007.990 1381.915 2008.270 1382.285 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2007.990 1381.960 2008.270 1382.240 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 1997.465 1382.250 2001.465 1382.400 ;
        RECT 2007.965 1382.250 2008.295 1382.265 ;
        RECT 1997.465 1381.950 2008.295 1382.250 ;
        RECT 1997.465 1381.800 2001.465 1381.950 ;
        RECT 2007.965 1381.935 2008.295 1381.950 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2804.690 2194.600 2805.010 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2804.690 2194.460 2901.150 2194.600 ;
        RECT 2804.690 2194.400 2805.010 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 2007.970 1490.460 2008.290 1490.520 ;
        RECT 2804.690 1490.460 2805.010 1490.520 ;
        RECT 2007.970 1490.320 2805.010 1490.460 ;
        RECT 2007.970 1490.260 2008.290 1490.320 ;
        RECT 2804.690 1490.260 2805.010 1490.320 ;
      LAYER via ;
        RECT 2804.720 2194.400 2804.980 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 2008.000 1490.260 2008.260 1490.520 ;
        RECT 2804.720 1490.260 2804.980 1490.520 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2804.720 2194.370 2804.980 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2804.780 1490.550 2804.920 2194.370 ;
        RECT 2008.000 1490.230 2008.260 1490.550 ;
        RECT 2804.720 1490.230 2804.980 1490.550 ;
        RECT 2008.060 1489.045 2008.200 1490.230 ;
        RECT 2007.990 1488.675 2008.270 1489.045 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2007.990 1488.720 2008.270 1489.000 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 1997.465 1489.010 2001.465 1489.160 ;
        RECT 2007.965 1489.010 2008.295 1489.025 ;
        RECT 1997.465 1488.710 2008.295 1489.010 ;
        RECT 1997.465 1488.560 2001.465 1488.710 ;
        RECT 2007.965 1488.695 2008.295 1488.710 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.650 206.960 2011.970 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2011.650 206.820 2901.150 206.960 ;
        RECT 2011.650 206.760 2011.970 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2011.680 206.760 2011.940 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2011.670 598.555 2011.950 598.925 ;
        RECT 2011.740 207.050 2011.880 598.555 ;
        RECT 2011.680 206.730 2011.940 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2011.670 598.600 2011.950 598.880 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 1997.465 598.890 2001.465 599.040 ;
        RECT 2011.645 598.890 2011.975 598.905 ;
        RECT 1997.465 598.590 2011.975 598.890 ;
        RECT 1997.465 598.440 2001.465 598.590 ;
        RECT 2011.645 598.575 2011.975 598.590 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2756.390 2546.500 2756.710 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2756.390 2546.360 2901.150 2546.500 ;
        RECT 2756.390 2546.300 2756.710 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
        RECT 2007.970 1669.640 2008.290 1669.700 ;
        RECT 2756.390 1669.640 2756.710 1669.700 ;
        RECT 2007.970 1669.500 2756.710 1669.640 ;
        RECT 2007.970 1669.440 2008.290 1669.500 ;
        RECT 2756.390 1669.440 2756.710 1669.500 ;
      LAYER via ;
        RECT 2756.420 2546.300 2756.680 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
        RECT 2008.000 1669.440 2008.260 1669.700 ;
        RECT 2756.420 1669.440 2756.680 1669.700 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2756.420 2546.270 2756.680 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2756.480 1669.730 2756.620 2546.270 ;
        RECT 2008.000 1669.410 2008.260 1669.730 ;
        RECT 2756.420 1669.410 2756.680 1669.730 ;
        RECT 2008.060 1667.205 2008.200 1669.410 ;
        RECT 2007.990 1666.835 2008.270 1667.205 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2007.990 1666.880 2008.270 1667.160 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 1997.465 1667.170 2001.465 1667.320 ;
        RECT 2007.965 1667.170 2008.295 1667.185 ;
        RECT 1997.465 1666.870 2008.295 1667.170 ;
        RECT 1997.465 1666.720 2001.465 1666.870 ;
        RECT 2007.965 1666.855 2008.295 1666.870 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2818.490 2781.100 2818.810 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2818.490 2780.960 2901.150 2781.100 ;
        RECT 2818.490 2780.900 2818.810 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2007.970 1780.140 2008.290 1780.200 ;
        RECT 2818.490 1780.140 2818.810 1780.200 ;
        RECT 2007.970 1780.000 2818.810 1780.140 ;
        RECT 2007.970 1779.940 2008.290 1780.000 ;
        RECT 2818.490 1779.940 2818.810 1780.000 ;
      LAYER via ;
        RECT 2818.520 2780.900 2818.780 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2008.000 1779.940 2008.260 1780.200 ;
        RECT 2818.520 1779.940 2818.780 1780.200 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2818.520 2780.870 2818.780 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2818.580 1780.230 2818.720 2780.870 ;
        RECT 2008.000 1779.910 2008.260 1780.230 ;
        RECT 2818.520 1779.910 2818.780 1780.230 ;
        RECT 2008.060 1773.965 2008.200 1779.910 ;
        RECT 2007.990 1773.595 2008.270 1773.965 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2007.990 1773.640 2008.270 1773.920 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 1997.465 1773.930 2001.465 1774.080 ;
        RECT 2007.965 1773.930 2008.295 1773.945 ;
        RECT 1997.465 1773.630 2008.295 1773.930 ;
        RECT 1997.465 1773.480 2001.465 1773.630 ;
        RECT 2007.965 1773.615 2008.295 1773.630 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2825.390 3015.700 2825.710 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2825.390 3015.560 2901.150 3015.700 ;
        RECT 2825.390 3015.500 2825.710 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2007.970 1883.500 2008.290 1883.560 ;
        RECT 2825.390 1883.500 2825.710 1883.560 ;
        RECT 2007.970 1883.360 2825.710 1883.500 ;
        RECT 2007.970 1883.300 2008.290 1883.360 ;
        RECT 2825.390 1883.300 2825.710 1883.360 ;
      LAYER via ;
        RECT 2825.420 3015.500 2825.680 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2008.000 1883.300 2008.260 1883.560 ;
        RECT 2825.420 1883.300 2825.680 1883.560 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2825.420 3015.470 2825.680 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2825.480 1883.590 2825.620 3015.470 ;
        RECT 2008.000 1883.270 2008.260 1883.590 ;
        RECT 2825.420 1883.270 2825.680 1883.590 ;
        RECT 2008.060 1880.725 2008.200 1883.270 ;
        RECT 2007.990 1880.355 2008.270 1880.725 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2007.990 1880.400 2008.270 1880.680 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 1997.465 1880.690 2001.465 1880.840 ;
        RECT 2007.965 1880.690 2008.295 1880.705 ;
        RECT 1997.465 1880.390 2008.295 1880.690 ;
        RECT 1997.465 1880.240 2001.465 1880.390 ;
        RECT 2007.965 1880.375 2008.295 1880.390 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2832.290 3250.300 2832.610 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2832.290 3250.160 2901.150 3250.300 ;
        RECT 2832.290 3250.100 2832.610 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2007.970 1994.000 2008.290 1994.060 ;
        RECT 2832.290 1994.000 2832.610 1994.060 ;
        RECT 2007.970 1993.860 2832.610 1994.000 ;
        RECT 2007.970 1993.800 2008.290 1993.860 ;
        RECT 2832.290 1993.800 2832.610 1993.860 ;
      LAYER via ;
        RECT 2832.320 3250.100 2832.580 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2008.000 1993.800 2008.260 1994.060 ;
        RECT 2832.320 1993.800 2832.580 1994.060 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2832.320 3250.070 2832.580 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2832.380 1994.090 2832.520 3250.070 ;
        RECT 2008.000 1993.770 2008.260 1994.090 ;
        RECT 2832.320 1993.770 2832.580 1994.090 ;
        RECT 2008.060 1987.485 2008.200 1993.770 ;
        RECT 2007.990 1987.115 2008.270 1987.485 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2007.990 1987.160 2008.270 1987.440 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 1997.465 1987.450 2001.465 1987.600 ;
        RECT 2007.965 1987.450 2008.295 1987.465 ;
        RECT 1997.465 1987.150 2008.295 1987.450 ;
        RECT 1997.465 1987.000 2001.465 1987.150 ;
        RECT 2007.965 1987.135 2008.295 1987.150 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2839.190 3484.900 2839.510 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2839.190 3484.760 2901.150 3484.900 ;
        RECT 2839.190 3484.700 2839.510 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2007.970 2097.360 2008.290 2097.420 ;
        RECT 2839.190 2097.360 2839.510 2097.420 ;
        RECT 2007.970 2097.220 2839.510 2097.360 ;
        RECT 2007.970 2097.160 2008.290 2097.220 ;
        RECT 2839.190 2097.160 2839.510 2097.220 ;
      LAYER via ;
        RECT 2839.220 3484.700 2839.480 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2008.000 2097.160 2008.260 2097.420 ;
        RECT 2839.220 2097.160 2839.480 2097.420 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2839.220 3484.670 2839.480 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2839.280 2097.450 2839.420 3484.670 ;
        RECT 2008.000 2097.130 2008.260 2097.450 ;
        RECT 2839.220 2097.130 2839.480 2097.450 ;
        RECT 2008.060 2094.245 2008.200 2097.130 ;
        RECT 2007.990 2093.875 2008.270 2094.245 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2007.990 2093.920 2008.270 2094.200 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 1997.465 2094.210 2001.465 2094.360 ;
        RECT 2007.965 2094.210 2008.295 2094.225 ;
        RECT 1997.465 2093.910 2008.295 2094.210 ;
        RECT 1997.465 2093.760 2001.465 2093.910 ;
        RECT 2007.965 2093.895 2008.295 2093.910 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1853.870 2122.520 1854.190 2122.580 ;
        RECT 2635.870 2122.520 2636.190 2122.580 ;
        RECT 1853.870 2122.380 2636.190 2122.520 ;
        RECT 1853.870 2122.320 1854.190 2122.380 ;
        RECT 2635.870 2122.320 2636.190 2122.380 ;
      LAYER via ;
        RECT 1853.900 2122.320 1854.160 2122.580 ;
        RECT 2635.900 2122.320 2636.160 2122.580 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 2122.610 2636.100 3517.600 ;
        RECT 1853.900 2122.290 1854.160 2122.610 ;
        RECT 2635.900 2122.290 2636.160 2122.610 ;
        RECT 1853.960 2112.185 1854.100 2122.290 ;
        RECT 1853.960 2111.740 1854.310 2112.185 ;
        RECT 1854.030 2108.185 1854.310 2111.740 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1677.230 2123.540 1677.550 2123.600 ;
        RECT 2311.570 2123.540 2311.890 2123.600 ;
        RECT 1677.230 2123.400 2311.890 2123.540 ;
        RECT 1677.230 2123.340 1677.550 2123.400 ;
        RECT 2311.570 2123.340 2311.890 2123.400 ;
      LAYER via ;
        RECT 1677.260 2123.340 1677.520 2123.600 ;
        RECT 2311.600 2123.340 2311.860 2123.600 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 2123.630 2311.800 3517.600 ;
        RECT 1677.260 2123.310 1677.520 2123.630 ;
        RECT 2311.600 2123.310 2311.860 2123.630 ;
        RECT 1677.320 2112.185 1677.460 2123.310 ;
        RECT 1677.320 2111.740 1677.670 2112.185 ;
        RECT 1677.390 2108.185 1677.670 2111.740 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1500.130 2124.560 1500.450 2124.620 ;
        RECT 1987.270 2124.560 1987.590 2124.620 ;
        RECT 1500.130 2124.420 1987.590 2124.560 ;
        RECT 1500.130 2124.360 1500.450 2124.420 ;
        RECT 1987.270 2124.360 1987.590 2124.420 ;
      LAYER via ;
        RECT 1500.160 2124.360 1500.420 2124.620 ;
        RECT 1987.300 2124.360 1987.560 2124.620 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 2124.650 1987.500 3517.600 ;
        RECT 1500.160 2124.330 1500.420 2124.650 ;
        RECT 1987.300 2124.330 1987.560 2124.650 ;
        RECT 1500.220 2112.185 1500.360 2124.330 ;
        RECT 1500.220 2111.740 1500.570 2112.185 ;
        RECT 1500.290 2108.185 1500.570 2111.740 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.070 3487.960 1656.390 3488.020 ;
        RECT 1662.510 3487.960 1662.830 3488.020 ;
        RECT 1656.070 3487.820 1662.830 3487.960 ;
        RECT 1656.070 3487.760 1656.390 3487.820 ;
        RECT 1662.510 3487.760 1662.830 3487.820 ;
        RECT 1323.490 2122.520 1323.810 2122.580 ;
        RECT 1656.070 2122.520 1656.390 2122.580 ;
        RECT 1323.490 2122.380 1656.390 2122.520 ;
        RECT 1323.490 2122.320 1323.810 2122.380 ;
        RECT 1656.070 2122.320 1656.390 2122.380 ;
      LAYER via ;
        RECT 1656.100 3487.760 1656.360 3488.020 ;
        RECT 1662.540 3487.760 1662.800 3488.020 ;
        RECT 1323.520 2122.320 1323.780 2122.580 ;
        RECT 1656.100 2122.320 1656.360 2122.580 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3488.050 1662.740 3517.600 ;
        RECT 1656.100 3487.730 1656.360 3488.050 ;
        RECT 1662.540 3487.730 1662.800 3488.050 ;
        RECT 1656.160 2122.610 1656.300 3487.730 ;
        RECT 1323.520 2122.290 1323.780 2122.610 ;
        RECT 1656.100 2122.290 1656.360 2122.610 ;
        RECT 1323.580 2112.185 1323.720 2122.290 ;
        RECT 1323.580 2111.740 1323.930 2112.185 ;
        RECT 1323.650 2108.185 1323.930 2111.740 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.770 3487.960 1332.090 3488.020 ;
        RECT 1338.210 3487.960 1338.530 3488.020 ;
        RECT 1331.770 3487.820 1338.530 3487.960 ;
        RECT 1331.770 3487.760 1332.090 3487.820 ;
        RECT 1338.210 3487.760 1338.530 3487.820 ;
        RECT 1146.390 2122.180 1146.710 2122.240 ;
        RECT 1331.770 2122.180 1332.090 2122.240 ;
        RECT 1146.390 2122.040 1332.090 2122.180 ;
        RECT 1146.390 2121.980 1146.710 2122.040 ;
        RECT 1331.770 2121.980 1332.090 2122.040 ;
      LAYER via ;
        RECT 1331.800 3487.760 1332.060 3488.020 ;
        RECT 1338.240 3487.760 1338.500 3488.020 ;
        RECT 1146.420 2121.980 1146.680 2122.240 ;
        RECT 1331.800 2121.980 1332.060 2122.240 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3488.050 1338.440 3517.600 ;
        RECT 1331.800 3487.730 1332.060 3488.050 ;
        RECT 1338.240 3487.730 1338.500 3488.050 ;
        RECT 1331.860 2122.270 1332.000 3487.730 ;
        RECT 1146.420 2121.950 1146.680 2122.270 ;
        RECT 1331.800 2121.950 1332.060 2122.270 ;
        RECT 1146.480 2112.185 1146.620 2121.950 ;
        RECT 1146.480 2111.740 1146.830 2112.185 ;
        RECT 1146.550 2108.185 1146.830 2111.740 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2012.570 441.560 2012.890 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2012.570 441.420 2901.150 441.560 ;
        RECT 2012.570 441.360 2012.890 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2012.600 441.360 2012.860 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2012.590 705.315 2012.870 705.685 ;
        RECT 2012.660 441.650 2012.800 705.315 ;
        RECT 2012.600 441.330 2012.860 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2012.590 705.360 2012.870 705.640 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 1997.465 705.650 2001.465 705.800 ;
        RECT 2012.565 705.650 2012.895 705.665 ;
        RECT 1997.465 705.350 2012.895 705.650 ;
        RECT 1997.465 705.200 2001.465 705.350 ;
        RECT 2012.565 705.335 2012.895 705.350 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1007.470 3487.960 1007.790 3488.020 ;
        RECT 1013.910 3487.960 1014.230 3488.020 ;
        RECT 1007.470 3487.820 1014.230 3487.960 ;
        RECT 1007.470 3487.760 1007.790 3487.820 ;
        RECT 1013.910 3487.760 1014.230 3487.820 ;
        RECT 969.750 2118.440 970.070 2118.500 ;
        RECT 1007.470 2118.440 1007.790 2118.500 ;
        RECT 969.750 2118.300 1007.790 2118.440 ;
        RECT 969.750 2118.240 970.070 2118.300 ;
        RECT 1007.470 2118.240 1007.790 2118.300 ;
      LAYER via ;
        RECT 1007.500 3487.760 1007.760 3488.020 ;
        RECT 1013.940 3487.760 1014.200 3488.020 ;
        RECT 969.780 2118.240 970.040 2118.500 ;
        RECT 1007.500 2118.240 1007.760 2118.500 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3488.050 1014.140 3517.600 ;
        RECT 1007.500 3487.730 1007.760 3488.050 ;
        RECT 1013.940 3487.730 1014.200 3488.050 ;
        RECT 1007.560 2118.530 1007.700 3487.730 ;
        RECT 969.780 2118.210 970.040 2118.530 ;
        RECT 1007.500 2118.210 1007.760 2118.530 ;
        RECT 969.840 2112.185 969.980 2118.210 ;
        RECT 969.840 2111.740 970.190 2112.185 ;
        RECT 969.910 2108.185 970.190 2111.740 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
        RECT 688.765 2898.585 688.935 2946.355 ;
        RECT 687.845 2849.625 688.015 2898.075 ;
        RECT 688.305 2753.065 688.475 2801.175 ;
        RECT 689.225 2186.965 689.395 2221.815 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
        RECT 688.765 2946.185 688.935 2946.355 ;
        RECT 687.845 2897.905 688.015 2898.075 ;
        RECT 688.305 2801.005 688.475 2801.175 ;
        RECT 689.225 2221.645 689.395 2221.815 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3270.700 689.010 3270.760 ;
        RECT 689.610 3270.700 689.930 3270.760 ;
        RECT 688.690 3270.560 689.930 3270.700 ;
        RECT 688.690 3270.500 689.010 3270.560 ;
        RECT 689.610 3270.500 689.930 3270.560 ;
        RECT 688.690 3174.140 689.010 3174.200 ;
        RECT 689.610 3174.140 689.930 3174.200 ;
        RECT 688.690 3174.000 689.930 3174.140 ;
        RECT 688.690 3173.940 689.010 3174.000 ;
        RECT 689.610 3173.940 689.930 3174.000 ;
        RECT 688.690 3077.580 689.010 3077.640 ;
        RECT 689.610 3077.580 689.930 3077.640 ;
        RECT 688.690 3077.440 689.930 3077.580 ;
        RECT 688.690 3077.380 689.010 3077.440 ;
        RECT 689.610 3077.380 689.930 3077.440 ;
        RECT 688.690 2981.020 689.010 2981.080 ;
        RECT 689.610 2981.020 689.930 2981.080 ;
        RECT 688.690 2980.880 689.930 2981.020 ;
        RECT 688.690 2980.820 689.010 2980.880 ;
        RECT 689.610 2980.820 689.930 2980.880 ;
        RECT 688.690 2946.340 689.010 2946.400 ;
        RECT 688.495 2946.200 689.010 2946.340 ;
        RECT 688.690 2946.140 689.010 2946.200 ;
        RECT 688.690 2898.740 689.010 2898.800 ;
        RECT 688.495 2898.600 689.010 2898.740 ;
        RECT 688.690 2898.540 689.010 2898.600 ;
        RECT 687.785 2898.060 688.075 2898.105 ;
        RECT 688.230 2898.060 688.550 2898.120 ;
        RECT 687.785 2897.920 688.550 2898.060 ;
        RECT 687.785 2897.875 688.075 2897.920 ;
        RECT 688.230 2897.860 688.550 2897.920 ;
        RECT 687.770 2849.780 688.090 2849.840 ;
        RECT 687.575 2849.640 688.090 2849.780 ;
        RECT 687.770 2849.580 688.090 2849.640 ;
        RECT 687.770 2815.240 688.090 2815.500 ;
        RECT 687.860 2814.760 688.000 2815.240 ;
        RECT 688.230 2814.760 688.550 2814.820 ;
        RECT 687.860 2814.620 688.550 2814.760 ;
        RECT 688.230 2814.560 688.550 2814.620 ;
        RECT 688.230 2801.160 688.550 2801.220 ;
        RECT 688.035 2801.020 688.550 2801.160 ;
        RECT 688.230 2800.960 688.550 2801.020 ;
        RECT 688.245 2753.220 688.535 2753.265 ;
        RECT 689.150 2753.220 689.470 2753.280 ;
        RECT 688.245 2753.080 689.470 2753.220 ;
        RECT 688.245 2753.035 688.535 2753.080 ;
        RECT 689.150 2753.020 689.470 2753.080 ;
        RECT 688.230 2718.200 688.550 2718.260 ;
        RECT 689.150 2718.200 689.470 2718.260 ;
        RECT 688.230 2718.060 689.470 2718.200 ;
        RECT 688.230 2718.000 688.550 2718.060 ;
        RECT 689.150 2718.000 689.470 2718.060 ;
        RECT 688.230 2670.260 688.550 2670.320 ;
        RECT 689.150 2670.260 689.470 2670.320 ;
        RECT 688.230 2670.120 689.470 2670.260 ;
        RECT 688.230 2670.060 688.550 2670.120 ;
        RECT 689.150 2670.060 689.470 2670.120 ;
        RECT 689.610 2608.380 689.930 2608.440 ;
        RECT 690.530 2608.380 690.850 2608.440 ;
        RECT 689.610 2608.240 690.850 2608.380 ;
        RECT 689.610 2608.180 689.930 2608.240 ;
        RECT 690.530 2608.180 690.850 2608.240 ;
        RECT 689.610 2511.820 689.930 2511.880 ;
        RECT 690.530 2511.820 690.850 2511.880 ;
        RECT 689.610 2511.680 690.850 2511.820 ;
        RECT 689.610 2511.620 689.930 2511.680 ;
        RECT 690.530 2511.620 690.850 2511.680 ;
        RECT 688.230 2463.200 688.550 2463.260 ;
        RECT 689.150 2463.200 689.470 2463.260 ;
        RECT 688.230 2463.060 689.470 2463.200 ;
        RECT 688.230 2463.000 688.550 2463.060 ;
        RECT 689.150 2463.000 689.470 2463.060 ;
        RECT 687.310 2366.640 687.630 2366.700 ;
        RECT 688.690 2366.640 689.010 2366.700 ;
        RECT 687.310 2366.500 689.010 2366.640 ;
        RECT 687.310 2366.440 687.630 2366.500 ;
        RECT 688.690 2366.440 689.010 2366.500 ;
        RECT 688.690 2235.540 689.010 2235.800 ;
        RECT 688.780 2235.400 688.920 2235.540 ;
        RECT 689.150 2235.400 689.470 2235.460 ;
        RECT 688.780 2235.260 689.470 2235.400 ;
        RECT 689.150 2235.200 689.470 2235.260 ;
        RECT 689.150 2221.800 689.470 2221.860 ;
        RECT 688.955 2221.660 689.470 2221.800 ;
        RECT 689.150 2221.600 689.470 2221.660 ;
        RECT 689.150 2187.120 689.470 2187.180 ;
        RECT 688.955 2186.980 689.470 2187.120 ;
        RECT 689.150 2186.920 689.470 2186.980 ;
        RECT 688.690 2125.580 689.010 2125.640 ;
        RECT 689.610 2125.580 689.930 2125.640 ;
        RECT 688.690 2125.440 689.930 2125.580 ;
        RECT 688.690 2125.380 689.010 2125.440 ;
        RECT 689.610 2125.380 689.930 2125.440 ;
        RECT 688.690 2121.840 689.010 2121.900 ;
        RECT 792.650 2121.840 792.970 2121.900 ;
        RECT 688.690 2121.700 792.970 2121.840 ;
        RECT 688.690 2121.640 689.010 2121.700 ;
        RECT 792.650 2121.640 792.970 2121.700 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3270.500 688.980 3270.760 ;
        RECT 689.640 3270.500 689.900 3270.760 ;
        RECT 688.720 3173.940 688.980 3174.200 ;
        RECT 689.640 3173.940 689.900 3174.200 ;
        RECT 688.720 3077.380 688.980 3077.640 ;
        RECT 689.640 3077.380 689.900 3077.640 ;
        RECT 688.720 2980.820 688.980 2981.080 ;
        RECT 689.640 2980.820 689.900 2981.080 ;
        RECT 688.720 2946.140 688.980 2946.400 ;
        RECT 688.720 2898.540 688.980 2898.800 ;
        RECT 688.260 2897.860 688.520 2898.120 ;
        RECT 687.800 2849.580 688.060 2849.840 ;
        RECT 687.800 2815.240 688.060 2815.500 ;
        RECT 688.260 2814.560 688.520 2814.820 ;
        RECT 688.260 2800.960 688.520 2801.220 ;
        RECT 689.180 2753.020 689.440 2753.280 ;
        RECT 688.260 2718.000 688.520 2718.260 ;
        RECT 689.180 2718.000 689.440 2718.260 ;
        RECT 688.260 2670.060 688.520 2670.320 ;
        RECT 689.180 2670.060 689.440 2670.320 ;
        RECT 689.640 2608.180 689.900 2608.440 ;
        RECT 690.560 2608.180 690.820 2608.440 ;
        RECT 689.640 2511.620 689.900 2511.880 ;
        RECT 690.560 2511.620 690.820 2511.880 ;
        RECT 688.260 2463.000 688.520 2463.260 ;
        RECT 689.180 2463.000 689.440 2463.260 ;
        RECT 687.340 2366.440 687.600 2366.700 ;
        RECT 688.720 2366.440 688.980 2366.700 ;
        RECT 688.720 2235.540 688.980 2235.800 ;
        RECT 689.180 2235.200 689.440 2235.460 ;
        RECT 689.180 2221.600 689.440 2221.860 ;
        RECT 689.180 2186.920 689.440 2187.180 ;
        RECT 688.720 2125.380 688.980 2125.640 ;
        RECT 689.640 2125.380 689.900 2125.640 ;
        RECT 688.720 2121.640 688.980 2121.900 ;
        RECT 792.680 2121.640 792.940 2121.900 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3270.790 688.920 3318.670 ;
        RECT 688.720 3270.470 688.980 3270.790 ;
        RECT 689.640 3270.470 689.900 3270.790 ;
        RECT 689.700 3222.250 689.840 3270.470 ;
        RECT 688.780 3222.110 689.840 3222.250 ;
        RECT 688.780 3174.230 688.920 3222.110 ;
        RECT 688.720 3173.910 688.980 3174.230 ;
        RECT 689.640 3173.910 689.900 3174.230 ;
        RECT 689.700 3125.690 689.840 3173.910 ;
        RECT 688.780 3125.550 689.840 3125.690 ;
        RECT 688.780 3077.670 688.920 3125.550 ;
        RECT 688.720 3077.350 688.980 3077.670 ;
        RECT 689.640 3077.350 689.900 3077.670 ;
        RECT 689.700 3029.130 689.840 3077.350 ;
        RECT 688.780 3028.990 689.840 3029.130 ;
        RECT 688.780 2981.110 688.920 3028.990 ;
        RECT 688.720 2980.790 688.980 2981.110 ;
        RECT 689.640 2980.850 689.900 2981.110 ;
        RECT 689.240 2980.790 689.900 2980.850 ;
        RECT 689.240 2980.710 689.840 2980.790 ;
        RECT 689.240 2959.770 689.380 2980.710 ;
        RECT 688.780 2959.630 689.380 2959.770 ;
        RECT 688.780 2946.430 688.920 2959.630 ;
        RECT 688.720 2946.110 688.980 2946.430 ;
        RECT 688.720 2898.570 688.980 2898.830 ;
        RECT 688.320 2898.510 688.980 2898.570 ;
        RECT 688.320 2898.430 688.920 2898.510 ;
        RECT 688.320 2898.150 688.460 2898.430 ;
        RECT 688.260 2897.830 688.520 2898.150 ;
        RECT 687.800 2849.550 688.060 2849.870 ;
        RECT 687.860 2815.530 688.000 2849.550 ;
        RECT 687.800 2815.210 688.060 2815.530 ;
        RECT 688.260 2814.530 688.520 2814.850 ;
        RECT 688.320 2801.250 688.460 2814.530 ;
        RECT 688.260 2800.930 688.520 2801.250 ;
        RECT 689.180 2752.990 689.440 2753.310 ;
        RECT 689.240 2718.290 689.380 2752.990 ;
        RECT 688.260 2717.970 688.520 2718.290 ;
        RECT 689.180 2717.970 689.440 2718.290 ;
        RECT 688.320 2670.350 688.460 2717.970 ;
        RECT 688.260 2670.030 688.520 2670.350 ;
        RECT 689.180 2670.030 689.440 2670.350 ;
        RECT 689.240 2656.605 689.380 2670.030 ;
        RECT 689.170 2656.235 689.450 2656.605 ;
        RECT 690.550 2656.235 690.830 2656.605 ;
        RECT 690.620 2608.470 690.760 2656.235 ;
        RECT 689.640 2608.150 689.900 2608.470 ;
        RECT 690.560 2608.150 690.820 2608.470 ;
        RECT 689.700 2573.530 689.840 2608.150 ;
        RECT 689.240 2573.390 689.840 2573.530 ;
        RECT 689.240 2560.045 689.380 2573.390 ;
        RECT 689.170 2559.675 689.450 2560.045 ;
        RECT 690.550 2559.675 690.830 2560.045 ;
        RECT 690.620 2511.910 690.760 2559.675 ;
        RECT 689.640 2511.590 689.900 2511.910 ;
        RECT 690.560 2511.590 690.820 2511.910 ;
        RECT 689.700 2476.970 689.840 2511.590 ;
        RECT 689.240 2476.830 689.840 2476.970 ;
        RECT 689.240 2463.290 689.380 2476.830 ;
        RECT 688.260 2462.970 688.520 2463.290 ;
        RECT 689.180 2462.970 689.440 2463.290 ;
        RECT 688.320 2415.205 688.460 2462.970 ;
        RECT 688.250 2414.835 688.530 2415.205 ;
        RECT 689.630 2414.835 689.910 2415.205 ;
        RECT 689.700 2380.410 689.840 2414.835 ;
        RECT 688.780 2380.270 689.840 2380.410 ;
        RECT 688.780 2366.730 688.920 2380.270 ;
        RECT 687.340 2366.410 687.600 2366.730 ;
        RECT 688.720 2366.410 688.980 2366.730 ;
        RECT 687.400 2318.645 687.540 2366.410 ;
        RECT 687.330 2318.275 687.610 2318.645 ;
        RECT 688.250 2318.275 688.530 2318.645 ;
        RECT 688.320 2283.850 688.460 2318.275 ;
        RECT 688.320 2283.710 688.920 2283.850 ;
        RECT 688.780 2235.830 688.920 2283.710 ;
        RECT 688.720 2235.510 688.980 2235.830 ;
        RECT 689.180 2235.170 689.440 2235.490 ;
        RECT 689.240 2221.890 689.380 2235.170 ;
        RECT 689.180 2221.570 689.440 2221.890 ;
        RECT 689.180 2186.890 689.440 2187.210 ;
        RECT 689.240 2173.690 689.380 2186.890 ;
        RECT 689.240 2173.550 689.840 2173.690 ;
        RECT 689.700 2125.670 689.840 2173.550 ;
        RECT 688.720 2125.350 688.980 2125.670 ;
        RECT 689.640 2125.350 689.900 2125.670 ;
        RECT 688.780 2121.930 688.920 2125.350 ;
        RECT 688.720 2121.610 688.980 2121.930 ;
        RECT 792.680 2121.610 792.940 2121.930 ;
        RECT 792.740 2112.185 792.880 2121.610 ;
        RECT 792.740 2111.740 793.090 2112.185 ;
        RECT 792.810 2108.185 793.090 2111.740 ;
      LAYER via2 ;
        RECT 689.170 2656.280 689.450 2656.560 ;
        RECT 690.550 2656.280 690.830 2656.560 ;
        RECT 689.170 2559.720 689.450 2560.000 ;
        RECT 690.550 2559.720 690.830 2560.000 ;
        RECT 688.250 2414.880 688.530 2415.160 ;
        RECT 689.630 2414.880 689.910 2415.160 ;
        RECT 687.330 2318.320 687.610 2318.600 ;
        RECT 688.250 2318.320 688.530 2318.600 ;
      LAYER met3 ;
        RECT 689.145 2656.570 689.475 2656.585 ;
        RECT 690.525 2656.570 690.855 2656.585 ;
        RECT 689.145 2656.270 690.855 2656.570 ;
        RECT 689.145 2656.255 689.475 2656.270 ;
        RECT 690.525 2656.255 690.855 2656.270 ;
        RECT 689.145 2560.010 689.475 2560.025 ;
        RECT 690.525 2560.010 690.855 2560.025 ;
        RECT 689.145 2559.710 690.855 2560.010 ;
        RECT 689.145 2559.695 689.475 2559.710 ;
        RECT 690.525 2559.695 690.855 2559.710 ;
        RECT 688.225 2415.170 688.555 2415.185 ;
        RECT 689.605 2415.170 689.935 2415.185 ;
        RECT 688.225 2414.870 689.935 2415.170 ;
        RECT 688.225 2414.855 688.555 2414.870 ;
        RECT 689.605 2414.855 689.935 2414.870 ;
        RECT 687.305 2318.610 687.635 2318.625 ;
        RECT 688.225 2318.610 688.555 2318.625 ;
        RECT 687.305 2318.310 688.555 2318.610 ;
        RECT 687.305 2318.295 687.635 2318.310 ;
        RECT 688.225 2318.295 688.555 2318.310 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
        RECT 364.925 3236.205 365.095 3284.315 ;
        RECT 365.385 3084.225 365.555 3132.675 ;
        RECT 364.465 2946.525 364.635 2994.635 ;
        RECT 363.085 2849.625 363.255 2898.075 ;
        RECT 363.085 2753.065 363.255 2767.175 ;
        RECT 363.085 2656.505 363.255 2670.615 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
        RECT 364.925 3284.145 365.095 3284.315 ;
        RECT 365.385 3132.505 365.555 3132.675 ;
        RECT 364.465 2994.465 364.635 2994.635 ;
        RECT 363.085 2897.905 363.255 2898.075 ;
        RECT 363.085 2767.005 363.255 2767.175 ;
        RECT 363.085 2670.445 363.255 2670.615 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 364.390 3298.240 364.710 3298.300 ;
        RECT 365.310 3298.240 365.630 3298.300 ;
        RECT 364.390 3298.100 365.630 3298.240 ;
        RECT 364.390 3298.040 364.710 3298.100 ;
        RECT 365.310 3298.040 365.630 3298.100 ;
        RECT 364.865 3284.300 365.155 3284.345 ;
        RECT 365.310 3284.300 365.630 3284.360 ;
        RECT 364.865 3284.160 365.630 3284.300 ;
        RECT 364.865 3284.115 365.155 3284.160 ;
        RECT 365.310 3284.100 365.630 3284.160 ;
        RECT 364.850 3236.360 365.170 3236.420 ;
        RECT 364.655 3236.220 365.170 3236.360 ;
        RECT 364.850 3236.160 365.170 3236.220 ;
        RECT 364.850 3202.020 365.170 3202.080 ;
        RECT 364.020 3201.880 365.170 3202.020 ;
        RECT 364.020 3201.400 364.160 3201.880 ;
        RECT 364.850 3201.820 365.170 3201.880 ;
        RECT 363.930 3201.140 364.250 3201.400 ;
        RECT 363.930 3187.740 364.250 3187.800 ;
        RECT 364.390 3187.740 364.710 3187.800 ;
        RECT 363.930 3187.600 364.710 3187.740 ;
        RECT 363.930 3187.540 364.250 3187.600 ;
        RECT 364.390 3187.540 364.710 3187.600 ;
        RECT 365.310 3132.660 365.630 3132.720 ;
        RECT 365.115 3132.520 365.630 3132.660 ;
        RECT 365.310 3132.460 365.630 3132.520 ;
        RECT 365.310 3084.380 365.630 3084.440 ;
        RECT 365.115 3084.240 365.630 3084.380 ;
        RECT 365.310 3084.180 365.630 3084.240 ;
        RECT 365.310 3057.180 365.630 3057.240 ;
        RECT 364.480 3057.040 365.630 3057.180 ;
        RECT 364.480 3056.560 364.620 3057.040 ;
        RECT 365.310 3056.980 365.630 3057.040 ;
        RECT 364.390 3056.300 364.710 3056.560 ;
        RECT 364.850 3007.880 365.170 3007.940 ;
        RECT 365.770 3007.880 366.090 3007.940 ;
        RECT 364.850 3007.740 366.090 3007.880 ;
        RECT 364.850 3007.680 365.170 3007.740 ;
        RECT 365.770 3007.680 366.090 3007.740 ;
        RECT 364.405 2994.620 364.695 2994.665 ;
        RECT 364.850 2994.620 365.170 2994.680 ;
        RECT 364.405 2994.480 365.170 2994.620 ;
        RECT 364.405 2994.435 364.695 2994.480 ;
        RECT 364.850 2994.420 365.170 2994.480 ;
        RECT 364.390 2946.680 364.710 2946.740 ;
        RECT 364.195 2946.540 364.710 2946.680 ;
        RECT 364.390 2946.480 364.710 2946.540 ;
        RECT 363.470 2912.000 363.790 2912.060 ;
        RECT 364.390 2912.000 364.710 2912.060 ;
        RECT 363.470 2911.860 364.710 2912.000 ;
        RECT 363.470 2911.800 363.790 2911.860 ;
        RECT 364.390 2911.800 364.710 2911.860 ;
        RECT 363.025 2898.060 363.315 2898.105 ;
        RECT 363.470 2898.060 363.790 2898.120 ;
        RECT 363.025 2897.920 363.790 2898.060 ;
        RECT 363.025 2897.875 363.315 2897.920 ;
        RECT 363.470 2897.860 363.790 2897.920 ;
        RECT 363.010 2849.780 363.330 2849.840 ;
        RECT 362.815 2849.640 363.330 2849.780 ;
        RECT 363.010 2849.580 363.330 2849.640 ;
        RECT 363.010 2815.240 363.330 2815.500 ;
        RECT 363.100 2814.760 363.240 2815.240 ;
        RECT 363.470 2814.760 363.790 2814.820 ;
        RECT 363.100 2814.620 363.790 2814.760 ;
        RECT 363.470 2814.560 363.790 2814.620 ;
        RECT 363.010 2767.160 363.330 2767.220 ;
        RECT 362.815 2767.020 363.330 2767.160 ;
        RECT 363.010 2766.960 363.330 2767.020 ;
        RECT 363.010 2753.220 363.330 2753.280 ;
        RECT 362.815 2753.080 363.330 2753.220 ;
        RECT 363.010 2753.020 363.330 2753.080 ;
        RECT 363.010 2718.680 363.330 2718.940 ;
        RECT 363.100 2718.200 363.240 2718.680 ;
        RECT 363.470 2718.200 363.790 2718.260 ;
        RECT 363.100 2718.060 363.790 2718.200 ;
        RECT 363.470 2718.000 363.790 2718.060 ;
        RECT 363.010 2670.600 363.330 2670.660 ;
        RECT 362.815 2670.460 363.330 2670.600 ;
        RECT 363.010 2670.400 363.330 2670.460 ;
        RECT 363.010 2656.660 363.330 2656.720 ;
        RECT 362.815 2656.520 363.330 2656.660 ;
        RECT 363.010 2656.460 363.330 2656.520 ;
        RECT 363.470 2621.640 363.790 2621.700 ;
        RECT 364.390 2621.640 364.710 2621.700 ;
        RECT 363.470 2621.500 364.710 2621.640 ;
        RECT 363.470 2621.440 363.790 2621.500 ;
        RECT 364.390 2621.440 364.710 2621.500 ;
        RECT 363.010 2511.820 363.330 2511.880 ;
        RECT 365.310 2511.820 365.630 2511.880 ;
        RECT 363.010 2511.680 365.630 2511.820 ;
        RECT 363.010 2511.620 363.330 2511.680 ;
        RECT 365.310 2511.620 365.630 2511.680 ;
        RECT 364.390 2401.320 364.710 2401.380 ;
        RECT 365.310 2401.320 365.630 2401.380 ;
        RECT 364.390 2401.180 365.630 2401.320 ;
        RECT 364.390 2401.120 364.710 2401.180 ;
        RECT 365.310 2401.120 365.630 2401.180 ;
        RECT 364.390 2304.760 364.710 2304.820 ;
        RECT 365.310 2304.760 365.630 2304.820 ;
        RECT 364.390 2304.620 365.630 2304.760 ;
        RECT 364.390 2304.560 364.710 2304.620 ;
        RECT 365.310 2304.560 365.630 2304.620 ;
        RECT 363.930 2187.460 364.250 2187.520 ;
        RECT 364.850 2187.460 365.170 2187.520 ;
        RECT 363.930 2187.320 365.170 2187.460 ;
        RECT 363.930 2187.260 364.250 2187.320 ;
        RECT 364.850 2187.260 365.170 2187.320 ;
        RECT 363.930 2122.860 364.250 2122.920 ;
        RECT 616.010 2122.860 616.330 2122.920 ;
        RECT 363.930 2122.720 616.330 2122.860 ;
        RECT 363.930 2122.660 364.250 2122.720 ;
        RECT 616.010 2122.660 616.330 2122.720 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 364.420 3298.040 364.680 3298.300 ;
        RECT 365.340 3298.040 365.600 3298.300 ;
        RECT 365.340 3284.100 365.600 3284.360 ;
        RECT 364.880 3236.160 365.140 3236.420 ;
        RECT 364.880 3201.820 365.140 3202.080 ;
        RECT 363.960 3201.140 364.220 3201.400 ;
        RECT 363.960 3187.540 364.220 3187.800 ;
        RECT 364.420 3187.540 364.680 3187.800 ;
        RECT 365.340 3132.460 365.600 3132.720 ;
        RECT 365.340 3084.180 365.600 3084.440 ;
        RECT 365.340 3056.980 365.600 3057.240 ;
        RECT 364.420 3056.300 364.680 3056.560 ;
        RECT 364.880 3007.680 365.140 3007.940 ;
        RECT 365.800 3007.680 366.060 3007.940 ;
        RECT 364.880 2994.420 365.140 2994.680 ;
        RECT 364.420 2946.480 364.680 2946.740 ;
        RECT 363.500 2911.800 363.760 2912.060 ;
        RECT 364.420 2911.800 364.680 2912.060 ;
        RECT 363.500 2897.860 363.760 2898.120 ;
        RECT 363.040 2849.580 363.300 2849.840 ;
        RECT 363.040 2815.240 363.300 2815.500 ;
        RECT 363.500 2814.560 363.760 2814.820 ;
        RECT 363.040 2766.960 363.300 2767.220 ;
        RECT 363.040 2753.020 363.300 2753.280 ;
        RECT 363.040 2718.680 363.300 2718.940 ;
        RECT 363.500 2718.000 363.760 2718.260 ;
        RECT 363.040 2670.400 363.300 2670.660 ;
        RECT 363.040 2656.460 363.300 2656.720 ;
        RECT 363.500 2621.440 363.760 2621.700 ;
        RECT 364.420 2621.440 364.680 2621.700 ;
        RECT 363.040 2511.620 363.300 2511.880 ;
        RECT 365.340 2511.620 365.600 2511.880 ;
        RECT 364.420 2401.120 364.680 2401.380 ;
        RECT 365.340 2401.120 365.600 2401.380 ;
        RECT 364.420 2304.560 364.680 2304.820 ;
        RECT 365.340 2304.560 365.600 2304.820 ;
        RECT 363.960 2187.260 364.220 2187.520 ;
        RECT 364.880 2187.260 365.140 2187.520 ;
        RECT 363.960 2122.660 364.220 2122.920 ;
        RECT 616.040 2122.660 616.300 2122.920 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.330 364.620 3298.410 ;
        RECT 364.020 3298.270 364.680 3298.330 ;
        RECT 364.420 3298.010 364.680 3298.270 ;
        RECT 365.340 3298.010 365.600 3298.330 ;
        RECT 365.400 3284.390 365.540 3298.010 ;
        RECT 365.340 3284.070 365.600 3284.390 ;
        RECT 364.880 3236.130 365.140 3236.450 ;
        RECT 364.940 3202.110 365.080 3236.130 ;
        RECT 364.880 3201.790 365.140 3202.110 ;
        RECT 363.960 3201.110 364.220 3201.430 ;
        RECT 364.020 3187.830 364.160 3201.110 ;
        RECT 363.960 3187.510 364.220 3187.830 ;
        RECT 364.420 3187.510 364.680 3187.830 ;
        RECT 364.480 3152.890 364.620 3187.510 ;
        RECT 364.480 3152.750 365.540 3152.890 ;
        RECT 365.400 3132.750 365.540 3152.750 ;
        RECT 365.340 3132.430 365.600 3132.750 ;
        RECT 365.340 3084.150 365.600 3084.470 ;
        RECT 365.400 3057.270 365.540 3084.150 ;
        RECT 365.340 3056.950 365.600 3057.270 ;
        RECT 364.420 3056.270 364.680 3056.590 ;
        RECT 364.480 3042.730 364.620 3056.270 ;
        RECT 364.870 3042.730 365.150 3042.845 ;
        RECT 364.480 3042.590 365.150 3042.730 ;
        RECT 364.870 3042.475 365.150 3042.590 ;
        RECT 365.790 3042.475 366.070 3042.845 ;
        RECT 365.860 3007.970 366.000 3042.475 ;
        RECT 364.880 3007.650 365.140 3007.970 ;
        RECT 365.800 3007.650 366.060 3007.970 ;
        RECT 364.940 2994.710 365.080 3007.650 ;
        RECT 364.880 2994.390 365.140 2994.710 ;
        RECT 364.420 2946.450 364.680 2946.770 ;
        RECT 364.480 2912.090 364.620 2946.450 ;
        RECT 363.500 2911.770 363.760 2912.090 ;
        RECT 364.420 2911.770 364.680 2912.090 ;
        RECT 363.560 2898.150 363.700 2911.770 ;
        RECT 363.500 2897.830 363.760 2898.150 ;
        RECT 363.040 2849.550 363.300 2849.870 ;
        RECT 363.100 2815.530 363.240 2849.550 ;
        RECT 363.040 2815.210 363.300 2815.530 ;
        RECT 363.500 2814.530 363.760 2814.850 ;
        RECT 363.560 2801.330 363.700 2814.530 ;
        RECT 363.100 2801.190 363.700 2801.330 ;
        RECT 363.100 2767.250 363.240 2801.190 ;
        RECT 363.040 2766.930 363.300 2767.250 ;
        RECT 363.040 2752.990 363.300 2753.310 ;
        RECT 363.100 2718.970 363.240 2752.990 ;
        RECT 363.040 2718.650 363.300 2718.970 ;
        RECT 363.500 2717.970 363.760 2718.290 ;
        RECT 363.560 2704.770 363.700 2717.970 ;
        RECT 363.100 2704.630 363.700 2704.770 ;
        RECT 363.100 2670.690 363.240 2704.630 ;
        RECT 363.040 2670.370 363.300 2670.690 ;
        RECT 363.100 2656.750 363.240 2656.905 ;
        RECT 363.040 2656.490 363.300 2656.750 ;
        RECT 363.490 2656.490 363.770 2656.605 ;
        RECT 363.040 2656.430 363.770 2656.490 ;
        RECT 363.100 2656.350 363.770 2656.430 ;
        RECT 363.490 2656.235 363.770 2656.350 ;
        RECT 364.410 2656.235 364.690 2656.605 ;
        RECT 364.480 2621.730 364.620 2656.235 ;
        RECT 363.500 2621.410 363.760 2621.730 ;
        RECT 364.420 2621.410 364.680 2621.730 ;
        RECT 363.560 2573.530 363.700 2621.410 ;
        RECT 363.560 2573.390 364.160 2573.530 ;
        RECT 364.020 2560.045 364.160 2573.390 ;
        RECT 363.030 2559.675 363.310 2560.045 ;
        RECT 363.950 2559.675 364.230 2560.045 ;
        RECT 363.100 2511.910 363.240 2559.675 ;
        RECT 363.040 2511.590 363.300 2511.910 ;
        RECT 365.340 2511.590 365.600 2511.910 ;
        RECT 365.400 2476.970 365.540 2511.590 ;
        RECT 364.940 2476.830 365.540 2476.970 ;
        RECT 364.940 2429.370 365.080 2476.830 ;
        RECT 364.480 2429.230 365.080 2429.370 ;
        RECT 364.480 2401.410 364.620 2429.230 ;
        RECT 364.420 2401.090 364.680 2401.410 ;
        RECT 365.340 2401.090 365.600 2401.410 ;
        RECT 365.400 2400.810 365.540 2401.090 ;
        RECT 364.940 2400.670 365.540 2400.810 ;
        RECT 364.940 2353.210 365.080 2400.670 ;
        RECT 364.480 2353.070 365.080 2353.210 ;
        RECT 364.480 2304.850 364.620 2353.070 ;
        RECT 364.420 2304.530 364.680 2304.850 ;
        RECT 365.340 2304.530 365.600 2304.850 ;
        RECT 365.400 2304.250 365.540 2304.530 ;
        RECT 364.940 2304.110 365.540 2304.250 ;
        RECT 364.940 2187.550 365.080 2304.110 ;
        RECT 363.960 2187.230 364.220 2187.550 ;
        RECT 364.880 2187.230 365.140 2187.550 ;
        RECT 364.020 2122.950 364.160 2187.230 ;
        RECT 363.960 2122.630 364.220 2122.950 ;
        RECT 616.040 2122.630 616.300 2122.950 ;
        RECT 616.100 2112.185 616.240 2122.630 ;
        RECT 616.100 2111.740 616.450 2112.185 ;
        RECT 616.170 2108.185 616.450 2111.740 ;
      LAYER via2 ;
        RECT 364.870 3042.520 365.150 3042.800 ;
        RECT 365.790 3042.520 366.070 3042.800 ;
        RECT 363.490 2656.280 363.770 2656.560 ;
        RECT 364.410 2656.280 364.690 2656.560 ;
        RECT 363.030 2559.720 363.310 2560.000 ;
        RECT 363.950 2559.720 364.230 2560.000 ;
      LAYER met3 ;
        RECT 364.845 3042.810 365.175 3042.825 ;
        RECT 365.765 3042.810 366.095 3042.825 ;
        RECT 364.845 3042.510 366.095 3042.810 ;
        RECT 364.845 3042.495 365.175 3042.510 ;
        RECT 365.765 3042.495 366.095 3042.510 ;
        RECT 363.465 2656.570 363.795 2656.585 ;
        RECT 364.385 2656.570 364.715 2656.585 ;
        RECT 363.465 2656.270 364.715 2656.570 ;
        RECT 363.465 2656.255 363.795 2656.270 ;
        RECT 364.385 2656.255 364.715 2656.270 ;
        RECT 363.005 2560.010 363.335 2560.025 ;
        RECT 363.925 2560.010 364.255 2560.025 ;
        RECT 363.005 2559.710 364.255 2560.010 ;
        RECT 363.005 2559.695 363.335 2559.710 ;
        RECT 363.925 2559.695 364.255 2559.710 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
        RECT 40.165 2898.585 40.335 2946.355 ;
        RECT 40.165 2704.785 40.335 2752.895 ;
        RECT 40.625 2186.965 40.795 2221.815 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
        RECT 40.165 2946.185 40.335 2946.355 ;
        RECT 40.165 2752.725 40.335 2752.895 ;
        RECT 40.625 2221.645 40.795 2221.815 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 40.090 2946.340 40.410 2946.400 ;
        RECT 39.895 2946.200 40.410 2946.340 ;
        RECT 40.090 2946.140 40.410 2946.200 ;
        RECT 40.090 2898.740 40.410 2898.800 ;
        RECT 39.895 2898.600 40.410 2898.740 ;
        RECT 40.090 2898.540 40.410 2898.600 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 40.550 2898.060 40.870 2898.120 ;
        RECT 39.630 2897.920 40.870 2898.060 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 40.550 2897.860 40.870 2897.920 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 40.550 2814.760 40.870 2814.820 ;
        RECT 39.630 2814.620 40.870 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.550 2814.560 40.870 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 39.895 2752.740 40.410 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.105 2704.940 40.395 2704.985 ;
        RECT 41.010 2704.940 41.330 2705.000 ;
        RECT 40.105 2704.800 41.330 2704.940 ;
        RECT 40.105 2704.755 40.395 2704.800 ;
        RECT 41.010 2704.740 41.330 2704.800 ;
        RECT 41.010 2608.380 41.330 2608.440 ;
        RECT 41.930 2608.380 42.250 2608.440 ;
        RECT 41.010 2608.240 42.250 2608.380 ;
        RECT 41.010 2608.180 41.330 2608.240 ;
        RECT 41.930 2608.180 42.250 2608.240 ;
        RECT 41.010 2511.820 41.330 2511.880 ;
        RECT 41.930 2511.820 42.250 2511.880 ;
        RECT 41.010 2511.680 42.250 2511.820 ;
        RECT 41.010 2511.620 41.330 2511.680 ;
        RECT 41.930 2511.620 42.250 2511.680 ;
        RECT 39.630 2463.200 39.950 2463.260 ;
        RECT 40.550 2463.200 40.870 2463.260 ;
        RECT 39.630 2463.060 40.870 2463.200 ;
        RECT 39.630 2463.000 39.950 2463.060 ;
        RECT 40.550 2463.000 40.870 2463.060 ;
        RECT 40.090 2366.640 40.410 2366.700 ;
        RECT 40.550 2366.640 40.870 2366.700 ;
        RECT 40.090 2366.500 40.870 2366.640 ;
        RECT 40.090 2366.440 40.410 2366.500 ;
        RECT 40.550 2366.440 40.870 2366.500 ;
        RECT 40.090 2235.540 40.410 2235.800 ;
        RECT 40.180 2235.400 40.320 2235.540 ;
        RECT 40.550 2235.400 40.870 2235.460 ;
        RECT 40.180 2235.260 40.870 2235.400 ;
        RECT 40.550 2235.200 40.870 2235.260 ;
        RECT 40.550 2221.800 40.870 2221.860 ;
        RECT 40.355 2221.660 40.870 2221.800 ;
        RECT 40.550 2221.600 40.870 2221.660 ;
        RECT 40.550 2187.120 40.870 2187.180 ;
        RECT 40.355 2186.980 40.870 2187.120 ;
        RECT 40.550 2186.920 40.870 2186.980 ;
        RECT 40.090 2125.580 40.410 2125.640 ;
        RECT 41.010 2125.580 41.330 2125.640 ;
        RECT 40.090 2125.440 41.330 2125.580 ;
        RECT 40.090 2125.380 40.410 2125.440 ;
        RECT 41.010 2125.380 41.330 2125.440 ;
        RECT 40.090 2121.840 40.410 2121.900 ;
        RECT 439.370 2121.840 439.690 2121.900 ;
        RECT 40.090 2121.700 439.690 2121.840 ;
        RECT 40.090 2121.640 40.410 2121.700 ;
        RECT 439.370 2121.640 439.690 2121.700 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 40.120 2946.140 40.380 2946.400 ;
        RECT 40.120 2898.540 40.380 2898.800 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 40.580 2897.860 40.840 2898.120 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.580 2814.560 40.840 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 41.040 2704.740 41.300 2705.000 ;
        RECT 41.040 2608.180 41.300 2608.440 ;
        RECT 41.960 2608.180 42.220 2608.440 ;
        RECT 41.040 2511.620 41.300 2511.880 ;
        RECT 41.960 2511.620 42.220 2511.880 ;
        RECT 39.660 2463.000 39.920 2463.260 ;
        RECT 40.580 2463.000 40.840 2463.260 ;
        RECT 40.120 2366.440 40.380 2366.700 ;
        RECT 40.580 2366.440 40.840 2366.700 ;
        RECT 40.120 2235.540 40.380 2235.800 ;
        RECT 40.580 2235.200 40.840 2235.460 ;
        RECT 40.580 2221.600 40.840 2221.860 ;
        RECT 40.580 2186.920 40.840 2187.180 ;
        RECT 40.120 2125.380 40.380 2125.640 ;
        RECT 41.040 2125.380 41.300 2125.640 ;
        RECT 40.120 2121.640 40.380 2121.900 ;
        RECT 439.400 2121.640 439.660 2121.900 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2946.430 40.320 2959.630 ;
        RECT 40.120 2946.110 40.380 2946.430 ;
        RECT 40.120 2898.570 40.380 2898.830 ;
        RECT 39.720 2898.510 40.380 2898.570 ;
        RECT 39.720 2898.430 40.320 2898.510 ;
        RECT 39.720 2898.150 39.860 2898.430 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 40.580 2897.830 40.840 2898.150 ;
        RECT 40.640 2814.850 40.780 2897.830 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 40.580 2814.530 40.840 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 41.040 2704.710 41.300 2705.030 ;
        RECT 41.100 2670.090 41.240 2704.710 ;
        RECT 40.640 2669.950 41.240 2670.090 ;
        RECT 40.640 2656.605 40.780 2669.950 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.950 2656.235 42.230 2656.605 ;
        RECT 42.020 2608.470 42.160 2656.235 ;
        RECT 41.040 2608.150 41.300 2608.470 ;
        RECT 41.960 2608.150 42.220 2608.470 ;
        RECT 41.100 2573.530 41.240 2608.150 ;
        RECT 40.640 2573.390 41.240 2573.530 ;
        RECT 40.640 2560.045 40.780 2573.390 ;
        RECT 40.570 2559.675 40.850 2560.045 ;
        RECT 41.950 2559.675 42.230 2560.045 ;
        RECT 42.020 2511.910 42.160 2559.675 ;
        RECT 41.040 2511.590 41.300 2511.910 ;
        RECT 41.960 2511.590 42.220 2511.910 ;
        RECT 41.100 2476.970 41.240 2511.590 ;
        RECT 40.640 2476.830 41.240 2476.970 ;
        RECT 40.640 2463.290 40.780 2476.830 ;
        RECT 39.660 2462.970 39.920 2463.290 ;
        RECT 40.580 2462.970 40.840 2463.290 ;
        RECT 39.720 2415.205 39.860 2462.970 ;
        RECT 39.650 2414.835 39.930 2415.205 ;
        RECT 41.030 2414.835 41.310 2415.205 ;
        RECT 41.100 2380.410 41.240 2414.835 ;
        RECT 40.180 2380.270 41.240 2380.410 ;
        RECT 40.180 2366.730 40.320 2380.270 ;
        RECT 40.120 2366.410 40.380 2366.730 ;
        RECT 40.580 2366.410 40.840 2366.730 ;
        RECT 40.640 2318.530 40.780 2366.410 ;
        RECT 40.640 2318.390 41.240 2318.530 ;
        RECT 41.100 2283.850 41.240 2318.390 ;
        RECT 40.180 2283.710 41.240 2283.850 ;
        RECT 40.180 2235.830 40.320 2283.710 ;
        RECT 40.120 2235.510 40.380 2235.830 ;
        RECT 40.580 2235.170 40.840 2235.490 ;
        RECT 40.640 2221.890 40.780 2235.170 ;
        RECT 40.580 2221.570 40.840 2221.890 ;
        RECT 40.580 2186.890 40.840 2187.210 ;
        RECT 40.640 2173.690 40.780 2186.890 ;
        RECT 40.640 2173.550 41.240 2173.690 ;
        RECT 41.100 2125.670 41.240 2173.550 ;
        RECT 40.120 2125.350 40.380 2125.670 ;
        RECT 41.040 2125.350 41.300 2125.670 ;
        RECT 40.180 2121.930 40.320 2125.350 ;
        RECT 40.120 2121.610 40.380 2121.930 ;
        RECT 439.400 2121.610 439.660 2121.930 ;
        RECT 439.460 2112.185 439.600 2121.610 ;
        RECT 439.460 2111.740 439.810 2112.185 ;
        RECT 439.530 2108.185 439.810 2111.740 ;
      LAYER via2 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.950 2656.280 42.230 2656.560 ;
        RECT 40.570 2559.720 40.850 2560.000 ;
        RECT 41.950 2559.720 42.230 2560.000 ;
        RECT 39.650 2414.880 39.930 2415.160 ;
        RECT 41.030 2414.880 41.310 2415.160 ;
      LAYER met3 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.925 2656.570 42.255 2656.585 ;
        RECT 40.545 2656.270 42.255 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.925 2656.255 42.255 2656.270 ;
        RECT 40.545 2560.010 40.875 2560.025 ;
        RECT 41.925 2560.010 42.255 2560.025 ;
        RECT 40.545 2559.710 42.255 2560.010 ;
        RECT 40.545 2559.695 40.875 2559.710 ;
        RECT 41.925 2559.695 42.255 2559.710 ;
        RECT 39.625 2415.170 39.955 2415.185 ;
        RECT 41.005 2415.170 41.335 2415.185 ;
        RECT 39.625 2414.870 41.335 2415.170 ;
        RECT 39.625 2414.855 39.955 2414.870 ;
        RECT 41.005 2414.855 41.335 2414.870 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 72.290 3263.900 72.610 3263.960 ;
        RECT 15.250 3263.760 72.610 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 72.290 3263.700 72.610 3263.760 ;
        RECT 72.290 2021.540 72.610 2021.600 ;
        RECT 393.370 2021.540 393.690 2021.600 ;
        RECT 72.290 2021.400 393.690 2021.540 ;
        RECT 72.290 2021.340 72.610 2021.400 ;
        RECT 393.370 2021.340 393.690 2021.400 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 72.320 3263.700 72.580 3263.960 ;
        RECT 72.320 2021.340 72.580 2021.600 ;
        RECT 393.400 2021.340 393.660 2021.600 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 72.320 3263.670 72.580 3263.990 ;
        RECT 72.380 2021.630 72.520 3263.670 ;
        RECT 72.320 2021.310 72.580 2021.630 ;
        RECT 393.400 2021.310 393.660 2021.630 ;
        RECT 393.460 2016.725 393.600 2021.310 ;
        RECT 393.390 2016.355 393.670 2016.725 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 393.390 2016.400 393.670 2016.680 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 393.365 2016.690 393.695 2016.705 ;
        RECT 410.000 2016.690 414.000 2016.840 ;
        RECT 393.365 2016.390 414.000 2016.690 ;
        RECT 393.365 2016.375 393.695 2016.390 ;
        RECT 410.000 2016.240 414.000 2016.390 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 224.090 2974.220 224.410 2974.280 ;
        RECT 16.630 2974.080 224.410 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 224.090 2974.020 224.410 2974.080 ;
        RECT 224.090 1904.240 224.410 1904.300 ;
        RECT 393.370 1904.240 393.690 1904.300 ;
        RECT 224.090 1904.100 393.690 1904.240 ;
        RECT 224.090 1904.040 224.410 1904.100 ;
        RECT 393.370 1904.040 393.690 1904.100 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 224.120 2974.020 224.380 2974.280 ;
        RECT 224.120 1904.040 224.380 1904.300 ;
        RECT 393.400 1904.040 393.660 1904.300 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 224.120 2973.990 224.380 2974.310 ;
        RECT 224.180 1904.330 224.320 2973.990 ;
        RECT 224.120 1904.010 224.380 1904.330 ;
        RECT 393.400 1904.010 393.660 1904.330 ;
        RECT 393.460 1902.485 393.600 1904.010 ;
        RECT 393.390 1902.115 393.670 1902.485 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
        RECT 393.390 1902.160 393.670 1902.440 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
        RECT 393.365 1902.450 393.695 1902.465 ;
        RECT 410.000 1902.450 414.000 1902.600 ;
        RECT 393.365 1902.150 414.000 1902.450 ;
        RECT 393.365 1902.135 393.695 1902.150 ;
        RECT 410.000 1902.000 414.000 1902.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2691.340 20.630 2691.400 ;
        RECT 86.090 2691.340 86.410 2691.400 ;
        RECT 20.310 2691.200 86.410 2691.340 ;
        RECT 20.310 2691.140 20.630 2691.200 ;
        RECT 86.090 2691.140 86.410 2691.200 ;
        RECT 86.090 1793.740 86.410 1793.800 ;
        RECT 393.370 1793.740 393.690 1793.800 ;
        RECT 86.090 1793.600 393.690 1793.740 ;
        RECT 86.090 1793.540 86.410 1793.600 ;
        RECT 393.370 1793.540 393.690 1793.600 ;
      LAYER via ;
        RECT 20.340 2691.140 20.600 2691.400 ;
        RECT 86.120 2691.140 86.380 2691.400 ;
        RECT 86.120 1793.540 86.380 1793.800 ;
        RECT 393.400 1793.540 393.660 1793.800 ;
      LAYER met2 ;
        RECT 20.330 2692.955 20.610 2693.325 ;
        RECT 20.400 2691.430 20.540 2692.955 ;
        RECT 20.340 2691.110 20.600 2691.430 ;
        RECT 86.120 2691.110 86.380 2691.430 ;
        RECT 86.180 1793.830 86.320 2691.110 ;
        RECT 86.120 1793.510 86.380 1793.830 ;
        RECT 393.400 1793.510 393.660 1793.830 ;
        RECT 393.460 1788.245 393.600 1793.510 ;
        RECT 393.390 1787.875 393.670 1788.245 ;
      LAYER via2 ;
        RECT 20.330 2693.000 20.610 2693.280 ;
        RECT 393.390 1787.920 393.670 1788.200 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 20.305 2693.290 20.635 2693.305 ;
        RECT -4.800 2692.990 20.635 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 20.305 2692.975 20.635 2692.990 ;
        RECT 393.365 1788.210 393.695 1788.225 ;
        RECT 410.000 1788.210 414.000 1788.360 ;
        RECT 393.365 1787.910 414.000 1788.210 ;
        RECT 393.365 1787.895 393.695 1787.910 ;
        RECT 410.000 1787.760 414.000 1787.910 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2401.320 16.030 2401.380 ;
        RECT 51.590 2401.320 51.910 2401.380 ;
        RECT 15.710 2401.180 51.910 2401.320 ;
        RECT 15.710 2401.120 16.030 2401.180 ;
        RECT 51.590 2401.120 51.910 2401.180 ;
        RECT 51.590 1676.440 51.910 1676.500 ;
        RECT 393.370 1676.440 393.690 1676.500 ;
        RECT 51.590 1676.300 393.690 1676.440 ;
        RECT 51.590 1676.240 51.910 1676.300 ;
        RECT 393.370 1676.240 393.690 1676.300 ;
      LAYER via ;
        RECT 15.740 2401.120 16.000 2401.380 ;
        RECT 51.620 2401.120 51.880 2401.380 ;
        RECT 51.620 1676.240 51.880 1676.500 ;
        RECT 393.400 1676.240 393.660 1676.500 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.800 2401.410 15.940 2405.315 ;
        RECT 15.740 2401.090 16.000 2401.410 ;
        RECT 51.620 2401.090 51.880 2401.410 ;
        RECT 51.680 1676.530 51.820 2401.090 ;
        RECT 51.620 1676.210 51.880 1676.530 ;
        RECT 393.400 1676.210 393.660 1676.530 ;
        RECT 393.460 1673.325 393.600 1676.210 ;
        RECT 393.390 1672.955 393.670 1673.325 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
        RECT 393.390 1673.000 393.670 1673.280 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
        RECT 393.365 1673.290 393.695 1673.305 ;
        RECT 410.000 1673.290 414.000 1673.440 ;
        RECT 393.365 1672.990 414.000 1673.290 ;
        RECT 393.365 1672.975 393.695 1672.990 ;
        RECT 410.000 1672.840 414.000 1672.990 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2118.440 16.950 2118.500 ;
        RECT 37.790 2118.440 38.110 2118.500 ;
        RECT 16.630 2118.300 38.110 2118.440 ;
        RECT 16.630 2118.240 16.950 2118.300 ;
        RECT 37.790 2118.240 38.110 2118.300 ;
        RECT 37.790 1559.140 38.110 1559.200 ;
        RECT 393.370 1559.140 393.690 1559.200 ;
        RECT 37.790 1559.000 393.690 1559.140 ;
        RECT 37.790 1558.940 38.110 1559.000 ;
        RECT 393.370 1558.940 393.690 1559.000 ;
      LAYER via ;
        RECT 16.660 2118.240 16.920 2118.500 ;
        RECT 37.820 2118.240 38.080 2118.500 ;
        RECT 37.820 1558.940 38.080 1559.200 ;
        RECT 393.400 1558.940 393.660 1559.200 ;
      LAYER met2 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
        RECT 16.660 2118.210 16.920 2118.355 ;
        RECT 37.820 2118.210 38.080 2118.530 ;
        RECT 37.880 1559.230 38.020 2118.210 ;
        RECT 37.820 1558.910 38.080 1559.230 ;
        RECT 393.400 1559.085 393.660 1559.230 ;
        RECT 393.390 1558.715 393.670 1559.085 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
        RECT 393.390 1558.760 393.670 1559.040 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
        RECT 393.365 1559.050 393.695 1559.065 ;
        RECT 410.000 1559.050 414.000 1559.200 ;
        RECT 393.365 1558.750 414.000 1559.050 ;
        RECT 393.365 1558.735 393.695 1558.750 ;
        RECT 410.000 1558.600 414.000 1558.750 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1448.980 17.870 1449.040 ;
        RECT 393.370 1448.980 393.690 1449.040 ;
        RECT 17.550 1448.840 393.690 1448.980 ;
        RECT 17.550 1448.780 17.870 1448.840 ;
        RECT 393.370 1448.780 393.690 1448.840 ;
      LAYER via ;
        RECT 17.580 1448.780 17.840 1449.040 ;
        RECT 393.400 1448.780 393.660 1449.040 ;
      LAYER met2 ;
        RECT 17.570 1830.715 17.850 1831.085 ;
        RECT 17.640 1449.070 17.780 1830.715 ;
        RECT 17.580 1448.750 17.840 1449.070 ;
        RECT 393.400 1448.750 393.660 1449.070 ;
        RECT 393.460 1444.845 393.600 1448.750 ;
        RECT 393.390 1444.475 393.670 1444.845 ;
      LAYER via2 ;
        RECT 17.570 1830.760 17.850 1831.040 ;
        RECT 393.390 1444.520 393.670 1444.800 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 17.545 1831.050 17.875 1831.065 ;
        RECT -4.800 1830.750 17.875 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 17.545 1830.735 17.875 1830.750 ;
        RECT 393.365 1444.810 393.695 1444.825 ;
        RECT 410.000 1444.810 414.000 1444.960 ;
        RECT 393.365 1444.510 414.000 1444.810 ;
        RECT 393.365 1444.495 393.695 1444.510 ;
        RECT 410.000 1444.360 414.000 1444.510 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.650 676.160 2011.970 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2011.650 676.020 2901.150 676.160 ;
        RECT 2011.650 675.960 2011.970 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2011.680 675.960 2011.940 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2011.670 812.075 2011.950 812.445 ;
        RECT 2011.740 676.250 2011.880 812.075 ;
        RECT 2011.680 675.930 2011.940 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2011.670 812.120 2011.950 812.400 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 1997.465 812.410 2001.465 812.560 ;
        RECT 2011.645 812.410 2011.975 812.425 ;
        RECT 1997.465 812.110 2011.975 812.410 ;
        RECT 1997.465 811.960 2001.465 812.110 ;
        RECT 2011.645 812.095 2011.975 812.110 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 1331.680 18.790 1331.740 ;
        RECT 393.370 1331.680 393.690 1331.740 ;
        RECT 18.470 1331.540 393.690 1331.680 ;
        RECT 18.470 1331.480 18.790 1331.540 ;
        RECT 393.370 1331.480 393.690 1331.540 ;
      LAYER via ;
        RECT 18.500 1331.480 18.760 1331.740 ;
        RECT 393.400 1331.480 393.660 1331.740 ;
      LAYER met2 ;
        RECT 18.490 1543.755 18.770 1544.125 ;
        RECT 18.560 1331.770 18.700 1543.755 ;
        RECT 18.500 1331.450 18.760 1331.770 ;
        RECT 393.400 1331.450 393.660 1331.770 ;
        RECT 393.460 1330.605 393.600 1331.450 ;
        RECT 393.390 1330.235 393.670 1330.605 ;
      LAYER via2 ;
        RECT 18.490 1543.800 18.770 1544.080 ;
        RECT 393.390 1330.280 393.670 1330.560 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 18.465 1544.090 18.795 1544.105 ;
        RECT -4.800 1543.790 18.795 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 18.465 1543.775 18.795 1543.790 ;
        RECT 393.365 1330.570 393.695 1330.585 ;
        RECT 410.000 1330.570 414.000 1330.720 ;
        RECT 393.365 1330.270 414.000 1330.570 ;
        RECT 393.365 1330.255 393.695 1330.270 ;
        RECT 410.000 1330.120 414.000 1330.270 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 1221.180 18.330 1221.240 ;
        RECT 393.370 1221.180 393.690 1221.240 ;
        RECT 18.010 1221.040 393.690 1221.180 ;
        RECT 18.010 1220.980 18.330 1221.040 ;
        RECT 393.370 1220.980 393.690 1221.040 ;
      LAYER via ;
        RECT 18.040 1220.980 18.300 1221.240 ;
        RECT 393.400 1220.980 393.660 1221.240 ;
      LAYER met2 ;
        RECT 18.030 1328.195 18.310 1328.565 ;
        RECT 18.100 1221.270 18.240 1328.195 ;
        RECT 18.040 1220.950 18.300 1221.270 ;
        RECT 393.400 1220.950 393.660 1221.270 ;
        RECT 393.460 1215.685 393.600 1220.950 ;
        RECT 393.390 1215.315 393.670 1215.685 ;
      LAYER via2 ;
        RECT 18.030 1328.240 18.310 1328.520 ;
        RECT 393.390 1215.360 393.670 1215.640 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 18.005 1328.530 18.335 1328.545 ;
        RECT -4.800 1328.230 18.335 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 18.005 1328.215 18.335 1328.230 ;
        RECT 393.365 1215.650 393.695 1215.665 ;
        RECT 410.000 1215.650 414.000 1215.800 ;
        RECT 393.365 1215.350 414.000 1215.650 ;
        RECT 393.365 1215.335 393.695 1215.350 ;
        RECT 410.000 1215.200 414.000 1215.350 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1103.880 15.110 1103.940 ;
        RECT 393.370 1103.880 393.690 1103.940 ;
        RECT 14.790 1103.740 393.690 1103.880 ;
        RECT 14.790 1103.680 15.110 1103.740 ;
        RECT 393.370 1103.680 393.690 1103.740 ;
      LAYER via ;
        RECT 14.820 1103.680 15.080 1103.940 ;
        RECT 393.400 1103.680 393.660 1103.940 ;
      LAYER met2 ;
        RECT 14.810 1112.635 15.090 1113.005 ;
        RECT 14.880 1103.970 15.020 1112.635 ;
        RECT 14.820 1103.650 15.080 1103.970 ;
        RECT 393.400 1103.650 393.660 1103.970 ;
        RECT 393.460 1101.445 393.600 1103.650 ;
        RECT 393.390 1101.075 393.670 1101.445 ;
      LAYER via2 ;
        RECT 14.810 1112.680 15.090 1112.960 ;
        RECT 393.390 1101.120 393.670 1101.400 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 14.785 1112.970 15.115 1112.985 ;
        RECT -4.800 1112.670 15.115 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 14.785 1112.655 15.115 1112.670 ;
        RECT 393.365 1101.410 393.695 1101.425 ;
        RECT 410.000 1101.410 414.000 1101.560 ;
        RECT 393.365 1101.110 414.000 1101.410 ;
        RECT 393.365 1101.095 393.695 1101.110 ;
        RECT 410.000 1100.960 414.000 1101.110 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 397.050 903.960 397.370 904.020 ;
        RECT 16.170 903.820 397.370 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 397.050 903.760 397.370 903.820 ;
      LAYER via ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 397.080 903.760 397.340 904.020 ;
      LAYER met2 ;
        RECT 397.070 986.835 397.350 987.205 ;
        RECT 397.140 904.050 397.280 986.835 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 397.080 903.730 397.340 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 397.070 986.880 397.350 987.160 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 397.045 987.170 397.375 987.185 ;
        RECT 410.000 987.170 414.000 987.320 ;
        RECT 397.045 986.870 414.000 987.170 ;
        RECT 397.045 986.855 397.375 986.870 ;
        RECT 410.000 986.720 414.000 986.870 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 397.050 682.960 397.370 683.020 ;
        RECT 16.170 682.820 397.370 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 397.050 682.760 397.370 682.820 ;
      LAYER via ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 397.080 682.760 397.340 683.020 ;
      LAYER met2 ;
        RECT 397.070 871.915 397.350 872.285 ;
        RECT 397.140 683.050 397.280 871.915 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 397.080 682.730 397.340 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 397.070 871.960 397.350 872.240 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 397.045 872.250 397.375 872.265 ;
        RECT 410.000 872.250 414.000 872.400 ;
        RECT 397.045 871.950 414.000 872.250 ;
        RECT 397.045 871.935 397.375 871.950 ;
        RECT 410.000 871.800 414.000 871.950 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 398.430 469.100 398.750 469.160 ;
        RECT 17.090 468.960 398.750 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 398.430 468.900 398.750 468.960 ;
      LAYER via ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 398.460 468.900 398.720 469.160 ;
      LAYER met2 ;
        RECT 398.450 757.675 398.730 758.045 ;
        RECT 398.520 469.190 398.660 757.675 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 398.460 468.870 398.720 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 398.450 757.720 398.730 758.000 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 398.425 758.010 398.755 758.025 ;
        RECT 410.000 758.010 414.000 758.160 ;
        RECT 398.425 757.710 414.000 758.010 ;
        RECT 398.425 757.695 398.755 757.710 ;
        RECT 410.000 757.560 414.000 757.710 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 397.510 255.240 397.830 255.300 ;
        RECT 17.090 255.100 397.830 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 397.510 255.040 397.830 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 397.540 255.040 397.800 255.300 ;
      LAYER met2 ;
        RECT 397.530 643.435 397.810 643.805 ;
        RECT 397.600 255.330 397.740 643.435 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 397.540 255.010 397.800 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 397.530 643.480 397.810 643.760 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 397.505 643.770 397.835 643.785 ;
        RECT 410.000 643.770 414.000 643.920 ;
        RECT 397.505 643.470 414.000 643.770 ;
        RECT 397.505 643.455 397.835 643.470 ;
        RECT 410.000 643.320 414.000 643.470 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 396.590 41.380 396.910 41.440 ;
        RECT 17.090 41.240 396.910 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 396.590 41.180 396.910 41.240 ;
      LAYER via ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 396.620 41.180 396.880 41.440 ;
      LAYER met2 ;
        RECT 396.610 529.195 396.890 529.565 ;
        RECT 396.680 41.470 396.820 529.195 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 396.620 41.150 396.880 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 396.610 529.240 396.890 529.520 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 396.585 529.530 396.915 529.545 ;
        RECT 410.000 529.530 414.000 529.680 ;
        RECT 396.585 529.230 414.000 529.530 ;
        RECT 396.585 529.215 396.915 529.230 ;
        RECT 410.000 529.080 414.000 529.230 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 910.760 2008.290 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2007.970 910.620 2901.150 910.760 ;
        RECT 2007.970 910.560 2008.290 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2008.000 910.560 2008.260 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2007.990 918.835 2008.270 919.205 ;
        RECT 2008.060 910.850 2008.200 918.835 ;
        RECT 2008.000 910.530 2008.260 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2007.990 918.880 2008.270 919.160 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 1997.465 919.170 2001.465 919.320 ;
        RECT 2007.965 919.170 2008.295 919.185 ;
        RECT 1997.465 918.870 2008.295 919.170 ;
        RECT 1997.465 918.720 2001.465 918.870 ;
        RECT 2007.965 918.855 2008.295 918.870 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2024.990 1138.900 2025.310 1138.960 ;
        RECT 2900.830 1138.900 2901.150 1138.960 ;
        RECT 2024.990 1138.760 2901.150 1138.900 ;
        RECT 2024.990 1138.700 2025.310 1138.760 ;
        RECT 2900.830 1138.700 2901.150 1138.760 ;
        RECT 2007.970 1028.060 2008.290 1028.120 ;
        RECT 2024.990 1028.060 2025.310 1028.120 ;
        RECT 2007.970 1027.920 2025.310 1028.060 ;
        RECT 2007.970 1027.860 2008.290 1027.920 ;
        RECT 2024.990 1027.860 2025.310 1027.920 ;
      LAYER via ;
        RECT 2025.020 1138.700 2025.280 1138.960 ;
        RECT 2900.860 1138.700 2901.120 1138.960 ;
        RECT 2008.000 1027.860 2008.260 1028.120 ;
        RECT 2025.020 1027.860 2025.280 1028.120 ;
      LAYER met2 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
        RECT 2900.920 1138.990 2901.060 1143.915 ;
        RECT 2025.020 1138.670 2025.280 1138.990 ;
        RECT 2900.860 1138.670 2901.120 1138.990 ;
        RECT 2025.080 1028.150 2025.220 1138.670 ;
        RECT 2008.000 1027.830 2008.260 1028.150 ;
        RECT 2025.020 1027.830 2025.280 1028.150 ;
        RECT 2008.060 1025.965 2008.200 1027.830 ;
        RECT 2007.990 1025.595 2008.270 1025.965 ;
      LAYER via2 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
        RECT 2007.990 1025.640 2008.270 1025.920 ;
      LAYER met3 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 1997.465 1025.930 2001.465 1026.080 ;
        RECT 2007.965 1025.930 2008.295 1025.945 ;
        RECT 1997.465 1025.630 2008.295 1025.930 ;
        RECT 1997.465 1025.480 2001.465 1025.630 ;
        RECT 2007.965 1025.615 2008.295 1025.630 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2128.490 1373.500 2128.810 1373.560 ;
        RECT 2900.830 1373.500 2901.150 1373.560 ;
        RECT 2128.490 1373.360 2901.150 1373.500 ;
        RECT 2128.490 1373.300 2128.810 1373.360 ;
        RECT 2900.830 1373.300 2901.150 1373.360 ;
        RECT 2007.970 1138.560 2008.290 1138.620 ;
        RECT 2128.490 1138.560 2128.810 1138.620 ;
        RECT 2007.970 1138.420 2128.810 1138.560 ;
        RECT 2007.970 1138.360 2008.290 1138.420 ;
        RECT 2128.490 1138.360 2128.810 1138.420 ;
      LAYER via ;
        RECT 2128.520 1373.300 2128.780 1373.560 ;
        RECT 2900.860 1373.300 2901.120 1373.560 ;
        RECT 2008.000 1138.360 2008.260 1138.620 ;
        RECT 2128.520 1138.360 2128.780 1138.620 ;
      LAYER met2 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
        RECT 2900.920 1373.590 2901.060 1378.515 ;
        RECT 2128.520 1373.270 2128.780 1373.590 ;
        RECT 2900.860 1373.270 2901.120 1373.590 ;
        RECT 2128.580 1138.650 2128.720 1373.270 ;
        RECT 2008.000 1138.330 2008.260 1138.650 ;
        RECT 2128.520 1138.330 2128.780 1138.650 ;
        RECT 2008.060 1133.405 2008.200 1138.330 ;
        RECT 2007.990 1133.035 2008.270 1133.405 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
        RECT 2007.990 1133.080 2008.270 1133.360 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 1997.465 1133.370 2001.465 1133.520 ;
        RECT 2007.965 1133.370 2008.295 1133.385 ;
        RECT 1997.465 1133.070 2008.295 1133.370 ;
        RECT 1997.465 1132.920 2001.465 1133.070 ;
        RECT 2007.965 1133.055 2008.295 1133.070 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.190 1528.200 2011.510 1528.260 ;
        RECT 2894.390 1528.200 2894.710 1528.260 ;
        RECT 2011.190 1528.060 2894.710 1528.200 ;
        RECT 2011.190 1528.000 2011.510 1528.060 ;
        RECT 2894.390 1528.000 2894.710 1528.060 ;
      LAYER via ;
        RECT 2011.220 1528.000 2011.480 1528.260 ;
        RECT 2894.420 1528.000 2894.680 1528.260 ;
      LAYER met2 ;
        RECT 2894.410 1613.115 2894.690 1613.485 ;
        RECT 2894.480 1528.290 2894.620 1613.115 ;
        RECT 2011.220 1527.970 2011.480 1528.290 ;
        RECT 2894.420 1527.970 2894.680 1528.290 ;
        RECT 2011.280 1240.165 2011.420 1527.970 ;
        RECT 2011.210 1239.795 2011.490 1240.165 ;
      LAYER via2 ;
        RECT 2894.410 1613.160 2894.690 1613.440 ;
        RECT 2011.210 1239.840 2011.490 1240.120 ;
      LAYER met3 ;
        RECT 2894.385 1613.450 2894.715 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2894.385 1613.150 2924.800 1613.450 ;
        RECT 2894.385 1613.135 2894.715 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 1997.465 1240.130 2001.465 1240.280 ;
        RECT 2011.185 1240.130 2011.515 1240.145 ;
        RECT 1997.465 1239.830 2011.515 1240.130 ;
        RECT 1997.465 1239.680 2001.465 1239.830 ;
        RECT 2011.185 1239.815 2011.515 1239.830 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2880.590 1842.700 2880.910 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2880.590 1842.560 2901.150 1842.700 ;
        RECT 2880.590 1842.500 2880.910 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
        RECT 2007.970 1352.420 2008.290 1352.480 ;
        RECT 2880.590 1352.420 2880.910 1352.480 ;
        RECT 2007.970 1352.280 2880.910 1352.420 ;
        RECT 2007.970 1352.220 2008.290 1352.280 ;
        RECT 2880.590 1352.220 2880.910 1352.280 ;
      LAYER via ;
        RECT 2880.620 1842.500 2880.880 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
        RECT 2008.000 1352.220 2008.260 1352.480 ;
        RECT 2880.620 1352.220 2880.880 1352.480 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2880.620 1842.470 2880.880 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 2880.680 1352.510 2880.820 1842.470 ;
        RECT 2008.000 1352.190 2008.260 1352.510 ;
        RECT 2880.620 1352.190 2880.880 1352.510 ;
        RECT 2008.060 1346.925 2008.200 1352.190 ;
        RECT 2007.990 1346.555 2008.270 1346.925 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
        RECT 2007.990 1346.600 2008.270 1346.880 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 1997.465 1346.890 2001.465 1347.040 ;
        RECT 2007.965 1346.890 2008.295 1346.905 ;
        RECT 1997.465 1346.590 2008.295 1346.890 ;
        RECT 1997.465 1346.440 2001.465 1346.590 ;
        RECT 2007.965 1346.575 2008.295 1346.590 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2128.490 2077.300 2128.810 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2128.490 2077.160 2901.150 2077.300 ;
        RECT 2128.490 2077.100 2128.810 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 2007.970 1455.780 2008.290 1455.840 ;
        RECT 2128.490 1455.780 2128.810 1455.840 ;
        RECT 2007.970 1455.640 2128.810 1455.780 ;
        RECT 2007.970 1455.580 2008.290 1455.640 ;
        RECT 2128.490 1455.580 2128.810 1455.640 ;
      LAYER via ;
        RECT 2128.520 2077.100 2128.780 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 2008.000 1455.580 2008.260 1455.840 ;
        RECT 2128.520 1455.580 2128.780 1455.840 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2128.520 2077.070 2128.780 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2128.580 1455.870 2128.720 2077.070 ;
        RECT 2008.000 1455.550 2008.260 1455.870 ;
        RECT 2128.520 1455.550 2128.780 1455.870 ;
        RECT 2008.060 1453.685 2008.200 1455.550 ;
        RECT 2007.990 1453.315 2008.270 1453.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2007.990 1453.360 2008.270 1453.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 1997.465 1453.650 2001.465 1453.800 ;
        RECT 2007.965 1453.650 2008.295 1453.665 ;
        RECT 1997.465 1453.350 2008.295 1453.650 ;
        RECT 1997.465 1453.200 2001.465 1453.350 ;
        RECT 2007.965 1453.335 2008.295 1453.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2859.890 2311.900 2860.210 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2859.890 2311.760 2901.150 2311.900 ;
        RECT 2859.890 2311.700 2860.210 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 2007.970 1566.280 2008.290 1566.340 ;
        RECT 2859.890 1566.280 2860.210 1566.340 ;
        RECT 2007.970 1566.140 2860.210 1566.280 ;
        RECT 2007.970 1566.080 2008.290 1566.140 ;
        RECT 2859.890 1566.080 2860.210 1566.140 ;
      LAYER via ;
        RECT 2859.920 2311.700 2860.180 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 2008.000 1566.080 2008.260 1566.340 ;
        RECT 2859.920 1566.080 2860.180 1566.340 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2859.920 2311.670 2860.180 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2859.980 1566.370 2860.120 2311.670 ;
        RECT 2008.000 1566.050 2008.260 1566.370 ;
        RECT 2859.920 1566.050 2860.180 1566.370 ;
        RECT 2008.060 1560.445 2008.200 1566.050 ;
        RECT 2007.990 1560.075 2008.270 1560.445 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2007.990 1560.120 2008.270 1560.400 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 1997.465 1560.410 2001.465 1560.560 ;
        RECT 2007.965 1560.410 2008.295 1560.425 ;
        RECT 1997.465 1560.110 2008.295 1560.410 ;
        RECT 1997.465 1559.960 2001.465 1560.110 ;
        RECT 2007.965 1560.095 2008.295 1560.110 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.190 151.540 2011.510 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2011.190 151.400 2901.150 151.540 ;
        RECT 2011.190 151.340 2011.510 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2011.220 151.340 2011.480 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2011.210 563.195 2011.490 563.565 ;
        RECT 2011.280 151.630 2011.420 563.195 ;
        RECT 2011.220 151.310 2011.480 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2011.210 563.240 2011.490 563.520 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 1997.465 563.530 2001.465 563.680 ;
        RECT 2011.185 563.530 2011.515 563.545 ;
        RECT 1997.465 563.230 2011.515 563.530 ;
        RECT 1997.465 563.080 2001.465 563.230 ;
        RECT 2011.185 563.215 2011.515 563.230 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2846.090 2491.080 2846.410 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2846.090 2490.940 2901.150 2491.080 ;
        RECT 2846.090 2490.880 2846.410 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 2007.970 1635.300 2008.290 1635.360 ;
        RECT 2846.090 1635.300 2846.410 1635.360 ;
        RECT 2007.970 1635.160 2846.410 1635.300 ;
        RECT 2007.970 1635.100 2008.290 1635.160 ;
        RECT 2846.090 1635.100 2846.410 1635.160 ;
      LAYER via ;
        RECT 2846.120 2490.880 2846.380 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 2008.000 1635.100 2008.260 1635.360 ;
        RECT 2846.120 1635.100 2846.380 1635.360 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2846.120 2490.850 2846.380 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2846.180 1635.390 2846.320 2490.850 ;
        RECT 2008.000 1635.070 2008.260 1635.390 ;
        RECT 2846.120 1635.070 2846.380 1635.390 ;
        RECT 2008.060 1631.845 2008.200 1635.070 ;
        RECT 2007.990 1631.475 2008.270 1631.845 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2007.990 1631.520 2008.270 1631.800 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 1997.465 1631.810 2001.465 1631.960 ;
        RECT 2007.965 1631.810 2008.295 1631.825 ;
        RECT 1997.465 1631.510 2008.295 1631.810 ;
        RECT 1997.465 1631.360 2001.465 1631.510 ;
        RECT 2007.965 1631.495 2008.295 1631.510 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2763.290 2725.680 2763.610 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2763.290 2725.540 2901.150 2725.680 ;
        RECT 2763.290 2725.480 2763.610 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 2007.970 1738.660 2008.290 1738.720 ;
        RECT 2763.290 1738.660 2763.610 1738.720 ;
        RECT 2007.970 1738.520 2763.610 1738.660 ;
        RECT 2007.970 1738.460 2008.290 1738.520 ;
        RECT 2763.290 1738.460 2763.610 1738.520 ;
      LAYER via ;
        RECT 2763.320 2725.480 2763.580 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 2008.000 1738.460 2008.260 1738.720 ;
        RECT 2763.320 1738.460 2763.580 1738.720 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2763.320 2725.450 2763.580 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2763.380 1738.750 2763.520 2725.450 ;
        RECT 2008.000 1738.605 2008.260 1738.750 ;
        RECT 2007.990 1738.235 2008.270 1738.605 ;
        RECT 2763.320 1738.430 2763.580 1738.750 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2007.990 1738.280 2008.270 1738.560 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 1997.465 1738.570 2001.465 1738.720 ;
        RECT 2007.965 1738.570 2008.295 1738.585 ;
        RECT 1997.465 1738.270 2008.295 1738.570 ;
        RECT 1997.465 1738.120 2001.465 1738.270 ;
        RECT 2007.965 1738.255 2008.295 1738.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2852.990 2960.280 2853.310 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 2852.990 2960.140 2901.150 2960.280 ;
        RECT 2852.990 2960.080 2853.310 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
        RECT 2007.970 1849.160 2008.290 1849.220 ;
        RECT 2852.990 1849.160 2853.310 1849.220 ;
        RECT 2007.970 1849.020 2853.310 1849.160 ;
        RECT 2007.970 1848.960 2008.290 1849.020 ;
        RECT 2852.990 1848.960 2853.310 1849.020 ;
      LAYER via ;
        RECT 2853.020 2960.080 2853.280 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
        RECT 2008.000 1848.960 2008.260 1849.220 ;
        RECT 2853.020 1848.960 2853.280 1849.220 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 2853.020 2960.050 2853.280 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 2853.080 1849.250 2853.220 2960.050 ;
        RECT 2008.000 1848.930 2008.260 1849.250 ;
        RECT 2853.020 1848.930 2853.280 1849.250 ;
        RECT 2008.060 1845.365 2008.200 1848.930 ;
        RECT 2007.990 1844.995 2008.270 1845.365 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 2007.990 1845.040 2008.270 1845.320 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 1997.465 1845.330 2001.465 1845.480 ;
        RECT 2007.965 1845.330 2008.295 1845.345 ;
        RECT 1997.465 1845.030 2008.295 1845.330 ;
        RECT 1997.465 1844.880 2001.465 1845.030 ;
        RECT 2007.965 1845.015 2008.295 1845.030 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2866.790 3194.880 2867.110 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2866.790 3194.740 2901.150 3194.880 ;
        RECT 2866.790 3194.680 2867.110 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
        RECT 2007.970 1952.520 2008.290 1952.580 ;
        RECT 2866.790 1952.520 2867.110 1952.580 ;
        RECT 2007.970 1952.380 2867.110 1952.520 ;
        RECT 2007.970 1952.320 2008.290 1952.380 ;
        RECT 2866.790 1952.320 2867.110 1952.380 ;
      LAYER via ;
        RECT 2866.820 3194.680 2867.080 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
        RECT 2008.000 1952.320 2008.260 1952.580 ;
        RECT 2866.820 1952.320 2867.080 1952.580 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2866.820 3194.650 2867.080 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2866.880 1952.610 2867.020 3194.650 ;
        RECT 2008.000 1952.290 2008.260 1952.610 ;
        RECT 2866.820 1952.290 2867.080 1952.610 ;
        RECT 2008.060 1952.125 2008.200 1952.290 ;
        RECT 2007.990 1951.755 2008.270 1952.125 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2007.990 1951.800 2008.270 1952.080 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 1997.465 1952.090 2001.465 1952.240 ;
        RECT 2007.965 1952.090 2008.295 1952.105 ;
        RECT 1997.465 1951.790 2008.295 1952.090 ;
        RECT 1997.465 1951.640 2001.465 1951.790 ;
        RECT 2007.965 1951.775 2008.295 1951.790 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 2063.020 2008.290 2063.080 ;
        RECT 2901.290 2063.020 2901.610 2063.080 ;
        RECT 2007.970 2062.880 2901.610 2063.020 ;
        RECT 2007.970 2062.820 2008.290 2062.880 ;
        RECT 2901.290 2062.820 2901.610 2062.880 ;
      LAYER via ;
        RECT 2008.000 2062.820 2008.260 2063.080 ;
        RECT 2901.320 2062.820 2901.580 2063.080 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 2901.380 2063.110 2901.520 3431.435 ;
        RECT 2008.000 2062.790 2008.260 2063.110 ;
        RECT 2901.320 2062.790 2901.580 2063.110 ;
        RECT 2008.060 2058.885 2008.200 2062.790 ;
        RECT 2007.990 2058.515 2008.270 2058.885 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
        RECT 2007.990 2058.560 2008.270 2058.840 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 1997.465 2058.850 2001.465 2059.000 ;
        RECT 2007.965 2058.850 2008.295 2058.865 ;
        RECT 1997.465 2058.550 2008.295 2058.850 ;
        RECT 1997.465 2058.400 2001.465 2058.550 ;
        RECT 2007.965 2058.535 2008.295 2058.550 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3415.555 ;
        RECT 2712.765 3008.405 2712.935 3042.915 ;
        RECT 2713.685 2946.525 2713.855 2994.635 ;
        RECT 2712.305 2753.065 2712.475 2801.175 ;
        RECT 2712.765 2428.705 2712.935 2463.215 ;
        RECT 2712.765 2331.805 2712.935 2366.655 ;
        RECT 2712.765 2138.685 2712.935 2173.535 ;
      LAYER mcon ;
        RECT 2713.685 3415.385 2713.855 3415.555 ;
        RECT 2712.765 3042.745 2712.935 3042.915 ;
        RECT 2713.685 2994.465 2713.855 2994.635 ;
        RECT 2712.305 2801.005 2712.475 2801.175 ;
        RECT 2712.765 2463.045 2712.935 2463.215 ;
        RECT 2712.765 2366.485 2712.935 2366.655 ;
        RECT 2712.765 2173.365 2712.935 2173.535 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2712.690 3470.620 2713.010 3470.680 ;
        RECT 2713.610 3470.620 2713.930 3470.680 ;
        RECT 2712.690 3470.480 2713.930 3470.620 ;
        RECT 2712.690 3470.420 2713.010 3470.480 ;
        RECT 2713.610 3470.420 2713.930 3470.480 ;
        RECT 2712.690 3463.820 2713.010 3463.880 ;
        RECT 2713.610 3463.820 2713.930 3463.880 ;
        RECT 2712.690 3463.680 2713.930 3463.820 ;
        RECT 2712.690 3463.620 2713.010 3463.680 ;
        RECT 2713.610 3463.620 2713.930 3463.680 ;
        RECT 2711.770 3415.540 2712.090 3415.600 ;
        RECT 2713.625 3415.540 2713.915 3415.585 ;
        RECT 2711.770 3415.400 2713.915 3415.540 ;
        RECT 2711.770 3415.340 2712.090 3415.400 ;
        RECT 2713.625 3415.355 2713.915 3415.400 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2712.690 3042.900 2713.010 3042.960 ;
        RECT 2712.495 3042.760 2713.010 3042.900 ;
        RECT 2712.690 3042.700 2713.010 3042.760 ;
        RECT 2712.705 3008.560 2712.995 3008.605 ;
        RECT 2713.610 3008.560 2713.930 3008.620 ;
        RECT 2712.705 3008.420 2713.930 3008.560 ;
        RECT 2712.705 3008.375 2712.995 3008.420 ;
        RECT 2713.610 3008.360 2713.930 3008.420 ;
        RECT 2713.610 2994.620 2713.930 2994.680 ;
        RECT 2713.415 2994.480 2713.930 2994.620 ;
        RECT 2713.610 2994.420 2713.930 2994.480 ;
        RECT 2713.625 2946.680 2713.915 2946.725 ;
        RECT 2714.070 2946.680 2714.390 2946.740 ;
        RECT 2713.625 2946.540 2714.390 2946.680 ;
        RECT 2713.625 2946.495 2713.915 2946.540 ;
        RECT 2714.070 2946.480 2714.390 2946.540 ;
        RECT 2714.070 2912.340 2714.390 2912.400 ;
        RECT 2713.700 2912.200 2714.390 2912.340 ;
        RECT 2713.700 2911.720 2713.840 2912.200 ;
        RECT 2714.070 2912.140 2714.390 2912.200 ;
        RECT 2713.610 2911.460 2713.930 2911.720 ;
        RECT 2712.230 2815.580 2712.550 2815.840 ;
        RECT 2712.320 2815.160 2712.460 2815.580 ;
        RECT 2712.230 2814.900 2712.550 2815.160 ;
        RECT 2712.230 2801.160 2712.550 2801.220 ;
        RECT 2712.035 2801.020 2712.550 2801.160 ;
        RECT 2712.230 2800.960 2712.550 2801.020 ;
        RECT 2712.245 2753.220 2712.535 2753.265 ;
        RECT 2713.150 2753.220 2713.470 2753.280 ;
        RECT 2712.245 2753.080 2713.470 2753.220 ;
        RECT 2712.245 2753.035 2712.535 2753.080 ;
        RECT 2713.150 2753.020 2713.470 2753.080 ;
        RECT 2712.230 2718.200 2712.550 2718.260 ;
        RECT 2713.150 2718.200 2713.470 2718.260 ;
        RECT 2712.230 2718.060 2713.470 2718.200 ;
        RECT 2712.230 2718.000 2712.550 2718.060 ;
        RECT 2713.150 2718.000 2713.470 2718.060 ;
        RECT 2712.230 2670.260 2712.550 2670.320 ;
        RECT 2713.150 2670.260 2713.470 2670.320 ;
        RECT 2712.230 2670.120 2713.470 2670.260 ;
        RECT 2712.230 2670.060 2712.550 2670.120 ;
        RECT 2713.150 2670.060 2713.470 2670.120 ;
        RECT 2713.150 2622.120 2713.470 2622.380 ;
        RECT 2713.240 2621.980 2713.380 2622.120 ;
        RECT 2713.610 2621.980 2713.930 2622.040 ;
        RECT 2713.240 2621.840 2713.930 2621.980 ;
        RECT 2713.610 2621.780 2713.930 2621.840 ;
        RECT 2712.690 2560.100 2713.010 2560.160 ;
        RECT 2714.070 2560.100 2714.390 2560.160 ;
        RECT 2712.690 2559.960 2714.390 2560.100 ;
        RECT 2712.690 2559.900 2713.010 2559.960 ;
        RECT 2714.070 2559.900 2714.390 2559.960 ;
        RECT 2713.150 2511.820 2713.470 2511.880 ;
        RECT 2714.070 2511.820 2714.390 2511.880 ;
        RECT 2713.150 2511.680 2714.390 2511.820 ;
        RECT 2713.150 2511.620 2713.470 2511.680 ;
        RECT 2714.070 2511.620 2714.390 2511.680 ;
        RECT 2712.690 2463.200 2713.010 2463.260 ;
        RECT 2712.495 2463.060 2713.010 2463.200 ;
        RECT 2712.690 2463.000 2713.010 2463.060 ;
        RECT 2712.690 2428.860 2713.010 2428.920 ;
        RECT 2712.495 2428.720 2713.010 2428.860 ;
        RECT 2712.690 2428.660 2713.010 2428.720 ;
        RECT 2712.230 2380.580 2712.550 2380.640 ;
        RECT 2713.150 2380.580 2713.470 2380.640 ;
        RECT 2712.230 2380.440 2713.470 2380.580 ;
        RECT 2712.230 2380.380 2712.550 2380.440 ;
        RECT 2713.150 2380.380 2713.470 2380.440 ;
        RECT 2712.690 2366.640 2713.010 2366.700 ;
        RECT 2712.495 2366.500 2713.010 2366.640 ;
        RECT 2712.690 2366.440 2713.010 2366.500 ;
        RECT 2712.690 2331.960 2713.010 2332.020 ;
        RECT 2712.495 2331.820 2713.010 2331.960 ;
        RECT 2712.690 2331.760 2713.010 2331.820 ;
        RECT 2711.770 2235.540 2712.090 2235.800 ;
        RECT 2711.860 2235.400 2712.000 2235.540 ;
        RECT 2712.230 2235.400 2712.550 2235.460 ;
        RECT 2711.860 2235.260 2712.550 2235.400 ;
        RECT 2712.230 2235.200 2712.550 2235.260 ;
        RECT 2712.690 2173.520 2713.010 2173.580 ;
        RECT 2712.495 2173.380 2713.010 2173.520 ;
        RECT 2712.690 2173.320 2713.010 2173.380 ;
        RECT 2712.690 2138.840 2713.010 2138.900 ;
        RECT 2712.495 2138.700 2713.010 2138.840 ;
        RECT 2712.690 2138.640 2713.010 2138.700 ;
        RECT 1912.750 2122.180 1913.070 2122.240 ;
        RECT 2713.150 2122.180 2713.470 2122.240 ;
        RECT 1912.750 2122.040 2713.470 2122.180 ;
        RECT 1912.750 2121.980 1913.070 2122.040 ;
        RECT 2713.150 2121.980 2713.470 2122.040 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2712.720 3470.420 2712.980 3470.680 ;
        RECT 2713.640 3470.420 2713.900 3470.680 ;
        RECT 2712.720 3463.620 2712.980 3463.880 ;
        RECT 2713.640 3463.620 2713.900 3463.880 ;
        RECT 2711.800 3415.340 2712.060 3415.600 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2712.720 3042.700 2712.980 3042.960 ;
        RECT 2713.640 3008.360 2713.900 3008.620 ;
        RECT 2713.640 2994.420 2713.900 2994.680 ;
        RECT 2714.100 2946.480 2714.360 2946.740 ;
        RECT 2714.100 2912.140 2714.360 2912.400 ;
        RECT 2713.640 2911.460 2713.900 2911.720 ;
        RECT 2712.260 2815.580 2712.520 2815.840 ;
        RECT 2712.260 2814.900 2712.520 2815.160 ;
        RECT 2712.260 2800.960 2712.520 2801.220 ;
        RECT 2713.180 2753.020 2713.440 2753.280 ;
        RECT 2712.260 2718.000 2712.520 2718.260 ;
        RECT 2713.180 2718.000 2713.440 2718.260 ;
        RECT 2712.260 2670.060 2712.520 2670.320 ;
        RECT 2713.180 2670.060 2713.440 2670.320 ;
        RECT 2713.180 2622.120 2713.440 2622.380 ;
        RECT 2713.640 2621.780 2713.900 2622.040 ;
        RECT 2712.720 2559.900 2712.980 2560.160 ;
        RECT 2714.100 2559.900 2714.360 2560.160 ;
        RECT 2713.180 2511.620 2713.440 2511.880 ;
        RECT 2714.100 2511.620 2714.360 2511.880 ;
        RECT 2712.720 2463.000 2712.980 2463.260 ;
        RECT 2712.720 2428.660 2712.980 2428.920 ;
        RECT 2712.260 2380.380 2712.520 2380.640 ;
        RECT 2713.180 2380.380 2713.440 2380.640 ;
        RECT 2712.720 2366.440 2712.980 2366.700 ;
        RECT 2712.720 2331.760 2712.980 2332.020 ;
        RECT 2711.800 2235.540 2712.060 2235.800 ;
        RECT 2712.260 2235.200 2712.520 2235.460 ;
        RECT 2712.720 2173.320 2712.980 2173.580 ;
        RECT 2712.720 2138.640 2712.980 2138.900 ;
        RECT 1912.780 2121.980 1913.040 2122.240 ;
        RECT 2713.180 2121.980 2713.440 2122.240 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3470.710 2713.840 3491.130 ;
        RECT 2712.720 3470.390 2712.980 3470.710 ;
        RECT 2713.640 3470.390 2713.900 3470.710 ;
        RECT 2712.780 3463.910 2712.920 3470.390 ;
        RECT 2712.720 3463.590 2712.980 3463.910 ;
        RECT 2713.640 3463.590 2713.900 3463.910 ;
        RECT 2713.700 3416.165 2713.840 3463.590 ;
        RECT 2711.790 3415.795 2712.070 3416.165 ;
        RECT 2713.630 3415.795 2713.910 3416.165 ;
        RECT 2711.860 3415.630 2712.000 3415.795 ;
        RECT 2711.800 3415.310 2712.060 3415.630 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3056.330 2712.460 3056.610 ;
        RECT 2712.320 3056.190 2712.920 3056.330 ;
        RECT 2712.780 3042.990 2712.920 3056.190 ;
        RECT 2712.720 3042.670 2712.980 3042.990 ;
        RECT 2713.640 3008.330 2713.900 3008.650 ;
        RECT 2713.700 2994.710 2713.840 3008.330 ;
        RECT 2713.640 2994.390 2713.900 2994.710 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.250 2712.460 2814.870 ;
        RECT 2712.260 2800.930 2712.520 2801.250 ;
        RECT 2713.180 2752.990 2713.440 2753.310 ;
        RECT 2713.240 2718.290 2713.380 2752.990 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2713.180 2717.970 2713.440 2718.290 ;
        RECT 2712.320 2670.350 2712.460 2717.970 ;
        RECT 2712.260 2670.030 2712.520 2670.350 ;
        RECT 2713.180 2670.030 2713.440 2670.350 ;
        RECT 2713.240 2622.410 2713.380 2670.030 ;
        RECT 2713.180 2622.090 2713.440 2622.410 ;
        RECT 2713.640 2621.750 2713.900 2622.070 ;
        RECT 2713.700 2608.325 2713.840 2621.750 ;
        RECT 2712.710 2607.955 2712.990 2608.325 ;
        RECT 2713.630 2607.955 2713.910 2608.325 ;
        RECT 2712.780 2560.190 2712.920 2607.955 ;
        RECT 2712.720 2559.870 2712.980 2560.190 ;
        RECT 2714.100 2559.870 2714.360 2560.190 ;
        RECT 2714.160 2511.910 2714.300 2559.870 ;
        RECT 2713.180 2511.765 2713.440 2511.910 ;
        RECT 2711.790 2511.395 2712.070 2511.765 ;
        RECT 2713.170 2511.395 2713.450 2511.765 ;
        RECT 2714.100 2511.590 2714.360 2511.910 ;
        RECT 2711.860 2463.485 2712.000 2511.395 ;
        RECT 2711.790 2463.115 2712.070 2463.485 ;
        RECT 2712.710 2463.115 2712.990 2463.485 ;
        RECT 2712.720 2462.970 2712.980 2463.115 ;
        RECT 2712.720 2428.630 2712.980 2428.950 ;
        RECT 2712.780 2415.090 2712.920 2428.630 ;
        RECT 2712.780 2414.950 2713.380 2415.090 ;
        RECT 2713.240 2380.670 2713.380 2414.950 ;
        RECT 2712.260 2380.410 2712.520 2380.670 ;
        RECT 2712.260 2380.350 2712.920 2380.410 ;
        RECT 2713.180 2380.350 2713.440 2380.670 ;
        RECT 2712.320 2380.270 2712.920 2380.350 ;
        RECT 2712.780 2366.730 2712.920 2380.270 ;
        RECT 2712.720 2366.410 2712.980 2366.730 ;
        RECT 2712.720 2331.730 2712.980 2332.050 ;
        RECT 2712.780 2318.530 2712.920 2331.730 ;
        RECT 2712.780 2318.390 2713.380 2318.530 ;
        RECT 2713.240 2270.365 2713.380 2318.390 ;
        RECT 2711.790 2269.995 2712.070 2270.365 ;
        RECT 2713.170 2269.995 2713.450 2270.365 ;
        RECT 2711.860 2235.830 2712.000 2269.995 ;
        RECT 2711.800 2235.510 2712.060 2235.830 ;
        RECT 2712.260 2235.170 2712.520 2235.490 ;
        RECT 2712.320 2187.290 2712.460 2235.170 ;
        RECT 2712.320 2187.150 2712.920 2187.290 ;
        RECT 2712.780 2173.610 2712.920 2187.150 ;
        RECT 2712.720 2173.290 2712.980 2173.610 ;
        RECT 2712.720 2138.610 2712.980 2138.930 ;
        RECT 2712.780 2125.410 2712.920 2138.610 ;
        RECT 2712.780 2125.270 2713.380 2125.410 ;
        RECT 2713.240 2122.270 2713.380 2125.270 ;
        RECT 1912.780 2121.950 1913.040 2122.270 ;
        RECT 2713.180 2121.950 2713.440 2122.270 ;
        RECT 1912.840 2112.185 1912.980 2121.950 ;
        RECT 1912.840 2111.740 1913.190 2112.185 ;
        RECT 1912.910 2108.185 1913.190 2111.740 ;
      LAYER via2 ;
        RECT 2711.790 3415.840 2712.070 3416.120 ;
        RECT 2713.630 3415.840 2713.910 3416.120 ;
        RECT 2712.710 2608.000 2712.990 2608.280 ;
        RECT 2713.630 2608.000 2713.910 2608.280 ;
        RECT 2711.790 2511.440 2712.070 2511.720 ;
        RECT 2713.170 2511.440 2713.450 2511.720 ;
        RECT 2711.790 2463.160 2712.070 2463.440 ;
        RECT 2712.710 2463.160 2712.990 2463.440 ;
        RECT 2711.790 2270.040 2712.070 2270.320 ;
        RECT 2713.170 2270.040 2713.450 2270.320 ;
      LAYER met3 ;
        RECT 2711.765 3416.130 2712.095 3416.145 ;
        RECT 2713.605 3416.130 2713.935 3416.145 ;
        RECT 2711.765 3415.830 2713.935 3416.130 ;
        RECT 2711.765 3415.815 2712.095 3415.830 ;
        RECT 2713.605 3415.815 2713.935 3415.830 ;
        RECT 2712.685 2608.290 2713.015 2608.305 ;
        RECT 2713.605 2608.290 2713.935 2608.305 ;
        RECT 2712.685 2607.990 2713.935 2608.290 ;
        RECT 2712.685 2607.975 2713.015 2607.990 ;
        RECT 2713.605 2607.975 2713.935 2607.990 ;
        RECT 2711.765 2511.730 2712.095 2511.745 ;
        RECT 2713.145 2511.730 2713.475 2511.745 ;
        RECT 2711.765 2511.430 2713.475 2511.730 ;
        RECT 2711.765 2511.415 2712.095 2511.430 ;
        RECT 2713.145 2511.415 2713.475 2511.430 ;
        RECT 2711.765 2463.450 2712.095 2463.465 ;
        RECT 2712.685 2463.450 2713.015 2463.465 ;
        RECT 2711.765 2463.150 2713.015 2463.450 ;
        RECT 2711.765 2463.135 2712.095 2463.150 ;
        RECT 2712.685 2463.135 2713.015 2463.150 ;
        RECT 2711.765 2270.330 2712.095 2270.345 ;
        RECT 2713.145 2270.330 2713.475 2270.345 ;
        RECT 2711.765 2270.030 2713.475 2270.330 ;
        RECT 2711.765 2270.015 2712.095 2270.030 ;
        RECT 2713.145 2270.015 2713.475 2270.030 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2387.545 2898.245 2387.715 2946.355 ;
        RECT 2388.005 2815.285 2388.175 2849.455 ;
      LAYER mcon ;
        RECT 2387.545 2946.185 2387.715 2946.355 ;
        RECT 2388.005 2849.285 2388.175 2849.455 ;
      LAYER met1 ;
        RECT 2387.470 3464.160 2387.790 3464.220 ;
        RECT 2392.990 3464.160 2393.310 3464.220 ;
        RECT 2387.470 3464.020 2393.310 3464.160 ;
        RECT 2387.470 3463.960 2387.790 3464.020 ;
        RECT 2392.990 3463.960 2393.310 3464.020 ;
        RECT 2387.470 3367.600 2387.790 3367.660 ;
        RECT 2388.390 3367.600 2388.710 3367.660 ;
        RECT 2387.470 3367.460 2388.710 3367.600 ;
        RECT 2387.470 3367.400 2387.790 3367.460 ;
        RECT 2388.390 3367.400 2388.710 3367.460 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 2387.470 3077.580 2387.790 3077.640 ;
        RECT 2388.390 3077.580 2388.710 3077.640 ;
        RECT 2387.470 3077.440 2388.710 3077.580 ;
        RECT 2387.470 3077.380 2387.790 3077.440 ;
        RECT 2388.390 3077.380 2388.710 3077.440 ;
        RECT 2387.470 2981.020 2387.790 2981.080 ;
        RECT 2388.390 2981.020 2388.710 2981.080 ;
        RECT 2387.470 2980.880 2388.710 2981.020 ;
        RECT 2387.470 2980.820 2387.790 2980.880 ;
        RECT 2388.390 2980.820 2388.710 2980.880 ;
        RECT 2387.485 2946.340 2387.775 2946.385 ;
        RECT 2387.930 2946.340 2388.250 2946.400 ;
        RECT 2387.485 2946.200 2388.250 2946.340 ;
        RECT 2387.485 2946.155 2387.775 2946.200 ;
        RECT 2387.930 2946.140 2388.250 2946.200 ;
        RECT 2387.470 2898.400 2387.790 2898.460 ;
        RECT 2387.275 2898.260 2387.790 2898.400 ;
        RECT 2387.470 2898.200 2387.790 2898.260 ;
        RECT 2387.930 2849.440 2388.250 2849.500 ;
        RECT 2387.735 2849.300 2388.250 2849.440 ;
        RECT 2387.930 2849.240 2388.250 2849.300 ;
        RECT 2387.945 2815.440 2388.235 2815.485 ;
        RECT 2388.850 2815.440 2389.170 2815.500 ;
        RECT 2387.945 2815.300 2389.170 2815.440 ;
        RECT 2387.945 2815.255 2388.235 2815.300 ;
        RECT 2388.850 2815.240 2389.170 2815.300 ;
        RECT 2387.930 2753.220 2388.250 2753.280 ;
        RECT 2389.310 2753.220 2389.630 2753.280 ;
        RECT 2387.930 2753.080 2389.630 2753.220 ;
        RECT 2387.930 2753.020 2388.250 2753.080 ;
        RECT 2389.310 2753.020 2389.630 2753.080 ;
        RECT 2389.310 2719.220 2389.630 2719.280 ;
        RECT 2388.940 2719.080 2389.630 2719.220 ;
        RECT 2388.940 2718.600 2389.080 2719.080 ;
        RECT 2389.310 2719.020 2389.630 2719.080 ;
        RECT 2388.850 2718.340 2389.170 2718.600 ;
        RECT 2387.930 2656.660 2388.250 2656.720 ;
        RECT 2389.310 2656.660 2389.630 2656.720 ;
        RECT 2387.930 2656.520 2389.630 2656.660 ;
        RECT 2387.930 2656.460 2388.250 2656.520 ;
        RECT 2389.310 2656.460 2389.630 2656.520 ;
        RECT 2389.310 2622.660 2389.630 2622.720 ;
        RECT 2388.940 2622.520 2389.630 2622.660 ;
        RECT 2388.940 2622.040 2389.080 2622.520 ;
        RECT 2389.310 2622.460 2389.630 2622.520 ;
        RECT 2388.850 2621.780 2389.170 2622.040 ;
        RECT 2387.930 2560.100 2388.250 2560.160 ;
        RECT 2389.310 2560.100 2389.630 2560.160 ;
        RECT 2387.930 2559.960 2389.630 2560.100 ;
        RECT 2387.930 2559.900 2388.250 2559.960 ;
        RECT 2389.310 2559.900 2389.630 2559.960 ;
        RECT 2388.390 2511.820 2388.710 2511.880 ;
        RECT 2389.310 2511.820 2389.630 2511.880 ;
        RECT 2388.390 2511.680 2389.630 2511.820 ;
        RECT 2388.390 2511.620 2388.710 2511.680 ;
        RECT 2389.310 2511.620 2389.630 2511.680 ;
        RECT 2387.470 2401.320 2387.790 2401.380 ;
        RECT 2388.390 2401.320 2388.710 2401.380 ;
        RECT 2387.470 2401.180 2388.710 2401.320 ;
        RECT 2387.470 2401.120 2387.790 2401.180 ;
        RECT 2388.390 2401.120 2388.710 2401.180 ;
        RECT 2387.470 2304.760 2387.790 2304.820 ;
        RECT 2388.390 2304.760 2388.710 2304.820 ;
        RECT 2387.470 2304.620 2388.710 2304.760 ;
        RECT 2387.470 2304.560 2387.790 2304.620 ;
        RECT 2388.390 2304.560 2388.710 2304.620 ;
        RECT 2387.470 2208.200 2387.790 2208.260 ;
        RECT 2388.390 2208.200 2388.710 2208.260 ;
        RECT 2387.470 2208.060 2388.710 2208.200 ;
        RECT 2387.470 2208.000 2387.790 2208.060 ;
        RECT 2388.390 2208.000 2388.710 2208.060 ;
        RECT 1736.110 2123.200 1736.430 2123.260 ;
        RECT 2388.390 2123.200 2388.710 2123.260 ;
        RECT 1736.110 2123.060 2388.710 2123.200 ;
        RECT 1736.110 2123.000 1736.430 2123.060 ;
        RECT 2388.390 2123.000 2388.710 2123.060 ;
      LAYER via ;
        RECT 2387.500 3463.960 2387.760 3464.220 ;
        RECT 2393.020 3463.960 2393.280 3464.220 ;
        RECT 2387.500 3367.400 2387.760 3367.660 ;
        RECT 2388.420 3367.400 2388.680 3367.660 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 2387.500 3077.380 2387.760 3077.640 ;
        RECT 2388.420 3077.380 2388.680 3077.640 ;
        RECT 2387.500 2980.820 2387.760 2981.080 ;
        RECT 2388.420 2980.820 2388.680 2981.080 ;
        RECT 2387.960 2946.140 2388.220 2946.400 ;
        RECT 2387.500 2898.200 2387.760 2898.460 ;
        RECT 2387.960 2849.240 2388.220 2849.500 ;
        RECT 2388.880 2815.240 2389.140 2815.500 ;
        RECT 2387.960 2753.020 2388.220 2753.280 ;
        RECT 2389.340 2753.020 2389.600 2753.280 ;
        RECT 2389.340 2719.020 2389.600 2719.280 ;
        RECT 2388.880 2718.340 2389.140 2718.600 ;
        RECT 2387.960 2656.460 2388.220 2656.720 ;
        RECT 2389.340 2656.460 2389.600 2656.720 ;
        RECT 2389.340 2622.460 2389.600 2622.720 ;
        RECT 2388.880 2621.780 2389.140 2622.040 ;
        RECT 2387.960 2559.900 2388.220 2560.160 ;
        RECT 2389.340 2559.900 2389.600 2560.160 ;
        RECT 2388.420 2511.620 2388.680 2511.880 ;
        RECT 2389.340 2511.620 2389.600 2511.880 ;
        RECT 2387.500 2401.120 2387.760 2401.380 ;
        RECT 2388.420 2401.120 2388.680 2401.380 ;
        RECT 2387.500 2304.560 2387.760 2304.820 ;
        RECT 2388.420 2304.560 2388.680 2304.820 ;
        RECT 2387.500 2208.000 2387.760 2208.260 ;
        RECT 2388.420 2208.000 2388.680 2208.260 ;
        RECT 1736.140 2123.000 1736.400 2123.260 ;
        RECT 2388.420 2123.000 2388.680 2123.260 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3464.250 2393.220 3517.230 ;
        RECT 2387.500 3463.930 2387.760 3464.250 ;
        RECT 2393.020 3463.930 2393.280 3464.250 ;
        RECT 2387.560 3415.370 2387.700 3463.930 ;
        RECT 2387.560 3415.230 2388.620 3415.370 ;
        RECT 2388.480 3367.690 2388.620 3415.230 ;
        RECT 2387.500 3367.370 2387.760 3367.690 ;
        RECT 2388.420 3367.370 2388.680 3367.690 ;
        RECT 2387.560 3318.810 2387.700 3367.370 ;
        RECT 2387.560 3318.670 2388.620 3318.810 ;
        RECT 2388.480 3270.790 2388.620 3318.670 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 2981.110 2388.620 3028.990 ;
        RECT 2387.500 2980.850 2387.760 2981.110 ;
        RECT 2387.500 2980.790 2388.160 2980.850 ;
        RECT 2388.420 2980.790 2388.680 2981.110 ;
        RECT 2387.560 2980.710 2388.160 2980.790 ;
        RECT 2388.020 2980.170 2388.160 2980.710 ;
        RECT 2388.020 2980.030 2388.620 2980.170 ;
        RECT 2388.480 2959.770 2388.620 2980.030 ;
        RECT 2388.020 2959.630 2388.620 2959.770 ;
        RECT 2388.020 2946.430 2388.160 2959.630 ;
        RECT 2387.960 2946.110 2388.220 2946.430 ;
        RECT 2387.500 2898.170 2387.760 2898.490 ;
        RECT 2387.560 2863.210 2387.700 2898.170 ;
        RECT 2387.560 2863.070 2388.160 2863.210 ;
        RECT 2388.020 2849.530 2388.160 2863.070 ;
        RECT 2387.960 2849.210 2388.220 2849.530 ;
        RECT 2388.880 2815.210 2389.140 2815.530 ;
        RECT 2388.940 2801.445 2389.080 2815.210 ;
        RECT 2387.950 2801.075 2388.230 2801.445 ;
        RECT 2388.870 2801.075 2389.150 2801.445 ;
        RECT 2388.020 2753.310 2388.160 2801.075 ;
        RECT 2387.960 2752.990 2388.220 2753.310 ;
        RECT 2389.340 2752.990 2389.600 2753.310 ;
        RECT 2389.400 2719.310 2389.540 2752.990 ;
        RECT 2389.340 2718.990 2389.600 2719.310 ;
        RECT 2388.880 2718.310 2389.140 2718.630 ;
        RECT 2388.940 2704.885 2389.080 2718.310 ;
        RECT 2387.950 2704.515 2388.230 2704.885 ;
        RECT 2388.870 2704.515 2389.150 2704.885 ;
        RECT 2388.020 2656.750 2388.160 2704.515 ;
        RECT 2387.960 2656.430 2388.220 2656.750 ;
        RECT 2389.340 2656.430 2389.600 2656.750 ;
        RECT 2389.400 2622.750 2389.540 2656.430 ;
        RECT 2389.340 2622.430 2389.600 2622.750 ;
        RECT 2388.880 2621.750 2389.140 2622.070 ;
        RECT 2388.940 2608.325 2389.080 2621.750 ;
        RECT 2387.950 2607.955 2388.230 2608.325 ;
        RECT 2388.870 2607.955 2389.150 2608.325 ;
        RECT 2388.020 2560.190 2388.160 2607.955 ;
        RECT 2387.960 2559.870 2388.220 2560.190 ;
        RECT 2389.340 2559.870 2389.600 2560.190 ;
        RECT 2389.400 2511.910 2389.540 2559.870 ;
        RECT 2388.420 2511.765 2388.680 2511.910 ;
        RECT 2387.030 2511.395 2387.310 2511.765 ;
        RECT 2388.410 2511.395 2388.690 2511.765 ;
        RECT 2389.340 2511.590 2389.600 2511.910 ;
        RECT 2387.100 2463.485 2387.240 2511.395 ;
        RECT 2387.030 2463.115 2387.310 2463.485 ;
        RECT 2387.950 2463.115 2388.230 2463.485 ;
        RECT 2388.020 2449.770 2388.160 2463.115 ;
        RECT 2388.020 2449.630 2388.620 2449.770 ;
        RECT 2388.480 2401.410 2388.620 2449.630 ;
        RECT 2387.500 2401.090 2387.760 2401.410 ;
        RECT 2388.420 2401.090 2388.680 2401.410 ;
        RECT 2387.560 2400.810 2387.700 2401.090 ;
        RECT 2387.560 2400.670 2388.160 2400.810 ;
        RECT 2388.020 2353.210 2388.160 2400.670 ;
        RECT 2388.020 2353.070 2388.620 2353.210 ;
        RECT 2388.480 2304.850 2388.620 2353.070 ;
        RECT 2387.500 2304.530 2387.760 2304.850 ;
        RECT 2388.420 2304.530 2388.680 2304.850 ;
        RECT 2387.560 2304.250 2387.700 2304.530 ;
        RECT 2387.560 2304.110 2388.160 2304.250 ;
        RECT 2388.020 2256.650 2388.160 2304.110 ;
        RECT 2388.020 2256.510 2388.620 2256.650 ;
        RECT 2388.480 2208.290 2388.620 2256.510 ;
        RECT 2387.500 2207.970 2387.760 2208.290 ;
        RECT 2388.420 2207.970 2388.680 2208.290 ;
        RECT 2387.560 2207.690 2387.700 2207.970 ;
        RECT 2387.560 2207.550 2388.160 2207.690 ;
        RECT 2388.020 2160.090 2388.160 2207.550 ;
        RECT 2388.020 2159.950 2388.620 2160.090 ;
        RECT 2388.480 2123.290 2388.620 2159.950 ;
        RECT 1736.140 2122.970 1736.400 2123.290 ;
        RECT 2388.420 2122.970 2388.680 2123.290 ;
        RECT 1736.200 2112.185 1736.340 2122.970 ;
        RECT 1736.200 2111.740 1736.550 2112.185 ;
        RECT 1736.270 2108.185 1736.550 2111.740 ;
      LAYER via2 ;
        RECT 2387.950 2801.120 2388.230 2801.400 ;
        RECT 2388.870 2801.120 2389.150 2801.400 ;
        RECT 2387.950 2704.560 2388.230 2704.840 ;
        RECT 2388.870 2704.560 2389.150 2704.840 ;
        RECT 2387.950 2608.000 2388.230 2608.280 ;
        RECT 2388.870 2608.000 2389.150 2608.280 ;
        RECT 2387.030 2511.440 2387.310 2511.720 ;
        RECT 2388.410 2511.440 2388.690 2511.720 ;
        RECT 2387.030 2463.160 2387.310 2463.440 ;
        RECT 2387.950 2463.160 2388.230 2463.440 ;
      LAYER met3 ;
        RECT 2387.925 2801.410 2388.255 2801.425 ;
        RECT 2388.845 2801.410 2389.175 2801.425 ;
        RECT 2387.925 2801.110 2389.175 2801.410 ;
        RECT 2387.925 2801.095 2388.255 2801.110 ;
        RECT 2388.845 2801.095 2389.175 2801.110 ;
        RECT 2387.925 2704.850 2388.255 2704.865 ;
        RECT 2388.845 2704.850 2389.175 2704.865 ;
        RECT 2387.925 2704.550 2389.175 2704.850 ;
        RECT 2387.925 2704.535 2388.255 2704.550 ;
        RECT 2388.845 2704.535 2389.175 2704.550 ;
        RECT 2387.925 2608.290 2388.255 2608.305 ;
        RECT 2388.845 2608.290 2389.175 2608.305 ;
        RECT 2387.925 2607.990 2389.175 2608.290 ;
        RECT 2387.925 2607.975 2388.255 2607.990 ;
        RECT 2388.845 2607.975 2389.175 2607.990 ;
        RECT 2387.005 2511.730 2387.335 2511.745 ;
        RECT 2388.385 2511.730 2388.715 2511.745 ;
        RECT 2387.005 2511.430 2388.715 2511.730 ;
        RECT 2387.005 2511.415 2387.335 2511.430 ;
        RECT 2388.385 2511.415 2388.715 2511.430 ;
        RECT 2387.005 2463.450 2387.335 2463.465 ;
        RECT 2387.925 2463.450 2388.255 2463.465 ;
        RECT 2387.005 2463.150 2388.255 2463.450 ;
        RECT 2387.005 2463.135 2387.335 2463.150 ;
        RECT 2387.925 2463.135 2388.255 2463.150 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2063.245 3416.065 2063.415 3463.835 ;
        RECT 2065.085 3332.765 2065.255 3415.555 ;
        RECT 2064.165 3008.405 2064.335 3042.915 ;
        RECT 2065.085 2946.525 2065.255 2994.635 ;
        RECT 2063.705 2753.065 2063.875 2801.175 ;
        RECT 2064.165 2428.705 2064.335 2463.215 ;
        RECT 2064.165 2331.805 2064.335 2366.655 ;
        RECT 2064.165 2138.685 2064.335 2173.535 ;
      LAYER mcon ;
        RECT 2063.245 3463.665 2063.415 3463.835 ;
        RECT 2065.085 3415.385 2065.255 3415.555 ;
        RECT 2064.165 3042.745 2064.335 3042.915 ;
        RECT 2065.085 2994.465 2065.255 2994.635 ;
        RECT 2063.705 2801.005 2063.875 2801.175 ;
        RECT 2064.165 2463.045 2064.335 2463.215 ;
        RECT 2064.165 2366.485 2064.335 2366.655 ;
        RECT 2064.165 2173.365 2064.335 2173.535 ;
      LAYER met1 ;
        RECT 2065.010 3491.360 2065.330 3491.420 ;
        RECT 2068.690 3491.360 2069.010 3491.420 ;
        RECT 2065.010 3491.220 2069.010 3491.360 ;
        RECT 2065.010 3491.160 2065.330 3491.220 ;
        RECT 2068.690 3491.160 2069.010 3491.220 ;
        RECT 2064.090 3470.620 2064.410 3470.680 ;
        RECT 2065.010 3470.620 2065.330 3470.680 ;
        RECT 2064.090 3470.480 2065.330 3470.620 ;
        RECT 2064.090 3470.420 2064.410 3470.480 ;
        RECT 2065.010 3470.420 2065.330 3470.480 ;
        RECT 2063.185 3463.820 2063.475 3463.865 ;
        RECT 2064.090 3463.820 2064.410 3463.880 ;
        RECT 2063.185 3463.680 2064.410 3463.820 ;
        RECT 2063.185 3463.635 2063.475 3463.680 ;
        RECT 2064.090 3463.620 2064.410 3463.680 ;
        RECT 2063.170 3416.220 2063.490 3416.280 ;
        RECT 2063.170 3416.080 2063.685 3416.220 ;
        RECT 2063.170 3416.020 2063.490 3416.080 ;
        RECT 2063.170 3415.540 2063.490 3415.600 ;
        RECT 2065.025 3415.540 2065.315 3415.585 ;
        RECT 2063.170 3415.400 2065.315 3415.540 ;
        RECT 2063.170 3415.340 2063.490 3415.400 ;
        RECT 2065.025 3415.355 2065.315 3415.400 ;
        RECT 2065.025 3332.920 2065.315 3332.965 ;
        RECT 2065.470 3332.920 2065.790 3332.980 ;
        RECT 2065.025 3332.780 2065.790 3332.920 ;
        RECT 2065.025 3332.735 2065.315 3332.780 ;
        RECT 2065.470 3332.720 2065.790 3332.780 ;
        RECT 2064.090 3236.360 2064.410 3236.420 ;
        RECT 2064.550 3236.360 2064.870 3236.420 ;
        RECT 2064.090 3236.220 2064.870 3236.360 ;
        RECT 2064.090 3236.160 2064.410 3236.220 ;
        RECT 2064.550 3236.160 2064.870 3236.220 ;
        RECT 2064.090 3202.020 2064.410 3202.080 ;
        RECT 2064.550 3202.020 2064.870 3202.080 ;
        RECT 2064.090 3201.880 2064.870 3202.020 ;
        RECT 2064.090 3201.820 2064.410 3201.880 ;
        RECT 2064.550 3201.820 2064.870 3201.880 ;
        RECT 2063.630 3153.400 2063.950 3153.460 ;
        RECT 2064.550 3153.400 2064.870 3153.460 ;
        RECT 2063.630 3153.260 2064.870 3153.400 ;
        RECT 2063.630 3153.200 2063.950 3153.260 ;
        RECT 2064.550 3153.200 2064.870 3153.260 ;
        RECT 2063.630 3056.840 2063.950 3056.900 ;
        RECT 2064.550 3056.840 2064.870 3056.900 ;
        RECT 2063.630 3056.700 2064.870 3056.840 ;
        RECT 2063.630 3056.640 2063.950 3056.700 ;
        RECT 2064.550 3056.640 2064.870 3056.700 ;
        RECT 2064.090 3042.900 2064.410 3042.960 ;
        RECT 2063.895 3042.760 2064.410 3042.900 ;
        RECT 2064.090 3042.700 2064.410 3042.760 ;
        RECT 2064.105 3008.560 2064.395 3008.605 ;
        RECT 2065.010 3008.560 2065.330 3008.620 ;
        RECT 2064.105 3008.420 2065.330 3008.560 ;
        RECT 2064.105 3008.375 2064.395 3008.420 ;
        RECT 2065.010 3008.360 2065.330 3008.420 ;
        RECT 2065.010 2994.620 2065.330 2994.680 ;
        RECT 2064.815 2994.480 2065.330 2994.620 ;
        RECT 2065.010 2994.420 2065.330 2994.480 ;
        RECT 2065.025 2946.680 2065.315 2946.725 ;
        RECT 2065.470 2946.680 2065.790 2946.740 ;
        RECT 2065.025 2946.540 2065.790 2946.680 ;
        RECT 2065.025 2946.495 2065.315 2946.540 ;
        RECT 2065.470 2946.480 2065.790 2946.540 ;
        RECT 2065.470 2912.340 2065.790 2912.400 ;
        RECT 2065.100 2912.200 2065.790 2912.340 ;
        RECT 2065.100 2911.720 2065.240 2912.200 ;
        RECT 2065.470 2912.140 2065.790 2912.200 ;
        RECT 2065.010 2911.460 2065.330 2911.720 ;
        RECT 2063.630 2815.580 2063.950 2815.840 ;
        RECT 2063.720 2815.160 2063.860 2815.580 ;
        RECT 2063.630 2814.900 2063.950 2815.160 ;
        RECT 2063.630 2801.160 2063.950 2801.220 ;
        RECT 2063.435 2801.020 2063.950 2801.160 ;
        RECT 2063.630 2800.960 2063.950 2801.020 ;
        RECT 2063.645 2753.220 2063.935 2753.265 ;
        RECT 2064.550 2753.220 2064.870 2753.280 ;
        RECT 2063.645 2753.080 2064.870 2753.220 ;
        RECT 2063.645 2753.035 2063.935 2753.080 ;
        RECT 2064.550 2753.020 2064.870 2753.080 ;
        RECT 2063.630 2718.200 2063.950 2718.260 ;
        RECT 2064.550 2718.200 2064.870 2718.260 ;
        RECT 2063.630 2718.060 2064.870 2718.200 ;
        RECT 2063.630 2718.000 2063.950 2718.060 ;
        RECT 2064.550 2718.000 2064.870 2718.060 ;
        RECT 2063.630 2670.260 2063.950 2670.320 ;
        RECT 2064.550 2670.260 2064.870 2670.320 ;
        RECT 2063.630 2670.120 2064.870 2670.260 ;
        RECT 2063.630 2670.060 2063.950 2670.120 ;
        RECT 2064.550 2670.060 2064.870 2670.120 ;
        RECT 2064.550 2622.120 2064.870 2622.380 ;
        RECT 2064.640 2621.980 2064.780 2622.120 ;
        RECT 2065.010 2621.980 2065.330 2622.040 ;
        RECT 2064.640 2621.840 2065.330 2621.980 ;
        RECT 2065.010 2621.780 2065.330 2621.840 ;
        RECT 2064.090 2560.100 2064.410 2560.160 ;
        RECT 2065.470 2560.100 2065.790 2560.160 ;
        RECT 2064.090 2559.960 2065.790 2560.100 ;
        RECT 2064.090 2559.900 2064.410 2559.960 ;
        RECT 2065.470 2559.900 2065.790 2559.960 ;
        RECT 2064.550 2511.820 2064.870 2511.880 ;
        RECT 2065.470 2511.820 2065.790 2511.880 ;
        RECT 2064.550 2511.680 2065.790 2511.820 ;
        RECT 2064.550 2511.620 2064.870 2511.680 ;
        RECT 2065.470 2511.620 2065.790 2511.680 ;
        RECT 2064.090 2463.200 2064.410 2463.260 ;
        RECT 2063.895 2463.060 2064.410 2463.200 ;
        RECT 2064.090 2463.000 2064.410 2463.060 ;
        RECT 2064.090 2428.860 2064.410 2428.920 ;
        RECT 2063.895 2428.720 2064.410 2428.860 ;
        RECT 2064.090 2428.660 2064.410 2428.720 ;
        RECT 2063.630 2380.580 2063.950 2380.640 ;
        RECT 2064.550 2380.580 2064.870 2380.640 ;
        RECT 2063.630 2380.440 2064.870 2380.580 ;
        RECT 2063.630 2380.380 2063.950 2380.440 ;
        RECT 2064.550 2380.380 2064.870 2380.440 ;
        RECT 2064.090 2366.640 2064.410 2366.700 ;
        RECT 2063.895 2366.500 2064.410 2366.640 ;
        RECT 2064.090 2366.440 2064.410 2366.500 ;
        RECT 2064.090 2331.960 2064.410 2332.020 ;
        RECT 2063.895 2331.820 2064.410 2331.960 ;
        RECT 2064.090 2331.760 2064.410 2331.820 ;
        RECT 2063.170 2235.540 2063.490 2235.800 ;
        RECT 2063.260 2235.400 2063.400 2235.540 ;
        RECT 2063.630 2235.400 2063.950 2235.460 ;
        RECT 2063.260 2235.260 2063.950 2235.400 ;
        RECT 2063.630 2235.200 2063.950 2235.260 ;
        RECT 2064.090 2173.520 2064.410 2173.580 ;
        RECT 2063.895 2173.380 2064.410 2173.520 ;
        RECT 2064.090 2173.320 2064.410 2173.380 ;
        RECT 2064.090 2138.840 2064.410 2138.900 ;
        RECT 2063.895 2138.700 2064.410 2138.840 ;
        RECT 2064.090 2138.640 2064.410 2138.700 ;
        RECT 1559.010 2124.220 1559.330 2124.280 ;
        RECT 2064.550 2124.220 2064.870 2124.280 ;
        RECT 1559.010 2124.080 2064.870 2124.220 ;
        RECT 1559.010 2124.020 1559.330 2124.080 ;
        RECT 2064.550 2124.020 2064.870 2124.080 ;
      LAYER via ;
        RECT 2065.040 3491.160 2065.300 3491.420 ;
        RECT 2068.720 3491.160 2068.980 3491.420 ;
        RECT 2064.120 3470.420 2064.380 3470.680 ;
        RECT 2065.040 3470.420 2065.300 3470.680 ;
        RECT 2064.120 3463.620 2064.380 3463.880 ;
        RECT 2063.200 3416.020 2063.460 3416.280 ;
        RECT 2063.200 3415.340 2063.460 3415.600 ;
        RECT 2065.500 3332.720 2065.760 3332.980 ;
        RECT 2064.120 3236.160 2064.380 3236.420 ;
        RECT 2064.580 3236.160 2064.840 3236.420 ;
        RECT 2064.120 3201.820 2064.380 3202.080 ;
        RECT 2064.580 3201.820 2064.840 3202.080 ;
        RECT 2063.660 3153.200 2063.920 3153.460 ;
        RECT 2064.580 3153.200 2064.840 3153.460 ;
        RECT 2063.660 3056.640 2063.920 3056.900 ;
        RECT 2064.580 3056.640 2064.840 3056.900 ;
        RECT 2064.120 3042.700 2064.380 3042.960 ;
        RECT 2065.040 3008.360 2065.300 3008.620 ;
        RECT 2065.040 2994.420 2065.300 2994.680 ;
        RECT 2065.500 2946.480 2065.760 2946.740 ;
        RECT 2065.500 2912.140 2065.760 2912.400 ;
        RECT 2065.040 2911.460 2065.300 2911.720 ;
        RECT 2063.660 2815.580 2063.920 2815.840 ;
        RECT 2063.660 2814.900 2063.920 2815.160 ;
        RECT 2063.660 2800.960 2063.920 2801.220 ;
        RECT 2064.580 2753.020 2064.840 2753.280 ;
        RECT 2063.660 2718.000 2063.920 2718.260 ;
        RECT 2064.580 2718.000 2064.840 2718.260 ;
        RECT 2063.660 2670.060 2063.920 2670.320 ;
        RECT 2064.580 2670.060 2064.840 2670.320 ;
        RECT 2064.580 2622.120 2064.840 2622.380 ;
        RECT 2065.040 2621.780 2065.300 2622.040 ;
        RECT 2064.120 2559.900 2064.380 2560.160 ;
        RECT 2065.500 2559.900 2065.760 2560.160 ;
        RECT 2064.580 2511.620 2064.840 2511.880 ;
        RECT 2065.500 2511.620 2065.760 2511.880 ;
        RECT 2064.120 2463.000 2064.380 2463.260 ;
        RECT 2064.120 2428.660 2064.380 2428.920 ;
        RECT 2063.660 2380.380 2063.920 2380.640 ;
        RECT 2064.580 2380.380 2064.840 2380.640 ;
        RECT 2064.120 2366.440 2064.380 2366.700 ;
        RECT 2064.120 2331.760 2064.380 2332.020 ;
        RECT 2063.200 2235.540 2063.460 2235.800 ;
        RECT 2063.660 2235.200 2063.920 2235.460 ;
        RECT 2064.120 2173.320 2064.380 2173.580 ;
        RECT 2064.120 2138.640 2064.380 2138.900 ;
        RECT 1559.040 2124.020 1559.300 2124.280 ;
        RECT 2064.580 2124.020 2064.840 2124.280 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3470.710 2065.240 3491.130 ;
        RECT 2064.120 3470.390 2064.380 3470.710 ;
        RECT 2065.040 3470.390 2065.300 3470.710 ;
        RECT 2064.180 3463.910 2064.320 3470.390 ;
        RECT 2064.120 3463.590 2064.380 3463.910 ;
        RECT 2063.200 3415.990 2063.460 3416.310 ;
        RECT 2063.260 3415.630 2063.400 3415.990 ;
        RECT 2063.200 3415.310 2063.460 3415.630 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3056.330 2063.860 3056.610 ;
        RECT 2063.720 3056.190 2064.320 3056.330 ;
        RECT 2064.180 3042.990 2064.320 3056.190 ;
        RECT 2064.120 3042.670 2064.380 3042.990 ;
        RECT 2065.040 3008.330 2065.300 3008.650 ;
        RECT 2065.100 2994.710 2065.240 3008.330 ;
        RECT 2065.040 2994.390 2065.300 2994.710 ;
        RECT 2065.500 2946.450 2065.760 2946.770 ;
        RECT 2065.560 2912.430 2065.700 2946.450 ;
        RECT 2065.500 2912.110 2065.760 2912.430 ;
        RECT 2065.040 2911.430 2065.300 2911.750 ;
        RECT 2065.100 2863.210 2065.240 2911.430 ;
        RECT 2064.180 2863.070 2065.240 2863.210 ;
        RECT 2064.180 2849.610 2064.320 2863.070 ;
        RECT 2063.720 2849.470 2064.320 2849.610 ;
        RECT 2063.720 2815.870 2063.860 2849.470 ;
        RECT 2063.660 2815.550 2063.920 2815.870 ;
        RECT 2063.660 2814.870 2063.920 2815.190 ;
        RECT 2063.720 2801.250 2063.860 2814.870 ;
        RECT 2063.660 2800.930 2063.920 2801.250 ;
        RECT 2064.580 2752.990 2064.840 2753.310 ;
        RECT 2064.640 2718.290 2064.780 2752.990 ;
        RECT 2063.660 2717.970 2063.920 2718.290 ;
        RECT 2064.580 2717.970 2064.840 2718.290 ;
        RECT 2063.720 2670.350 2063.860 2717.970 ;
        RECT 2063.660 2670.030 2063.920 2670.350 ;
        RECT 2064.580 2670.030 2064.840 2670.350 ;
        RECT 2064.640 2622.410 2064.780 2670.030 ;
        RECT 2064.580 2622.090 2064.840 2622.410 ;
        RECT 2065.040 2621.750 2065.300 2622.070 ;
        RECT 2065.100 2608.325 2065.240 2621.750 ;
        RECT 2064.110 2607.955 2064.390 2608.325 ;
        RECT 2065.030 2607.955 2065.310 2608.325 ;
        RECT 2064.180 2560.190 2064.320 2607.955 ;
        RECT 2064.120 2559.870 2064.380 2560.190 ;
        RECT 2065.500 2559.870 2065.760 2560.190 ;
        RECT 2065.560 2511.910 2065.700 2559.870 ;
        RECT 2064.580 2511.765 2064.840 2511.910 ;
        RECT 2063.190 2511.395 2063.470 2511.765 ;
        RECT 2064.570 2511.395 2064.850 2511.765 ;
        RECT 2065.500 2511.590 2065.760 2511.910 ;
        RECT 2063.260 2463.485 2063.400 2511.395 ;
        RECT 2063.190 2463.115 2063.470 2463.485 ;
        RECT 2064.110 2463.115 2064.390 2463.485 ;
        RECT 2064.120 2462.970 2064.380 2463.115 ;
        RECT 2064.120 2428.630 2064.380 2428.950 ;
        RECT 2064.180 2415.090 2064.320 2428.630 ;
        RECT 2064.180 2414.950 2064.780 2415.090 ;
        RECT 2064.640 2380.670 2064.780 2414.950 ;
        RECT 2063.660 2380.410 2063.920 2380.670 ;
        RECT 2063.660 2380.350 2064.320 2380.410 ;
        RECT 2064.580 2380.350 2064.840 2380.670 ;
        RECT 2063.720 2380.270 2064.320 2380.350 ;
        RECT 2064.180 2366.730 2064.320 2380.270 ;
        RECT 2064.120 2366.410 2064.380 2366.730 ;
        RECT 2064.120 2331.730 2064.380 2332.050 ;
        RECT 2064.180 2318.530 2064.320 2331.730 ;
        RECT 2064.180 2318.390 2064.780 2318.530 ;
        RECT 2064.640 2270.365 2064.780 2318.390 ;
        RECT 2063.190 2269.995 2063.470 2270.365 ;
        RECT 2064.570 2269.995 2064.850 2270.365 ;
        RECT 2063.260 2235.830 2063.400 2269.995 ;
        RECT 2063.200 2235.510 2063.460 2235.830 ;
        RECT 2063.660 2235.170 2063.920 2235.490 ;
        RECT 2063.720 2187.290 2063.860 2235.170 ;
        RECT 2063.720 2187.150 2064.320 2187.290 ;
        RECT 2064.180 2173.610 2064.320 2187.150 ;
        RECT 2064.120 2173.290 2064.380 2173.610 ;
        RECT 2064.120 2138.610 2064.380 2138.930 ;
        RECT 2064.180 2125.410 2064.320 2138.610 ;
        RECT 2064.180 2125.270 2064.780 2125.410 ;
        RECT 2064.640 2124.310 2064.780 2125.270 ;
        RECT 1559.040 2123.990 1559.300 2124.310 ;
        RECT 2064.580 2123.990 2064.840 2124.310 ;
        RECT 1559.100 2112.185 1559.240 2123.990 ;
        RECT 1559.100 2111.740 1559.450 2112.185 ;
        RECT 1559.170 2108.185 1559.450 2111.740 ;
      LAYER via2 ;
        RECT 2064.110 2608.000 2064.390 2608.280 ;
        RECT 2065.030 2608.000 2065.310 2608.280 ;
        RECT 2063.190 2511.440 2063.470 2511.720 ;
        RECT 2064.570 2511.440 2064.850 2511.720 ;
        RECT 2063.190 2463.160 2063.470 2463.440 ;
        RECT 2064.110 2463.160 2064.390 2463.440 ;
        RECT 2063.190 2270.040 2063.470 2270.320 ;
        RECT 2064.570 2270.040 2064.850 2270.320 ;
      LAYER met3 ;
        RECT 2064.085 2608.290 2064.415 2608.305 ;
        RECT 2065.005 2608.290 2065.335 2608.305 ;
        RECT 2064.085 2607.990 2065.335 2608.290 ;
        RECT 2064.085 2607.975 2064.415 2607.990 ;
        RECT 2065.005 2607.975 2065.335 2607.990 ;
        RECT 2063.165 2511.730 2063.495 2511.745 ;
        RECT 2064.545 2511.730 2064.875 2511.745 ;
        RECT 2063.165 2511.430 2064.875 2511.730 ;
        RECT 2063.165 2511.415 2063.495 2511.430 ;
        RECT 2064.545 2511.415 2064.875 2511.430 ;
        RECT 2063.165 2463.450 2063.495 2463.465 ;
        RECT 2064.085 2463.450 2064.415 2463.465 ;
        RECT 2063.165 2463.150 2064.415 2463.450 ;
        RECT 2063.165 2463.135 2063.495 2463.150 ;
        RECT 2064.085 2463.135 2064.415 2463.150 ;
        RECT 2063.165 2270.330 2063.495 2270.345 ;
        RECT 2064.545 2270.330 2064.875 2270.345 ;
        RECT 2063.165 2270.030 2064.875 2270.330 ;
        RECT 2063.165 2270.015 2063.495 2270.030 ;
        RECT 2064.545 2270.015 2064.875 2270.030 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1738.945 2898.245 1739.115 2946.355 ;
        RECT 1739.405 2815.285 1739.575 2849.455 ;
      LAYER mcon ;
        RECT 1738.945 2946.185 1739.115 2946.355 ;
        RECT 1739.405 2849.285 1739.575 2849.455 ;
      LAYER met1 ;
        RECT 1738.870 3464.160 1739.190 3464.220 ;
        RECT 1744.390 3464.160 1744.710 3464.220 ;
        RECT 1738.870 3464.020 1744.710 3464.160 ;
        RECT 1738.870 3463.960 1739.190 3464.020 ;
        RECT 1744.390 3463.960 1744.710 3464.020 ;
        RECT 1738.870 3367.600 1739.190 3367.660 ;
        RECT 1739.790 3367.600 1740.110 3367.660 ;
        RECT 1738.870 3367.460 1740.110 3367.600 ;
        RECT 1738.870 3367.400 1739.190 3367.460 ;
        RECT 1739.790 3367.400 1740.110 3367.460 ;
        RECT 1738.870 3270.700 1739.190 3270.760 ;
        RECT 1739.790 3270.700 1740.110 3270.760 ;
        RECT 1738.870 3270.560 1740.110 3270.700 ;
        RECT 1738.870 3270.500 1739.190 3270.560 ;
        RECT 1739.790 3270.500 1740.110 3270.560 ;
        RECT 1738.870 3174.140 1739.190 3174.200 ;
        RECT 1739.790 3174.140 1740.110 3174.200 ;
        RECT 1738.870 3174.000 1740.110 3174.140 ;
        RECT 1738.870 3173.940 1739.190 3174.000 ;
        RECT 1739.790 3173.940 1740.110 3174.000 ;
        RECT 1738.870 3077.580 1739.190 3077.640 ;
        RECT 1739.790 3077.580 1740.110 3077.640 ;
        RECT 1738.870 3077.440 1740.110 3077.580 ;
        RECT 1738.870 3077.380 1739.190 3077.440 ;
        RECT 1739.790 3077.380 1740.110 3077.440 ;
        RECT 1738.870 2981.020 1739.190 2981.080 ;
        RECT 1739.790 2981.020 1740.110 2981.080 ;
        RECT 1738.870 2980.880 1740.110 2981.020 ;
        RECT 1738.870 2980.820 1739.190 2980.880 ;
        RECT 1739.790 2980.820 1740.110 2980.880 ;
        RECT 1738.885 2946.340 1739.175 2946.385 ;
        RECT 1739.330 2946.340 1739.650 2946.400 ;
        RECT 1738.885 2946.200 1739.650 2946.340 ;
        RECT 1738.885 2946.155 1739.175 2946.200 ;
        RECT 1739.330 2946.140 1739.650 2946.200 ;
        RECT 1738.870 2898.400 1739.190 2898.460 ;
        RECT 1738.870 2898.260 1739.385 2898.400 ;
        RECT 1738.870 2898.200 1739.190 2898.260 ;
        RECT 1739.330 2849.440 1739.650 2849.500 ;
        RECT 1739.135 2849.300 1739.650 2849.440 ;
        RECT 1739.330 2849.240 1739.650 2849.300 ;
        RECT 1739.345 2815.440 1739.635 2815.485 ;
        RECT 1740.250 2815.440 1740.570 2815.500 ;
        RECT 1739.345 2815.300 1740.570 2815.440 ;
        RECT 1739.345 2815.255 1739.635 2815.300 ;
        RECT 1740.250 2815.240 1740.570 2815.300 ;
        RECT 1739.330 2753.220 1739.650 2753.280 ;
        RECT 1740.710 2753.220 1741.030 2753.280 ;
        RECT 1739.330 2753.080 1741.030 2753.220 ;
        RECT 1739.330 2753.020 1739.650 2753.080 ;
        RECT 1740.710 2753.020 1741.030 2753.080 ;
        RECT 1740.710 2719.220 1741.030 2719.280 ;
        RECT 1740.340 2719.080 1741.030 2719.220 ;
        RECT 1740.340 2718.600 1740.480 2719.080 ;
        RECT 1740.710 2719.020 1741.030 2719.080 ;
        RECT 1740.250 2718.340 1740.570 2718.600 ;
        RECT 1739.330 2656.660 1739.650 2656.720 ;
        RECT 1740.710 2656.660 1741.030 2656.720 ;
        RECT 1739.330 2656.520 1741.030 2656.660 ;
        RECT 1739.330 2656.460 1739.650 2656.520 ;
        RECT 1740.710 2656.460 1741.030 2656.520 ;
        RECT 1740.710 2622.660 1741.030 2622.720 ;
        RECT 1740.340 2622.520 1741.030 2622.660 ;
        RECT 1740.340 2622.040 1740.480 2622.520 ;
        RECT 1740.710 2622.460 1741.030 2622.520 ;
        RECT 1740.250 2621.780 1740.570 2622.040 ;
        RECT 1739.330 2560.100 1739.650 2560.160 ;
        RECT 1740.710 2560.100 1741.030 2560.160 ;
        RECT 1739.330 2559.960 1741.030 2560.100 ;
        RECT 1739.330 2559.900 1739.650 2559.960 ;
        RECT 1740.710 2559.900 1741.030 2559.960 ;
        RECT 1739.790 2511.820 1740.110 2511.880 ;
        RECT 1740.710 2511.820 1741.030 2511.880 ;
        RECT 1739.790 2511.680 1741.030 2511.820 ;
        RECT 1739.790 2511.620 1740.110 2511.680 ;
        RECT 1740.710 2511.620 1741.030 2511.680 ;
        RECT 1738.870 2401.320 1739.190 2401.380 ;
        RECT 1739.790 2401.320 1740.110 2401.380 ;
        RECT 1738.870 2401.180 1740.110 2401.320 ;
        RECT 1738.870 2401.120 1739.190 2401.180 ;
        RECT 1739.790 2401.120 1740.110 2401.180 ;
        RECT 1738.870 2304.760 1739.190 2304.820 ;
        RECT 1739.790 2304.760 1740.110 2304.820 ;
        RECT 1738.870 2304.620 1740.110 2304.760 ;
        RECT 1738.870 2304.560 1739.190 2304.620 ;
        RECT 1739.790 2304.560 1740.110 2304.620 ;
        RECT 1738.870 2208.200 1739.190 2208.260 ;
        RECT 1739.790 2208.200 1740.110 2208.260 ;
        RECT 1738.870 2208.060 1740.110 2208.200 ;
        RECT 1738.870 2208.000 1739.190 2208.060 ;
        RECT 1739.790 2208.000 1740.110 2208.060 ;
        RECT 1382.370 2122.180 1382.690 2122.240 ;
        RECT 1739.790 2122.180 1740.110 2122.240 ;
        RECT 1382.370 2122.040 1740.110 2122.180 ;
        RECT 1382.370 2121.980 1382.690 2122.040 ;
        RECT 1739.790 2121.980 1740.110 2122.040 ;
      LAYER via ;
        RECT 1738.900 3463.960 1739.160 3464.220 ;
        RECT 1744.420 3463.960 1744.680 3464.220 ;
        RECT 1738.900 3367.400 1739.160 3367.660 ;
        RECT 1739.820 3367.400 1740.080 3367.660 ;
        RECT 1738.900 3270.500 1739.160 3270.760 ;
        RECT 1739.820 3270.500 1740.080 3270.760 ;
        RECT 1738.900 3173.940 1739.160 3174.200 ;
        RECT 1739.820 3173.940 1740.080 3174.200 ;
        RECT 1738.900 3077.380 1739.160 3077.640 ;
        RECT 1739.820 3077.380 1740.080 3077.640 ;
        RECT 1738.900 2980.820 1739.160 2981.080 ;
        RECT 1739.820 2980.820 1740.080 2981.080 ;
        RECT 1739.360 2946.140 1739.620 2946.400 ;
        RECT 1738.900 2898.200 1739.160 2898.460 ;
        RECT 1739.360 2849.240 1739.620 2849.500 ;
        RECT 1740.280 2815.240 1740.540 2815.500 ;
        RECT 1739.360 2753.020 1739.620 2753.280 ;
        RECT 1740.740 2753.020 1741.000 2753.280 ;
        RECT 1740.740 2719.020 1741.000 2719.280 ;
        RECT 1740.280 2718.340 1740.540 2718.600 ;
        RECT 1739.360 2656.460 1739.620 2656.720 ;
        RECT 1740.740 2656.460 1741.000 2656.720 ;
        RECT 1740.740 2622.460 1741.000 2622.720 ;
        RECT 1740.280 2621.780 1740.540 2622.040 ;
        RECT 1739.360 2559.900 1739.620 2560.160 ;
        RECT 1740.740 2559.900 1741.000 2560.160 ;
        RECT 1739.820 2511.620 1740.080 2511.880 ;
        RECT 1740.740 2511.620 1741.000 2511.880 ;
        RECT 1738.900 2401.120 1739.160 2401.380 ;
        RECT 1739.820 2401.120 1740.080 2401.380 ;
        RECT 1738.900 2304.560 1739.160 2304.820 ;
        RECT 1739.820 2304.560 1740.080 2304.820 ;
        RECT 1738.900 2208.000 1739.160 2208.260 ;
        RECT 1739.820 2208.000 1740.080 2208.260 ;
        RECT 1382.400 2121.980 1382.660 2122.240 ;
        RECT 1739.820 2121.980 1740.080 2122.240 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3517.370 1744.160 3517.600 ;
        RECT 1744.020 3517.230 1744.620 3517.370 ;
        RECT 1744.480 3464.250 1744.620 3517.230 ;
        RECT 1738.900 3463.930 1739.160 3464.250 ;
        RECT 1744.420 3463.930 1744.680 3464.250 ;
        RECT 1738.960 3415.370 1739.100 3463.930 ;
        RECT 1738.960 3415.230 1740.020 3415.370 ;
        RECT 1739.880 3367.690 1740.020 3415.230 ;
        RECT 1738.900 3367.370 1739.160 3367.690 ;
        RECT 1739.820 3367.370 1740.080 3367.690 ;
        RECT 1738.960 3318.810 1739.100 3367.370 ;
        RECT 1738.960 3318.670 1740.020 3318.810 ;
        RECT 1739.880 3270.790 1740.020 3318.670 ;
        RECT 1738.900 3270.470 1739.160 3270.790 ;
        RECT 1739.820 3270.470 1740.080 3270.790 ;
        RECT 1738.960 3222.250 1739.100 3270.470 ;
        RECT 1738.960 3222.110 1740.020 3222.250 ;
        RECT 1739.880 3174.230 1740.020 3222.110 ;
        RECT 1738.900 3173.910 1739.160 3174.230 ;
        RECT 1739.820 3173.910 1740.080 3174.230 ;
        RECT 1738.960 3125.690 1739.100 3173.910 ;
        RECT 1738.960 3125.550 1740.020 3125.690 ;
        RECT 1739.880 3077.670 1740.020 3125.550 ;
        RECT 1738.900 3077.350 1739.160 3077.670 ;
        RECT 1739.820 3077.350 1740.080 3077.670 ;
        RECT 1738.960 3029.130 1739.100 3077.350 ;
        RECT 1738.960 3028.990 1740.020 3029.130 ;
        RECT 1739.880 2981.110 1740.020 3028.990 ;
        RECT 1738.900 2980.850 1739.160 2981.110 ;
        RECT 1738.900 2980.790 1739.560 2980.850 ;
        RECT 1739.820 2980.790 1740.080 2981.110 ;
        RECT 1738.960 2980.710 1739.560 2980.790 ;
        RECT 1739.420 2980.170 1739.560 2980.710 ;
        RECT 1739.420 2980.030 1740.020 2980.170 ;
        RECT 1739.880 2959.770 1740.020 2980.030 ;
        RECT 1739.420 2959.630 1740.020 2959.770 ;
        RECT 1739.420 2946.430 1739.560 2959.630 ;
        RECT 1739.360 2946.110 1739.620 2946.430 ;
        RECT 1738.900 2898.170 1739.160 2898.490 ;
        RECT 1738.960 2863.210 1739.100 2898.170 ;
        RECT 1738.960 2863.070 1739.560 2863.210 ;
        RECT 1739.420 2849.530 1739.560 2863.070 ;
        RECT 1739.360 2849.210 1739.620 2849.530 ;
        RECT 1740.280 2815.210 1740.540 2815.530 ;
        RECT 1740.340 2801.445 1740.480 2815.210 ;
        RECT 1739.350 2801.075 1739.630 2801.445 ;
        RECT 1740.270 2801.075 1740.550 2801.445 ;
        RECT 1739.420 2753.310 1739.560 2801.075 ;
        RECT 1739.360 2752.990 1739.620 2753.310 ;
        RECT 1740.740 2752.990 1741.000 2753.310 ;
        RECT 1740.800 2719.310 1740.940 2752.990 ;
        RECT 1740.740 2718.990 1741.000 2719.310 ;
        RECT 1740.280 2718.310 1740.540 2718.630 ;
        RECT 1740.340 2704.885 1740.480 2718.310 ;
        RECT 1739.350 2704.515 1739.630 2704.885 ;
        RECT 1740.270 2704.515 1740.550 2704.885 ;
        RECT 1739.420 2656.750 1739.560 2704.515 ;
        RECT 1739.360 2656.430 1739.620 2656.750 ;
        RECT 1740.740 2656.430 1741.000 2656.750 ;
        RECT 1740.800 2622.750 1740.940 2656.430 ;
        RECT 1740.740 2622.430 1741.000 2622.750 ;
        RECT 1740.280 2621.750 1740.540 2622.070 ;
        RECT 1740.340 2608.325 1740.480 2621.750 ;
        RECT 1739.350 2607.955 1739.630 2608.325 ;
        RECT 1740.270 2607.955 1740.550 2608.325 ;
        RECT 1739.420 2560.190 1739.560 2607.955 ;
        RECT 1739.360 2559.870 1739.620 2560.190 ;
        RECT 1740.740 2559.870 1741.000 2560.190 ;
        RECT 1740.800 2511.910 1740.940 2559.870 ;
        RECT 1739.820 2511.765 1740.080 2511.910 ;
        RECT 1739.810 2511.395 1740.090 2511.765 ;
        RECT 1740.740 2511.590 1741.000 2511.910 ;
        RECT 1739.350 2463.115 1739.630 2463.485 ;
        RECT 1739.420 2449.770 1739.560 2463.115 ;
        RECT 1739.420 2449.630 1740.020 2449.770 ;
        RECT 1739.880 2401.410 1740.020 2449.630 ;
        RECT 1738.900 2401.090 1739.160 2401.410 ;
        RECT 1739.820 2401.090 1740.080 2401.410 ;
        RECT 1738.960 2400.810 1739.100 2401.090 ;
        RECT 1738.960 2400.670 1739.560 2400.810 ;
        RECT 1739.420 2353.210 1739.560 2400.670 ;
        RECT 1739.420 2353.070 1740.020 2353.210 ;
        RECT 1739.880 2304.850 1740.020 2353.070 ;
        RECT 1738.900 2304.530 1739.160 2304.850 ;
        RECT 1739.820 2304.530 1740.080 2304.850 ;
        RECT 1738.960 2304.250 1739.100 2304.530 ;
        RECT 1738.960 2304.110 1739.560 2304.250 ;
        RECT 1739.420 2256.650 1739.560 2304.110 ;
        RECT 1739.420 2256.510 1740.020 2256.650 ;
        RECT 1739.880 2208.290 1740.020 2256.510 ;
        RECT 1738.900 2207.970 1739.160 2208.290 ;
        RECT 1739.820 2207.970 1740.080 2208.290 ;
        RECT 1738.960 2207.690 1739.100 2207.970 ;
        RECT 1738.960 2207.550 1739.560 2207.690 ;
        RECT 1739.420 2160.090 1739.560 2207.550 ;
        RECT 1739.420 2159.950 1740.020 2160.090 ;
        RECT 1739.880 2122.270 1740.020 2159.950 ;
        RECT 1382.400 2121.950 1382.660 2122.270 ;
        RECT 1739.820 2121.950 1740.080 2122.270 ;
        RECT 1382.460 2112.185 1382.600 2121.950 ;
        RECT 1382.460 2111.740 1382.810 2112.185 ;
        RECT 1382.530 2108.185 1382.810 2111.740 ;
      LAYER via2 ;
        RECT 1739.350 2801.120 1739.630 2801.400 ;
        RECT 1740.270 2801.120 1740.550 2801.400 ;
        RECT 1739.350 2704.560 1739.630 2704.840 ;
        RECT 1740.270 2704.560 1740.550 2704.840 ;
        RECT 1739.350 2608.000 1739.630 2608.280 ;
        RECT 1740.270 2608.000 1740.550 2608.280 ;
        RECT 1739.810 2511.440 1740.090 2511.720 ;
        RECT 1739.350 2463.160 1739.630 2463.440 ;
      LAYER met3 ;
        RECT 1739.325 2801.410 1739.655 2801.425 ;
        RECT 1740.245 2801.410 1740.575 2801.425 ;
        RECT 1739.325 2801.110 1740.575 2801.410 ;
        RECT 1739.325 2801.095 1739.655 2801.110 ;
        RECT 1740.245 2801.095 1740.575 2801.110 ;
        RECT 1739.325 2704.850 1739.655 2704.865 ;
        RECT 1740.245 2704.850 1740.575 2704.865 ;
        RECT 1739.325 2704.550 1740.575 2704.850 ;
        RECT 1739.325 2704.535 1739.655 2704.550 ;
        RECT 1740.245 2704.535 1740.575 2704.550 ;
        RECT 1739.325 2608.290 1739.655 2608.305 ;
        RECT 1740.245 2608.290 1740.575 2608.305 ;
        RECT 1739.325 2607.990 1740.575 2608.290 ;
        RECT 1739.325 2607.975 1739.655 2607.990 ;
        RECT 1740.245 2607.975 1740.575 2607.990 ;
        RECT 1739.070 2511.730 1739.450 2511.740 ;
        RECT 1739.785 2511.730 1740.115 2511.745 ;
        RECT 1739.070 2511.430 1740.115 2511.730 ;
        RECT 1739.070 2511.420 1739.450 2511.430 ;
        RECT 1739.785 2511.415 1740.115 2511.430 ;
        RECT 1739.325 2463.460 1739.655 2463.465 ;
        RECT 1739.070 2463.450 1739.655 2463.460 ;
        RECT 1739.070 2463.150 1739.880 2463.450 ;
        RECT 1739.070 2463.140 1739.655 2463.150 ;
        RECT 1739.325 2463.135 1739.655 2463.140 ;
      LAYER via3 ;
        RECT 1739.100 2511.420 1739.420 2511.740 ;
        RECT 1739.100 2463.140 1739.420 2463.460 ;
      LAYER met4 ;
        RECT 1739.095 2511.415 1739.425 2511.745 ;
        RECT 1739.110 2463.465 1739.410 2511.415 ;
        RECT 1739.095 2463.135 1739.425 2463.465 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1416.485 3332.765 1416.655 3415.555 ;
        RECT 1415.565 3008.405 1415.735 3042.915 ;
        RECT 1416.485 2946.525 1416.655 2994.635 ;
        RECT 1415.105 2753.065 1415.275 2801.175 ;
        RECT 1415.565 2428.705 1415.735 2463.215 ;
        RECT 1415.565 2331.805 1415.735 2366.655 ;
        RECT 1415.565 2138.685 1415.735 2173.535 ;
      LAYER mcon ;
        RECT 1416.485 3415.385 1416.655 3415.555 ;
        RECT 1415.565 3042.745 1415.735 3042.915 ;
        RECT 1416.485 2994.465 1416.655 2994.635 ;
        RECT 1415.105 2801.005 1415.275 2801.175 ;
        RECT 1415.565 2463.045 1415.735 2463.215 ;
        RECT 1415.565 2366.485 1415.735 2366.655 ;
        RECT 1415.565 2173.365 1415.735 2173.535 ;
      LAYER met1 ;
        RECT 1416.410 3491.360 1416.730 3491.420 ;
        RECT 1419.630 3491.360 1419.950 3491.420 ;
        RECT 1416.410 3491.220 1419.950 3491.360 ;
        RECT 1416.410 3491.160 1416.730 3491.220 ;
        RECT 1419.630 3491.160 1419.950 3491.220 ;
        RECT 1415.490 3470.620 1415.810 3470.680 ;
        RECT 1416.410 3470.620 1416.730 3470.680 ;
        RECT 1415.490 3470.480 1416.730 3470.620 ;
        RECT 1415.490 3470.420 1415.810 3470.480 ;
        RECT 1416.410 3470.420 1416.730 3470.480 ;
        RECT 1415.490 3463.820 1415.810 3463.880 ;
        RECT 1416.410 3463.820 1416.730 3463.880 ;
        RECT 1415.490 3463.680 1416.730 3463.820 ;
        RECT 1415.490 3463.620 1415.810 3463.680 ;
        RECT 1416.410 3463.620 1416.730 3463.680 ;
        RECT 1414.570 3415.540 1414.890 3415.600 ;
        RECT 1416.425 3415.540 1416.715 3415.585 ;
        RECT 1414.570 3415.400 1416.715 3415.540 ;
        RECT 1414.570 3415.340 1414.890 3415.400 ;
        RECT 1416.425 3415.355 1416.715 3415.400 ;
        RECT 1416.425 3332.920 1416.715 3332.965 ;
        RECT 1416.870 3332.920 1417.190 3332.980 ;
        RECT 1416.425 3332.780 1417.190 3332.920 ;
        RECT 1416.425 3332.735 1416.715 3332.780 ;
        RECT 1416.870 3332.720 1417.190 3332.780 ;
        RECT 1415.490 3236.360 1415.810 3236.420 ;
        RECT 1415.950 3236.360 1416.270 3236.420 ;
        RECT 1415.490 3236.220 1416.270 3236.360 ;
        RECT 1415.490 3236.160 1415.810 3236.220 ;
        RECT 1415.950 3236.160 1416.270 3236.220 ;
        RECT 1415.490 3202.020 1415.810 3202.080 ;
        RECT 1415.950 3202.020 1416.270 3202.080 ;
        RECT 1415.490 3201.880 1416.270 3202.020 ;
        RECT 1415.490 3201.820 1415.810 3201.880 ;
        RECT 1415.950 3201.820 1416.270 3201.880 ;
        RECT 1415.030 3153.400 1415.350 3153.460 ;
        RECT 1415.950 3153.400 1416.270 3153.460 ;
        RECT 1415.030 3153.260 1416.270 3153.400 ;
        RECT 1415.030 3153.200 1415.350 3153.260 ;
        RECT 1415.950 3153.200 1416.270 3153.260 ;
        RECT 1415.030 3056.840 1415.350 3056.900 ;
        RECT 1415.950 3056.840 1416.270 3056.900 ;
        RECT 1415.030 3056.700 1416.270 3056.840 ;
        RECT 1415.030 3056.640 1415.350 3056.700 ;
        RECT 1415.950 3056.640 1416.270 3056.700 ;
        RECT 1415.490 3042.900 1415.810 3042.960 ;
        RECT 1415.295 3042.760 1415.810 3042.900 ;
        RECT 1415.490 3042.700 1415.810 3042.760 ;
        RECT 1415.505 3008.560 1415.795 3008.605 ;
        RECT 1416.410 3008.560 1416.730 3008.620 ;
        RECT 1415.505 3008.420 1416.730 3008.560 ;
        RECT 1415.505 3008.375 1415.795 3008.420 ;
        RECT 1416.410 3008.360 1416.730 3008.420 ;
        RECT 1416.410 2994.620 1416.730 2994.680 ;
        RECT 1416.215 2994.480 1416.730 2994.620 ;
        RECT 1416.410 2994.420 1416.730 2994.480 ;
        RECT 1416.425 2946.680 1416.715 2946.725 ;
        RECT 1416.870 2946.680 1417.190 2946.740 ;
        RECT 1416.425 2946.540 1417.190 2946.680 ;
        RECT 1416.425 2946.495 1416.715 2946.540 ;
        RECT 1416.870 2946.480 1417.190 2946.540 ;
        RECT 1416.870 2912.340 1417.190 2912.400 ;
        RECT 1416.500 2912.200 1417.190 2912.340 ;
        RECT 1416.500 2911.720 1416.640 2912.200 ;
        RECT 1416.870 2912.140 1417.190 2912.200 ;
        RECT 1416.410 2911.460 1416.730 2911.720 ;
        RECT 1415.030 2815.580 1415.350 2815.840 ;
        RECT 1415.120 2815.160 1415.260 2815.580 ;
        RECT 1415.030 2814.900 1415.350 2815.160 ;
        RECT 1415.030 2801.160 1415.350 2801.220 ;
        RECT 1414.835 2801.020 1415.350 2801.160 ;
        RECT 1415.030 2800.960 1415.350 2801.020 ;
        RECT 1415.045 2753.220 1415.335 2753.265 ;
        RECT 1415.950 2753.220 1416.270 2753.280 ;
        RECT 1415.045 2753.080 1416.270 2753.220 ;
        RECT 1415.045 2753.035 1415.335 2753.080 ;
        RECT 1415.950 2753.020 1416.270 2753.080 ;
        RECT 1415.030 2718.200 1415.350 2718.260 ;
        RECT 1415.950 2718.200 1416.270 2718.260 ;
        RECT 1415.030 2718.060 1416.270 2718.200 ;
        RECT 1415.030 2718.000 1415.350 2718.060 ;
        RECT 1415.950 2718.000 1416.270 2718.060 ;
        RECT 1415.030 2670.260 1415.350 2670.320 ;
        RECT 1415.950 2670.260 1416.270 2670.320 ;
        RECT 1415.030 2670.120 1416.270 2670.260 ;
        RECT 1415.030 2670.060 1415.350 2670.120 ;
        RECT 1415.950 2670.060 1416.270 2670.120 ;
        RECT 1415.950 2622.120 1416.270 2622.380 ;
        RECT 1416.040 2621.980 1416.180 2622.120 ;
        RECT 1416.410 2621.980 1416.730 2622.040 ;
        RECT 1416.040 2621.840 1416.730 2621.980 ;
        RECT 1416.410 2621.780 1416.730 2621.840 ;
        RECT 1415.490 2560.100 1415.810 2560.160 ;
        RECT 1416.870 2560.100 1417.190 2560.160 ;
        RECT 1415.490 2559.960 1417.190 2560.100 ;
        RECT 1415.490 2559.900 1415.810 2559.960 ;
        RECT 1416.870 2559.900 1417.190 2559.960 ;
        RECT 1415.950 2511.820 1416.270 2511.880 ;
        RECT 1416.870 2511.820 1417.190 2511.880 ;
        RECT 1415.950 2511.680 1417.190 2511.820 ;
        RECT 1415.950 2511.620 1416.270 2511.680 ;
        RECT 1416.870 2511.620 1417.190 2511.680 ;
        RECT 1415.490 2463.200 1415.810 2463.260 ;
        RECT 1415.295 2463.060 1415.810 2463.200 ;
        RECT 1415.490 2463.000 1415.810 2463.060 ;
        RECT 1415.490 2428.860 1415.810 2428.920 ;
        RECT 1415.295 2428.720 1415.810 2428.860 ;
        RECT 1415.490 2428.660 1415.810 2428.720 ;
        RECT 1415.030 2380.580 1415.350 2380.640 ;
        RECT 1415.950 2380.580 1416.270 2380.640 ;
        RECT 1415.030 2380.440 1416.270 2380.580 ;
        RECT 1415.030 2380.380 1415.350 2380.440 ;
        RECT 1415.950 2380.380 1416.270 2380.440 ;
        RECT 1415.490 2366.640 1415.810 2366.700 ;
        RECT 1415.295 2366.500 1415.810 2366.640 ;
        RECT 1415.490 2366.440 1415.810 2366.500 ;
        RECT 1415.490 2331.960 1415.810 2332.020 ;
        RECT 1415.295 2331.820 1415.810 2331.960 ;
        RECT 1415.490 2331.760 1415.810 2331.820 ;
        RECT 1414.570 2235.540 1414.890 2235.800 ;
        RECT 1414.660 2235.400 1414.800 2235.540 ;
        RECT 1415.030 2235.400 1415.350 2235.460 ;
        RECT 1414.660 2235.260 1415.350 2235.400 ;
        RECT 1415.030 2235.200 1415.350 2235.260 ;
        RECT 1415.490 2173.520 1415.810 2173.580 ;
        RECT 1415.295 2173.380 1415.810 2173.520 ;
        RECT 1415.490 2173.320 1415.810 2173.380 ;
        RECT 1415.490 2138.840 1415.810 2138.900 ;
        RECT 1415.295 2138.700 1415.810 2138.840 ;
        RECT 1415.490 2138.640 1415.810 2138.700 ;
        RECT 1205.270 2121.840 1205.590 2121.900 ;
        RECT 1415.950 2121.840 1416.270 2121.900 ;
        RECT 1205.270 2121.700 1416.270 2121.840 ;
        RECT 1205.270 2121.640 1205.590 2121.700 ;
        RECT 1415.950 2121.640 1416.270 2121.700 ;
      LAYER via ;
        RECT 1416.440 3491.160 1416.700 3491.420 ;
        RECT 1419.660 3491.160 1419.920 3491.420 ;
        RECT 1415.520 3470.420 1415.780 3470.680 ;
        RECT 1416.440 3470.420 1416.700 3470.680 ;
        RECT 1415.520 3463.620 1415.780 3463.880 ;
        RECT 1416.440 3463.620 1416.700 3463.880 ;
        RECT 1414.600 3415.340 1414.860 3415.600 ;
        RECT 1416.900 3332.720 1417.160 3332.980 ;
        RECT 1415.520 3236.160 1415.780 3236.420 ;
        RECT 1415.980 3236.160 1416.240 3236.420 ;
        RECT 1415.520 3201.820 1415.780 3202.080 ;
        RECT 1415.980 3201.820 1416.240 3202.080 ;
        RECT 1415.060 3153.200 1415.320 3153.460 ;
        RECT 1415.980 3153.200 1416.240 3153.460 ;
        RECT 1415.060 3056.640 1415.320 3056.900 ;
        RECT 1415.980 3056.640 1416.240 3056.900 ;
        RECT 1415.520 3042.700 1415.780 3042.960 ;
        RECT 1416.440 3008.360 1416.700 3008.620 ;
        RECT 1416.440 2994.420 1416.700 2994.680 ;
        RECT 1416.900 2946.480 1417.160 2946.740 ;
        RECT 1416.900 2912.140 1417.160 2912.400 ;
        RECT 1416.440 2911.460 1416.700 2911.720 ;
        RECT 1415.060 2815.580 1415.320 2815.840 ;
        RECT 1415.060 2814.900 1415.320 2815.160 ;
        RECT 1415.060 2800.960 1415.320 2801.220 ;
        RECT 1415.980 2753.020 1416.240 2753.280 ;
        RECT 1415.060 2718.000 1415.320 2718.260 ;
        RECT 1415.980 2718.000 1416.240 2718.260 ;
        RECT 1415.060 2670.060 1415.320 2670.320 ;
        RECT 1415.980 2670.060 1416.240 2670.320 ;
        RECT 1415.980 2622.120 1416.240 2622.380 ;
        RECT 1416.440 2621.780 1416.700 2622.040 ;
        RECT 1415.520 2559.900 1415.780 2560.160 ;
        RECT 1416.900 2559.900 1417.160 2560.160 ;
        RECT 1415.980 2511.620 1416.240 2511.880 ;
        RECT 1416.900 2511.620 1417.160 2511.880 ;
        RECT 1415.520 2463.000 1415.780 2463.260 ;
        RECT 1415.520 2428.660 1415.780 2428.920 ;
        RECT 1415.060 2380.380 1415.320 2380.640 ;
        RECT 1415.980 2380.380 1416.240 2380.640 ;
        RECT 1415.520 2366.440 1415.780 2366.700 ;
        RECT 1415.520 2331.760 1415.780 2332.020 ;
        RECT 1414.600 2235.540 1414.860 2235.800 ;
        RECT 1415.060 2235.200 1415.320 2235.460 ;
        RECT 1415.520 2173.320 1415.780 2173.580 ;
        RECT 1415.520 2138.640 1415.780 2138.900 ;
        RECT 1205.300 2121.640 1205.560 2121.900 ;
        RECT 1415.980 2121.640 1416.240 2121.900 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3517.370 1419.400 3517.600 ;
        RECT 1419.260 3517.230 1419.860 3517.370 ;
        RECT 1419.720 3491.450 1419.860 3517.230 ;
        RECT 1416.440 3491.130 1416.700 3491.450 ;
        RECT 1419.660 3491.130 1419.920 3491.450 ;
        RECT 1416.500 3470.710 1416.640 3491.130 ;
        RECT 1415.520 3470.390 1415.780 3470.710 ;
        RECT 1416.440 3470.390 1416.700 3470.710 ;
        RECT 1415.580 3463.910 1415.720 3470.390 ;
        RECT 1415.520 3463.590 1415.780 3463.910 ;
        RECT 1416.440 3463.590 1416.700 3463.910 ;
        RECT 1416.500 3416.165 1416.640 3463.590 ;
        RECT 1414.590 3415.795 1414.870 3416.165 ;
        RECT 1416.430 3415.795 1416.710 3416.165 ;
        RECT 1414.660 3415.630 1414.800 3415.795 ;
        RECT 1414.600 3415.310 1414.860 3415.630 ;
        RECT 1416.900 3332.690 1417.160 3333.010 ;
        RECT 1416.960 3298.410 1417.100 3332.690 ;
        RECT 1416.040 3298.270 1417.100 3298.410 ;
        RECT 1416.040 3236.450 1416.180 3298.270 ;
        RECT 1415.520 3236.130 1415.780 3236.450 ;
        RECT 1415.980 3236.130 1416.240 3236.450 ;
        RECT 1415.580 3202.110 1415.720 3236.130 ;
        RECT 1415.520 3201.790 1415.780 3202.110 ;
        RECT 1415.980 3201.790 1416.240 3202.110 ;
        RECT 1416.040 3153.490 1416.180 3201.790 ;
        RECT 1415.060 3153.170 1415.320 3153.490 ;
        RECT 1415.980 3153.170 1416.240 3153.490 ;
        RECT 1415.120 3152.890 1415.260 3153.170 ;
        RECT 1415.120 3152.750 1415.720 3152.890 ;
        RECT 1415.580 3105.290 1415.720 3152.750 ;
        RECT 1415.580 3105.150 1416.180 3105.290 ;
        RECT 1416.040 3056.930 1416.180 3105.150 ;
        RECT 1415.060 3056.610 1415.320 3056.930 ;
        RECT 1415.980 3056.610 1416.240 3056.930 ;
        RECT 1415.120 3056.330 1415.260 3056.610 ;
        RECT 1415.120 3056.190 1415.720 3056.330 ;
        RECT 1415.580 3042.990 1415.720 3056.190 ;
        RECT 1415.520 3042.670 1415.780 3042.990 ;
        RECT 1416.440 3008.330 1416.700 3008.650 ;
        RECT 1416.500 2994.710 1416.640 3008.330 ;
        RECT 1416.440 2994.390 1416.700 2994.710 ;
        RECT 1416.900 2946.450 1417.160 2946.770 ;
        RECT 1416.960 2912.430 1417.100 2946.450 ;
        RECT 1416.900 2912.110 1417.160 2912.430 ;
        RECT 1416.440 2911.430 1416.700 2911.750 ;
        RECT 1416.500 2863.210 1416.640 2911.430 ;
        RECT 1415.580 2863.070 1416.640 2863.210 ;
        RECT 1415.580 2849.610 1415.720 2863.070 ;
        RECT 1415.120 2849.470 1415.720 2849.610 ;
        RECT 1415.120 2815.870 1415.260 2849.470 ;
        RECT 1415.060 2815.550 1415.320 2815.870 ;
        RECT 1415.060 2814.870 1415.320 2815.190 ;
        RECT 1415.120 2801.250 1415.260 2814.870 ;
        RECT 1415.060 2800.930 1415.320 2801.250 ;
        RECT 1415.980 2752.990 1416.240 2753.310 ;
        RECT 1416.040 2718.290 1416.180 2752.990 ;
        RECT 1415.060 2717.970 1415.320 2718.290 ;
        RECT 1415.980 2717.970 1416.240 2718.290 ;
        RECT 1415.120 2670.350 1415.260 2717.970 ;
        RECT 1415.060 2670.030 1415.320 2670.350 ;
        RECT 1415.980 2670.030 1416.240 2670.350 ;
        RECT 1416.040 2622.410 1416.180 2670.030 ;
        RECT 1415.980 2622.090 1416.240 2622.410 ;
        RECT 1416.440 2621.750 1416.700 2622.070 ;
        RECT 1416.500 2608.325 1416.640 2621.750 ;
        RECT 1415.510 2607.955 1415.790 2608.325 ;
        RECT 1416.430 2607.955 1416.710 2608.325 ;
        RECT 1415.580 2560.190 1415.720 2607.955 ;
        RECT 1415.520 2559.870 1415.780 2560.190 ;
        RECT 1416.900 2559.870 1417.160 2560.190 ;
        RECT 1416.960 2511.910 1417.100 2559.870 ;
        RECT 1415.980 2511.765 1416.240 2511.910 ;
        RECT 1414.590 2511.395 1414.870 2511.765 ;
        RECT 1415.970 2511.395 1416.250 2511.765 ;
        RECT 1416.900 2511.590 1417.160 2511.910 ;
        RECT 1414.660 2463.485 1414.800 2511.395 ;
        RECT 1414.590 2463.115 1414.870 2463.485 ;
        RECT 1415.510 2463.115 1415.790 2463.485 ;
        RECT 1415.520 2462.970 1415.780 2463.115 ;
        RECT 1415.520 2428.630 1415.780 2428.950 ;
        RECT 1415.580 2415.090 1415.720 2428.630 ;
        RECT 1415.580 2414.950 1416.180 2415.090 ;
        RECT 1416.040 2380.670 1416.180 2414.950 ;
        RECT 1415.060 2380.410 1415.320 2380.670 ;
        RECT 1415.060 2380.350 1415.720 2380.410 ;
        RECT 1415.980 2380.350 1416.240 2380.670 ;
        RECT 1415.120 2380.270 1415.720 2380.350 ;
        RECT 1415.580 2366.730 1415.720 2380.270 ;
        RECT 1415.520 2366.410 1415.780 2366.730 ;
        RECT 1415.520 2331.730 1415.780 2332.050 ;
        RECT 1415.580 2318.530 1415.720 2331.730 ;
        RECT 1415.580 2318.390 1416.180 2318.530 ;
        RECT 1416.040 2270.365 1416.180 2318.390 ;
        RECT 1414.590 2269.995 1414.870 2270.365 ;
        RECT 1415.970 2269.995 1416.250 2270.365 ;
        RECT 1414.660 2235.830 1414.800 2269.995 ;
        RECT 1414.600 2235.510 1414.860 2235.830 ;
        RECT 1415.060 2235.170 1415.320 2235.490 ;
        RECT 1415.120 2187.290 1415.260 2235.170 ;
        RECT 1415.120 2187.150 1415.720 2187.290 ;
        RECT 1415.580 2173.610 1415.720 2187.150 ;
        RECT 1415.520 2173.290 1415.780 2173.610 ;
        RECT 1415.520 2138.610 1415.780 2138.930 ;
        RECT 1415.580 2125.410 1415.720 2138.610 ;
        RECT 1415.580 2125.270 1416.180 2125.410 ;
        RECT 1416.040 2121.930 1416.180 2125.270 ;
        RECT 1205.300 2121.610 1205.560 2121.930 ;
        RECT 1415.980 2121.610 1416.240 2121.930 ;
        RECT 1205.360 2112.185 1205.500 2121.610 ;
        RECT 1205.360 2111.740 1205.710 2112.185 ;
        RECT 1205.430 2108.185 1205.710 2111.740 ;
      LAYER via2 ;
        RECT 1414.590 3415.840 1414.870 3416.120 ;
        RECT 1416.430 3415.840 1416.710 3416.120 ;
        RECT 1415.510 2608.000 1415.790 2608.280 ;
        RECT 1416.430 2608.000 1416.710 2608.280 ;
        RECT 1414.590 2511.440 1414.870 2511.720 ;
        RECT 1415.970 2511.440 1416.250 2511.720 ;
        RECT 1414.590 2463.160 1414.870 2463.440 ;
        RECT 1415.510 2463.160 1415.790 2463.440 ;
        RECT 1414.590 2270.040 1414.870 2270.320 ;
        RECT 1415.970 2270.040 1416.250 2270.320 ;
      LAYER met3 ;
        RECT 1414.565 3416.130 1414.895 3416.145 ;
        RECT 1416.405 3416.130 1416.735 3416.145 ;
        RECT 1414.565 3415.830 1416.735 3416.130 ;
        RECT 1414.565 3415.815 1414.895 3415.830 ;
        RECT 1416.405 3415.815 1416.735 3415.830 ;
        RECT 1415.485 2608.290 1415.815 2608.305 ;
        RECT 1416.405 2608.290 1416.735 2608.305 ;
        RECT 1415.485 2607.990 1416.735 2608.290 ;
        RECT 1415.485 2607.975 1415.815 2607.990 ;
        RECT 1416.405 2607.975 1416.735 2607.990 ;
        RECT 1414.565 2511.730 1414.895 2511.745 ;
        RECT 1415.945 2511.730 1416.275 2511.745 ;
        RECT 1414.565 2511.430 1416.275 2511.730 ;
        RECT 1414.565 2511.415 1414.895 2511.430 ;
        RECT 1415.945 2511.415 1416.275 2511.430 ;
        RECT 1414.565 2463.450 1414.895 2463.465 ;
        RECT 1415.485 2463.450 1415.815 2463.465 ;
        RECT 1414.565 2463.150 1415.815 2463.450 ;
        RECT 1414.565 2463.135 1414.895 2463.150 ;
        RECT 1415.485 2463.135 1415.815 2463.150 ;
        RECT 1414.565 2270.330 1414.895 2270.345 ;
        RECT 1415.945 2270.330 1416.275 2270.345 ;
        RECT 1414.565 2270.030 1416.275 2270.330 ;
        RECT 1414.565 2270.015 1414.895 2270.030 ;
        RECT 1415.945 2270.015 1416.275 2270.030 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2012.110 386.140 2012.430 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2012.110 386.000 2901.150 386.140 ;
        RECT 2012.110 385.940 2012.430 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2012.140 385.940 2012.400 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2012.130 669.955 2012.410 670.325 ;
        RECT 2012.200 386.230 2012.340 669.955 ;
        RECT 2012.140 385.910 2012.400 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2012.130 670.000 2012.410 670.280 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 1997.465 670.290 2001.465 670.440 ;
        RECT 2012.105 670.290 2012.435 670.305 ;
        RECT 1997.465 669.990 2012.435 670.290 ;
        RECT 1997.465 669.840 2001.465 669.990 ;
        RECT 2012.105 669.975 2012.435 669.990 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1090.345 2898.245 1090.515 2946.355 ;
        RECT 1090.805 2815.285 1090.975 2849.455 ;
      LAYER mcon ;
        RECT 1090.345 2946.185 1090.515 2946.355 ;
        RECT 1090.805 2849.285 1090.975 2849.455 ;
      LAYER met1 ;
        RECT 1090.270 3464.160 1090.590 3464.220 ;
        RECT 1095.330 3464.160 1095.650 3464.220 ;
        RECT 1090.270 3464.020 1095.650 3464.160 ;
        RECT 1090.270 3463.960 1090.590 3464.020 ;
        RECT 1095.330 3463.960 1095.650 3464.020 ;
        RECT 1090.270 3367.600 1090.590 3367.660 ;
        RECT 1091.190 3367.600 1091.510 3367.660 ;
        RECT 1090.270 3367.460 1091.510 3367.600 ;
        RECT 1090.270 3367.400 1090.590 3367.460 ;
        RECT 1091.190 3367.400 1091.510 3367.460 ;
        RECT 1090.270 3270.700 1090.590 3270.760 ;
        RECT 1091.190 3270.700 1091.510 3270.760 ;
        RECT 1090.270 3270.560 1091.510 3270.700 ;
        RECT 1090.270 3270.500 1090.590 3270.560 ;
        RECT 1091.190 3270.500 1091.510 3270.560 ;
        RECT 1090.270 3174.140 1090.590 3174.200 ;
        RECT 1091.190 3174.140 1091.510 3174.200 ;
        RECT 1090.270 3174.000 1091.510 3174.140 ;
        RECT 1090.270 3173.940 1090.590 3174.000 ;
        RECT 1091.190 3173.940 1091.510 3174.000 ;
        RECT 1090.270 3077.580 1090.590 3077.640 ;
        RECT 1091.190 3077.580 1091.510 3077.640 ;
        RECT 1090.270 3077.440 1091.510 3077.580 ;
        RECT 1090.270 3077.380 1090.590 3077.440 ;
        RECT 1091.190 3077.380 1091.510 3077.440 ;
        RECT 1090.270 2981.020 1090.590 2981.080 ;
        RECT 1091.190 2981.020 1091.510 2981.080 ;
        RECT 1090.270 2980.880 1091.510 2981.020 ;
        RECT 1090.270 2980.820 1090.590 2980.880 ;
        RECT 1091.190 2980.820 1091.510 2980.880 ;
        RECT 1090.285 2946.340 1090.575 2946.385 ;
        RECT 1090.730 2946.340 1091.050 2946.400 ;
        RECT 1090.285 2946.200 1091.050 2946.340 ;
        RECT 1090.285 2946.155 1090.575 2946.200 ;
        RECT 1090.730 2946.140 1091.050 2946.200 ;
        RECT 1090.270 2898.400 1090.590 2898.460 ;
        RECT 1090.075 2898.260 1090.590 2898.400 ;
        RECT 1090.270 2898.200 1090.590 2898.260 ;
        RECT 1090.730 2849.440 1091.050 2849.500 ;
        RECT 1090.535 2849.300 1091.050 2849.440 ;
        RECT 1090.730 2849.240 1091.050 2849.300 ;
        RECT 1090.745 2815.440 1091.035 2815.485 ;
        RECT 1091.650 2815.440 1091.970 2815.500 ;
        RECT 1090.745 2815.300 1091.970 2815.440 ;
        RECT 1090.745 2815.255 1091.035 2815.300 ;
        RECT 1091.650 2815.240 1091.970 2815.300 ;
        RECT 1090.730 2753.220 1091.050 2753.280 ;
        RECT 1092.110 2753.220 1092.430 2753.280 ;
        RECT 1090.730 2753.080 1092.430 2753.220 ;
        RECT 1090.730 2753.020 1091.050 2753.080 ;
        RECT 1092.110 2753.020 1092.430 2753.080 ;
        RECT 1092.110 2719.220 1092.430 2719.280 ;
        RECT 1091.740 2719.080 1092.430 2719.220 ;
        RECT 1091.740 2718.600 1091.880 2719.080 ;
        RECT 1092.110 2719.020 1092.430 2719.080 ;
        RECT 1091.650 2718.340 1091.970 2718.600 ;
        RECT 1090.730 2656.660 1091.050 2656.720 ;
        RECT 1092.110 2656.660 1092.430 2656.720 ;
        RECT 1090.730 2656.520 1092.430 2656.660 ;
        RECT 1090.730 2656.460 1091.050 2656.520 ;
        RECT 1092.110 2656.460 1092.430 2656.520 ;
        RECT 1092.110 2622.660 1092.430 2622.720 ;
        RECT 1091.740 2622.520 1092.430 2622.660 ;
        RECT 1091.740 2622.040 1091.880 2622.520 ;
        RECT 1092.110 2622.460 1092.430 2622.520 ;
        RECT 1091.650 2621.780 1091.970 2622.040 ;
        RECT 1090.730 2560.100 1091.050 2560.160 ;
        RECT 1092.110 2560.100 1092.430 2560.160 ;
        RECT 1090.730 2559.960 1092.430 2560.100 ;
        RECT 1090.730 2559.900 1091.050 2559.960 ;
        RECT 1092.110 2559.900 1092.430 2559.960 ;
        RECT 1091.190 2511.820 1091.510 2511.880 ;
        RECT 1092.110 2511.820 1092.430 2511.880 ;
        RECT 1091.190 2511.680 1092.430 2511.820 ;
        RECT 1091.190 2511.620 1091.510 2511.680 ;
        RECT 1092.110 2511.620 1092.430 2511.680 ;
        RECT 1090.270 2401.320 1090.590 2401.380 ;
        RECT 1091.190 2401.320 1091.510 2401.380 ;
        RECT 1090.270 2401.180 1091.510 2401.320 ;
        RECT 1090.270 2401.120 1090.590 2401.180 ;
        RECT 1091.190 2401.120 1091.510 2401.180 ;
        RECT 1090.270 2304.760 1090.590 2304.820 ;
        RECT 1091.190 2304.760 1091.510 2304.820 ;
        RECT 1090.270 2304.620 1091.510 2304.760 ;
        RECT 1090.270 2304.560 1090.590 2304.620 ;
        RECT 1091.190 2304.560 1091.510 2304.620 ;
        RECT 1090.270 2208.200 1090.590 2208.260 ;
        RECT 1091.190 2208.200 1091.510 2208.260 ;
        RECT 1090.270 2208.060 1091.510 2208.200 ;
        RECT 1090.270 2208.000 1090.590 2208.060 ;
        RECT 1091.190 2208.000 1091.510 2208.060 ;
        RECT 1028.630 2122.180 1028.950 2122.240 ;
        RECT 1091.190 2122.180 1091.510 2122.240 ;
        RECT 1028.630 2122.040 1091.510 2122.180 ;
        RECT 1028.630 2121.980 1028.950 2122.040 ;
        RECT 1091.190 2121.980 1091.510 2122.040 ;
      LAYER via ;
        RECT 1090.300 3463.960 1090.560 3464.220 ;
        RECT 1095.360 3463.960 1095.620 3464.220 ;
        RECT 1090.300 3367.400 1090.560 3367.660 ;
        RECT 1091.220 3367.400 1091.480 3367.660 ;
        RECT 1090.300 3270.500 1090.560 3270.760 ;
        RECT 1091.220 3270.500 1091.480 3270.760 ;
        RECT 1090.300 3173.940 1090.560 3174.200 ;
        RECT 1091.220 3173.940 1091.480 3174.200 ;
        RECT 1090.300 3077.380 1090.560 3077.640 ;
        RECT 1091.220 3077.380 1091.480 3077.640 ;
        RECT 1090.300 2980.820 1090.560 2981.080 ;
        RECT 1091.220 2980.820 1091.480 2981.080 ;
        RECT 1090.760 2946.140 1091.020 2946.400 ;
        RECT 1090.300 2898.200 1090.560 2898.460 ;
        RECT 1090.760 2849.240 1091.020 2849.500 ;
        RECT 1091.680 2815.240 1091.940 2815.500 ;
        RECT 1090.760 2753.020 1091.020 2753.280 ;
        RECT 1092.140 2753.020 1092.400 2753.280 ;
        RECT 1092.140 2719.020 1092.400 2719.280 ;
        RECT 1091.680 2718.340 1091.940 2718.600 ;
        RECT 1090.760 2656.460 1091.020 2656.720 ;
        RECT 1092.140 2656.460 1092.400 2656.720 ;
        RECT 1092.140 2622.460 1092.400 2622.720 ;
        RECT 1091.680 2621.780 1091.940 2622.040 ;
        RECT 1090.760 2559.900 1091.020 2560.160 ;
        RECT 1092.140 2559.900 1092.400 2560.160 ;
        RECT 1091.220 2511.620 1091.480 2511.880 ;
        RECT 1092.140 2511.620 1092.400 2511.880 ;
        RECT 1090.300 2401.120 1090.560 2401.380 ;
        RECT 1091.220 2401.120 1091.480 2401.380 ;
        RECT 1090.300 2304.560 1090.560 2304.820 ;
        RECT 1091.220 2304.560 1091.480 2304.820 ;
        RECT 1090.300 2208.000 1090.560 2208.260 ;
        RECT 1091.220 2208.000 1091.480 2208.260 ;
        RECT 1028.660 2121.980 1028.920 2122.240 ;
        RECT 1091.220 2121.980 1091.480 2122.240 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.960 3517.230 1095.560 3517.370 ;
        RECT 1095.420 3464.250 1095.560 3517.230 ;
        RECT 1090.300 3463.930 1090.560 3464.250 ;
        RECT 1095.360 3463.930 1095.620 3464.250 ;
        RECT 1090.360 3415.370 1090.500 3463.930 ;
        RECT 1090.360 3415.230 1091.420 3415.370 ;
        RECT 1091.280 3367.690 1091.420 3415.230 ;
        RECT 1090.300 3367.370 1090.560 3367.690 ;
        RECT 1091.220 3367.370 1091.480 3367.690 ;
        RECT 1090.360 3318.810 1090.500 3367.370 ;
        RECT 1090.360 3318.670 1091.420 3318.810 ;
        RECT 1091.280 3270.790 1091.420 3318.670 ;
        RECT 1090.300 3270.470 1090.560 3270.790 ;
        RECT 1091.220 3270.470 1091.480 3270.790 ;
        RECT 1090.360 3222.250 1090.500 3270.470 ;
        RECT 1090.360 3222.110 1091.420 3222.250 ;
        RECT 1091.280 3174.230 1091.420 3222.110 ;
        RECT 1090.300 3173.910 1090.560 3174.230 ;
        RECT 1091.220 3173.910 1091.480 3174.230 ;
        RECT 1090.360 3125.690 1090.500 3173.910 ;
        RECT 1090.360 3125.550 1091.420 3125.690 ;
        RECT 1091.280 3077.670 1091.420 3125.550 ;
        RECT 1090.300 3077.350 1090.560 3077.670 ;
        RECT 1091.220 3077.350 1091.480 3077.670 ;
        RECT 1090.360 3029.130 1090.500 3077.350 ;
        RECT 1090.360 3028.990 1091.420 3029.130 ;
        RECT 1091.280 2981.110 1091.420 3028.990 ;
        RECT 1090.300 2980.850 1090.560 2981.110 ;
        RECT 1090.300 2980.790 1090.960 2980.850 ;
        RECT 1091.220 2980.790 1091.480 2981.110 ;
        RECT 1090.360 2980.710 1090.960 2980.790 ;
        RECT 1090.820 2980.170 1090.960 2980.710 ;
        RECT 1090.820 2980.030 1091.420 2980.170 ;
        RECT 1091.280 2959.770 1091.420 2980.030 ;
        RECT 1090.820 2959.630 1091.420 2959.770 ;
        RECT 1090.820 2946.430 1090.960 2959.630 ;
        RECT 1090.760 2946.110 1091.020 2946.430 ;
        RECT 1090.300 2898.170 1090.560 2898.490 ;
        RECT 1090.360 2863.210 1090.500 2898.170 ;
        RECT 1090.360 2863.070 1090.960 2863.210 ;
        RECT 1090.820 2849.530 1090.960 2863.070 ;
        RECT 1090.760 2849.210 1091.020 2849.530 ;
        RECT 1091.680 2815.210 1091.940 2815.530 ;
        RECT 1091.740 2801.445 1091.880 2815.210 ;
        RECT 1090.750 2801.075 1091.030 2801.445 ;
        RECT 1091.670 2801.075 1091.950 2801.445 ;
        RECT 1090.820 2753.310 1090.960 2801.075 ;
        RECT 1090.760 2752.990 1091.020 2753.310 ;
        RECT 1092.140 2752.990 1092.400 2753.310 ;
        RECT 1092.200 2719.310 1092.340 2752.990 ;
        RECT 1092.140 2718.990 1092.400 2719.310 ;
        RECT 1091.680 2718.310 1091.940 2718.630 ;
        RECT 1091.740 2704.885 1091.880 2718.310 ;
        RECT 1090.750 2704.515 1091.030 2704.885 ;
        RECT 1091.670 2704.515 1091.950 2704.885 ;
        RECT 1090.820 2656.750 1090.960 2704.515 ;
        RECT 1090.760 2656.430 1091.020 2656.750 ;
        RECT 1092.140 2656.430 1092.400 2656.750 ;
        RECT 1092.200 2622.750 1092.340 2656.430 ;
        RECT 1092.140 2622.430 1092.400 2622.750 ;
        RECT 1091.680 2621.750 1091.940 2622.070 ;
        RECT 1091.740 2608.325 1091.880 2621.750 ;
        RECT 1090.750 2607.955 1091.030 2608.325 ;
        RECT 1091.670 2607.955 1091.950 2608.325 ;
        RECT 1090.820 2560.190 1090.960 2607.955 ;
        RECT 1090.760 2559.870 1091.020 2560.190 ;
        RECT 1092.140 2559.870 1092.400 2560.190 ;
        RECT 1092.200 2511.910 1092.340 2559.870 ;
        RECT 1091.220 2511.765 1091.480 2511.910 ;
        RECT 1089.830 2511.395 1090.110 2511.765 ;
        RECT 1091.210 2511.395 1091.490 2511.765 ;
        RECT 1092.140 2511.590 1092.400 2511.910 ;
        RECT 1089.900 2463.485 1090.040 2511.395 ;
        RECT 1089.830 2463.115 1090.110 2463.485 ;
        RECT 1090.750 2463.115 1091.030 2463.485 ;
        RECT 1090.820 2449.770 1090.960 2463.115 ;
        RECT 1090.820 2449.630 1091.420 2449.770 ;
        RECT 1091.280 2401.410 1091.420 2449.630 ;
        RECT 1090.300 2401.090 1090.560 2401.410 ;
        RECT 1091.220 2401.090 1091.480 2401.410 ;
        RECT 1090.360 2400.810 1090.500 2401.090 ;
        RECT 1090.360 2400.670 1090.960 2400.810 ;
        RECT 1090.820 2353.210 1090.960 2400.670 ;
        RECT 1090.820 2353.070 1091.420 2353.210 ;
        RECT 1091.280 2304.850 1091.420 2353.070 ;
        RECT 1090.300 2304.530 1090.560 2304.850 ;
        RECT 1091.220 2304.530 1091.480 2304.850 ;
        RECT 1090.360 2304.250 1090.500 2304.530 ;
        RECT 1090.360 2304.110 1090.960 2304.250 ;
        RECT 1090.820 2256.650 1090.960 2304.110 ;
        RECT 1090.820 2256.510 1091.420 2256.650 ;
        RECT 1091.280 2208.290 1091.420 2256.510 ;
        RECT 1090.300 2207.970 1090.560 2208.290 ;
        RECT 1091.220 2207.970 1091.480 2208.290 ;
        RECT 1090.360 2207.690 1090.500 2207.970 ;
        RECT 1090.360 2207.550 1090.960 2207.690 ;
        RECT 1090.820 2160.090 1090.960 2207.550 ;
        RECT 1090.820 2159.950 1091.420 2160.090 ;
        RECT 1091.280 2122.270 1091.420 2159.950 ;
        RECT 1028.660 2121.950 1028.920 2122.270 ;
        RECT 1091.220 2121.950 1091.480 2122.270 ;
        RECT 1028.720 2112.185 1028.860 2121.950 ;
        RECT 1028.720 2111.740 1029.070 2112.185 ;
        RECT 1028.790 2108.185 1029.070 2111.740 ;
      LAYER via2 ;
        RECT 1090.750 2801.120 1091.030 2801.400 ;
        RECT 1091.670 2801.120 1091.950 2801.400 ;
        RECT 1090.750 2704.560 1091.030 2704.840 ;
        RECT 1091.670 2704.560 1091.950 2704.840 ;
        RECT 1090.750 2608.000 1091.030 2608.280 ;
        RECT 1091.670 2608.000 1091.950 2608.280 ;
        RECT 1089.830 2511.440 1090.110 2511.720 ;
        RECT 1091.210 2511.440 1091.490 2511.720 ;
        RECT 1089.830 2463.160 1090.110 2463.440 ;
        RECT 1090.750 2463.160 1091.030 2463.440 ;
      LAYER met3 ;
        RECT 1090.725 2801.410 1091.055 2801.425 ;
        RECT 1091.645 2801.410 1091.975 2801.425 ;
        RECT 1090.725 2801.110 1091.975 2801.410 ;
        RECT 1090.725 2801.095 1091.055 2801.110 ;
        RECT 1091.645 2801.095 1091.975 2801.110 ;
        RECT 1090.725 2704.850 1091.055 2704.865 ;
        RECT 1091.645 2704.850 1091.975 2704.865 ;
        RECT 1090.725 2704.550 1091.975 2704.850 ;
        RECT 1090.725 2704.535 1091.055 2704.550 ;
        RECT 1091.645 2704.535 1091.975 2704.550 ;
        RECT 1090.725 2608.290 1091.055 2608.305 ;
        RECT 1091.645 2608.290 1091.975 2608.305 ;
        RECT 1090.725 2607.990 1091.975 2608.290 ;
        RECT 1090.725 2607.975 1091.055 2607.990 ;
        RECT 1091.645 2607.975 1091.975 2607.990 ;
        RECT 1089.805 2511.730 1090.135 2511.745 ;
        RECT 1091.185 2511.730 1091.515 2511.745 ;
        RECT 1089.805 2511.430 1091.515 2511.730 ;
        RECT 1089.805 2511.415 1090.135 2511.430 ;
        RECT 1091.185 2511.415 1091.515 2511.430 ;
        RECT 1089.805 2463.450 1090.135 2463.465 ;
        RECT 1090.725 2463.450 1091.055 2463.465 ;
        RECT 1089.805 2463.150 1091.055 2463.450 ;
        RECT 1089.805 2463.135 1090.135 2463.150 ;
        RECT 1090.725 2463.135 1091.055 2463.150 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
        RECT 771.565 2898.585 771.735 2946.355 ;
        RECT 772.025 2608.225 772.195 2656.335 ;
        RECT 772.025 2511.665 772.195 2559.775 ;
        RECT 772.025 2186.965 772.195 2221.815 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
        RECT 771.565 2946.185 771.735 2946.355 ;
        RECT 772.025 2656.165 772.195 2656.335 ;
        RECT 772.025 2559.605 772.195 2559.775 ;
        RECT 772.025 2221.645 772.195 2221.815 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 2981.020 771.810 2981.080 ;
        RECT 772.410 2981.020 772.730 2981.080 ;
        RECT 771.490 2980.880 772.730 2981.020 ;
        RECT 771.490 2980.820 771.810 2980.880 ;
        RECT 772.410 2980.820 772.730 2980.880 ;
        RECT 771.490 2946.340 771.810 2946.400 ;
        RECT 771.295 2946.200 771.810 2946.340 ;
        RECT 771.490 2946.140 771.810 2946.200 ;
        RECT 771.490 2898.740 771.810 2898.800 ;
        RECT 771.295 2898.600 771.810 2898.740 ;
        RECT 771.490 2898.540 771.810 2898.600 ;
        RECT 771.030 2898.060 771.350 2898.120 ;
        RECT 771.950 2898.060 772.270 2898.120 ;
        RECT 771.030 2897.920 772.270 2898.060 ;
        RECT 771.030 2897.860 771.350 2897.920 ;
        RECT 771.950 2897.860 772.270 2897.920 ;
        RECT 771.030 2814.760 771.350 2814.820 ;
        RECT 771.950 2814.760 772.270 2814.820 ;
        RECT 771.030 2814.620 772.270 2814.760 ;
        RECT 771.030 2814.560 771.350 2814.620 ;
        RECT 771.950 2814.560 772.270 2814.620 ;
        RECT 771.950 2656.320 772.270 2656.380 ;
        RECT 771.755 2656.180 772.270 2656.320 ;
        RECT 771.950 2656.120 772.270 2656.180 ;
        RECT 771.965 2608.380 772.255 2608.425 ;
        RECT 772.410 2608.380 772.730 2608.440 ;
        RECT 771.965 2608.240 772.730 2608.380 ;
        RECT 771.965 2608.195 772.255 2608.240 ;
        RECT 772.410 2608.180 772.730 2608.240 ;
        RECT 771.950 2559.760 772.270 2559.820 ;
        RECT 771.755 2559.620 772.270 2559.760 ;
        RECT 771.950 2559.560 772.270 2559.620 ;
        RECT 771.965 2511.820 772.255 2511.865 ;
        RECT 772.410 2511.820 772.730 2511.880 ;
        RECT 771.965 2511.680 772.730 2511.820 ;
        RECT 771.965 2511.635 772.255 2511.680 ;
        RECT 772.410 2511.620 772.730 2511.680 ;
        RECT 771.030 2463.200 771.350 2463.260 ;
        RECT 771.950 2463.200 772.270 2463.260 ;
        RECT 771.030 2463.060 772.270 2463.200 ;
        RECT 771.030 2463.000 771.350 2463.060 ;
        RECT 771.950 2463.000 772.270 2463.060 ;
        RECT 771.490 2332.300 771.810 2332.360 ;
        RECT 772.410 2332.300 772.730 2332.360 ;
        RECT 771.490 2332.160 772.730 2332.300 ;
        RECT 771.490 2332.100 771.810 2332.160 ;
        RECT 772.410 2332.100 772.730 2332.160 ;
        RECT 771.490 2235.540 771.810 2235.800 ;
        RECT 771.580 2235.400 771.720 2235.540 ;
        RECT 771.950 2235.400 772.270 2235.460 ;
        RECT 771.580 2235.260 772.270 2235.400 ;
        RECT 771.950 2235.200 772.270 2235.260 ;
        RECT 771.950 2221.800 772.270 2221.860 ;
        RECT 771.755 2221.660 772.270 2221.800 ;
        RECT 771.950 2221.600 772.270 2221.660 ;
        RECT 771.950 2187.120 772.270 2187.180 ;
        RECT 771.755 2186.980 772.270 2187.120 ;
        RECT 771.950 2186.920 772.270 2186.980 ;
        RECT 771.490 2125.580 771.810 2125.640 ;
        RECT 772.410 2125.580 772.730 2125.640 ;
        RECT 771.490 2125.440 772.730 2125.580 ;
        RECT 771.490 2125.380 771.810 2125.440 ;
        RECT 772.410 2125.380 772.730 2125.440 ;
        RECT 771.490 2122.180 771.810 2122.240 ;
        RECT 851.990 2122.180 852.310 2122.240 ;
        RECT 771.490 2122.040 852.310 2122.180 ;
        RECT 771.490 2121.980 771.810 2122.040 ;
        RECT 851.990 2121.980 852.310 2122.040 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 2980.820 771.780 2981.080 ;
        RECT 772.440 2980.820 772.700 2981.080 ;
        RECT 771.520 2946.140 771.780 2946.400 ;
        RECT 771.520 2898.540 771.780 2898.800 ;
        RECT 771.060 2897.860 771.320 2898.120 ;
        RECT 771.980 2897.860 772.240 2898.120 ;
        RECT 771.060 2814.560 771.320 2814.820 ;
        RECT 771.980 2814.560 772.240 2814.820 ;
        RECT 771.980 2656.120 772.240 2656.380 ;
        RECT 772.440 2608.180 772.700 2608.440 ;
        RECT 771.980 2559.560 772.240 2559.820 ;
        RECT 772.440 2511.620 772.700 2511.880 ;
        RECT 771.060 2463.000 771.320 2463.260 ;
        RECT 771.980 2463.000 772.240 2463.260 ;
        RECT 771.520 2332.100 771.780 2332.360 ;
        RECT 772.440 2332.100 772.700 2332.360 ;
        RECT 771.520 2235.540 771.780 2235.800 ;
        RECT 771.980 2235.200 772.240 2235.460 ;
        RECT 771.980 2221.600 772.240 2221.860 ;
        RECT 771.980 2186.920 772.240 2187.180 ;
        RECT 771.520 2125.380 771.780 2125.640 ;
        RECT 772.440 2125.380 772.700 2125.640 ;
        RECT 771.520 2121.980 771.780 2122.240 ;
        RECT 852.020 2121.980 852.280 2122.240 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 2981.110 771.720 3028.990 ;
        RECT 771.520 2980.790 771.780 2981.110 ;
        RECT 772.440 2980.850 772.700 2981.110 ;
        RECT 772.040 2980.790 772.700 2980.850 ;
        RECT 772.040 2980.710 772.640 2980.790 ;
        RECT 772.040 2959.770 772.180 2980.710 ;
        RECT 771.580 2959.630 772.180 2959.770 ;
        RECT 771.580 2946.430 771.720 2959.630 ;
        RECT 771.520 2946.110 771.780 2946.430 ;
        RECT 771.520 2898.570 771.780 2898.830 ;
        RECT 771.120 2898.510 771.780 2898.570 ;
        RECT 771.120 2898.430 771.720 2898.510 ;
        RECT 771.120 2898.150 771.260 2898.430 ;
        RECT 771.060 2897.830 771.320 2898.150 ;
        RECT 771.980 2897.830 772.240 2898.150 ;
        RECT 772.040 2814.850 772.180 2897.830 ;
        RECT 771.060 2814.530 771.320 2814.850 ;
        RECT 771.980 2814.530 772.240 2814.850 ;
        RECT 771.120 2766.650 771.260 2814.530 ;
        RECT 771.120 2766.510 771.720 2766.650 ;
        RECT 771.580 2719.050 771.720 2766.510 ;
        RECT 771.580 2718.910 772.640 2719.050 ;
        RECT 772.500 2670.090 772.640 2718.910 ;
        RECT 772.040 2669.950 772.640 2670.090 ;
        RECT 772.040 2656.410 772.180 2669.950 ;
        RECT 771.980 2656.090 772.240 2656.410 ;
        RECT 772.440 2608.150 772.700 2608.470 ;
        RECT 772.500 2573.530 772.640 2608.150 ;
        RECT 772.040 2573.390 772.640 2573.530 ;
        RECT 772.040 2559.850 772.180 2573.390 ;
        RECT 771.980 2559.530 772.240 2559.850 ;
        RECT 772.440 2511.590 772.700 2511.910 ;
        RECT 772.500 2476.970 772.640 2511.590 ;
        RECT 772.040 2476.830 772.640 2476.970 ;
        RECT 772.040 2463.290 772.180 2476.830 ;
        RECT 771.060 2462.970 771.320 2463.290 ;
        RECT 771.980 2462.970 772.240 2463.290 ;
        RECT 771.120 2415.205 771.260 2462.970 ;
        RECT 771.050 2414.835 771.330 2415.205 ;
        RECT 772.430 2414.835 772.710 2415.205 ;
        RECT 772.500 2380.410 772.640 2414.835 ;
        RECT 771.580 2380.270 772.640 2380.410 ;
        RECT 771.580 2332.390 771.720 2380.270 ;
        RECT 771.520 2332.070 771.780 2332.390 ;
        RECT 772.440 2332.070 772.700 2332.390 ;
        RECT 772.500 2283.850 772.640 2332.070 ;
        RECT 771.580 2283.710 772.640 2283.850 ;
        RECT 771.580 2235.830 771.720 2283.710 ;
        RECT 771.520 2235.510 771.780 2235.830 ;
        RECT 771.980 2235.170 772.240 2235.490 ;
        RECT 772.040 2221.890 772.180 2235.170 ;
        RECT 771.980 2221.570 772.240 2221.890 ;
        RECT 771.980 2186.890 772.240 2187.210 ;
        RECT 772.040 2173.690 772.180 2186.890 ;
        RECT 772.040 2173.550 772.640 2173.690 ;
        RECT 772.500 2125.670 772.640 2173.550 ;
        RECT 771.520 2125.350 771.780 2125.670 ;
        RECT 772.440 2125.350 772.700 2125.670 ;
        RECT 771.580 2122.270 771.720 2125.350 ;
        RECT 771.520 2121.950 771.780 2122.270 ;
        RECT 852.020 2121.950 852.280 2122.270 ;
        RECT 852.080 2112.185 852.220 2121.950 ;
        RECT 852.080 2111.740 852.430 2112.185 ;
        RECT 852.150 2108.185 852.430 2111.740 ;
      LAYER via2 ;
        RECT 771.050 2414.880 771.330 2415.160 ;
        RECT 772.430 2414.880 772.710 2415.160 ;
      LAYER met3 ;
        RECT 771.025 2415.170 771.355 2415.185 ;
        RECT 772.405 2415.170 772.735 2415.185 ;
        RECT 771.025 2414.870 772.735 2415.170 ;
        RECT 771.025 2414.855 771.355 2414.870 ;
        RECT 772.405 2414.855 772.735 2414.870 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2121.840 448.430 2121.900 ;
        RECT 674.890 2121.840 675.210 2121.900 ;
        RECT 448.110 2121.700 675.210 2121.840 ;
        RECT 448.110 2121.640 448.430 2121.700 ;
        RECT 674.890 2121.640 675.210 2121.700 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2121.640 448.400 2121.900 ;
        RECT 674.920 2121.640 675.180 2121.900 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2121.930 448.340 3498.270 ;
        RECT 448.140 2121.610 448.400 2121.930 ;
        RECT 674.920 2121.610 675.180 2121.930 ;
        RECT 674.980 2112.185 675.120 2121.610 ;
        RECT 674.980 2111.740 675.330 2112.185 ;
        RECT 675.050 2108.185 675.330 2111.740 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2122.180 124.130 2122.240 ;
        RECT 498.250 2122.180 498.570 2122.240 ;
        RECT 123.810 2122.040 498.570 2122.180 ;
        RECT 123.810 2121.980 124.130 2122.040 ;
        RECT 498.250 2121.980 498.570 2122.040 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2121.980 124.100 2122.240 ;
        RECT 498.280 2121.980 498.540 2122.240 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2122.270 124.040 3498.270 ;
        RECT 123.840 2121.950 124.100 2122.270 ;
        RECT 498.280 2121.950 498.540 2122.270 ;
        RECT 498.340 2112.185 498.480 2121.950 ;
        RECT 498.340 2111.740 498.690 2112.185 ;
        RECT 498.410 2108.185 498.690 2111.740 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2056.220 17.410 2056.280 ;
        RECT 393.370 2056.220 393.690 2056.280 ;
        RECT 17.090 2056.080 393.690 2056.220 ;
        RECT 17.090 2056.020 17.410 2056.080 ;
        RECT 393.370 2056.020 393.690 2056.080 ;
      LAYER via ;
        RECT 17.120 2056.020 17.380 2056.280 ;
        RECT 393.400 2056.020 393.660 2056.280 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 2056.310 17.320 3339.635 ;
        RECT 17.120 2055.990 17.380 2056.310 ;
        RECT 393.400 2055.990 393.660 2056.310 ;
        RECT 393.460 2054.805 393.600 2055.990 ;
        RECT 393.390 2054.435 393.670 2054.805 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 393.390 2054.480 393.670 2054.760 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 393.365 2054.770 393.695 2054.785 ;
        RECT 410.000 2054.770 414.000 2054.920 ;
        RECT 393.365 2054.470 414.000 2054.770 ;
        RECT 393.365 2054.455 393.695 2054.470 ;
        RECT 410.000 2054.320 414.000 2054.470 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1945.720 17.870 1945.780 ;
        RECT 393.370 1945.720 393.690 1945.780 ;
        RECT 17.550 1945.580 393.690 1945.720 ;
        RECT 17.550 1945.520 17.870 1945.580 ;
        RECT 393.370 1945.520 393.690 1945.580 ;
      LAYER via ;
        RECT 17.580 1945.520 17.840 1945.780 ;
        RECT 393.400 1945.520 393.660 1945.780 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 1945.810 17.780 3051.995 ;
        RECT 17.580 1945.490 17.840 1945.810 ;
        RECT 393.400 1945.490 393.660 1945.810 ;
        RECT 393.460 1940.565 393.600 1945.490 ;
        RECT 393.390 1940.195 393.670 1940.565 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 393.390 1940.240 393.670 1940.520 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 393.365 1940.530 393.695 1940.545 ;
        RECT 410.000 1940.530 414.000 1940.680 ;
        RECT 393.365 1940.230 414.000 1940.530 ;
        RECT 393.365 1940.215 393.695 1940.230 ;
        RECT 410.000 1940.080 414.000 1940.230 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 1828.420 18.330 1828.480 ;
        RECT 393.370 1828.420 393.690 1828.480 ;
        RECT 18.010 1828.280 393.690 1828.420 ;
        RECT 18.010 1828.220 18.330 1828.280 ;
        RECT 393.370 1828.220 393.690 1828.280 ;
      LAYER via ;
        RECT 18.040 1828.220 18.300 1828.480 ;
        RECT 393.400 1828.220 393.660 1828.480 ;
      LAYER met2 ;
        RECT 18.030 2765.035 18.310 2765.405 ;
        RECT 18.100 1828.510 18.240 2765.035 ;
        RECT 18.040 1828.190 18.300 1828.510 ;
        RECT 393.400 1828.190 393.660 1828.510 ;
        RECT 393.460 1826.325 393.600 1828.190 ;
        RECT 393.390 1825.955 393.670 1826.325 ;
      LAYER via2 ;
        RECT 18.030 2765.080 18.310 2765.360 ;
        RECT 393.390 1826.000 393.670 1826.280 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.005 2765.370 18.335 2765.385 ;
        RECT -4.800 2765.070 18.335 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.005 2765.055 18.335 2765.070 ;
        RECT 393.365 1826.290 393.695 1826.305 ;
        RECT 410.000 1826.290 414.000 1826.440 ;
        RECT 393.365 1825.990 414.000 1826.290 ;
        RECT 393.365 1825.975 393.695 1825.990 ;
        RECT 410.000 1825.840 414.000 1825.990 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 1717.920 18.790 1717.980 ;
        RECT 393.370 1717.920 393.690 1717.980 ;
        RECT 18.470 1717.780 393.690 1717.920 ;
        RECT 18.470 1717.720 18.790 1717.780 ;
        RECT 393.370 1717.720 393.690 1717.780 ;
      LAYER via ;
        RECT 18.500 1717.720 18.760 1717.980 ;
        RECT 393.400 1717.720 393.660 1717.980 ;
      LAYER met2 ;
        RECT 18.490 2477.395 18.770 2477.765 ;
        RECT 18.560 1718.010 18.700 2477.395 ;
        RECT 18.500 1717.690 18.760 1718.010 ;
        RECT 393.400 1717.690 393.660 1718.010 ;
        RECT 393.460 1711.405 393.600 1717.690 ;
        RECT 393.390 1711.035 393.670 1711.405 ;
      LAYER via2 ;
        RECT 18.490 2477.440 18.770 2477.720 ;
        RECT 393.390 1711.080 393.670 1711.360 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 18.465 2477.730 18.795 2477.745 ;
        RECT -4.800 2477.430 18.795 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 18.465 2477.415 18.795 2477.430 ;
        RECT 393.365 1711.370 393.695 1711.385 ;
        RECT 410.000 1711.370 414.000 1711.520 ;
        RECT 393.365 1711.070 414.000 1711.370 ;
        RECT 393.365 1711.055 393.695 1711.070 ;
        RECT 410.000 1710.920 414.000 1711.070 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 1600.620 19.250 1600.680 ;
        RECT 393.370 1600.620 393.690 1600.680 ;
        RECT 18.930 1600.480 393.690 1600.620 ;
        RECT 18.930 1600.420 19.250 1600.480 ;
        RECT 393.370 1600.420 393.690 1600.480 ;
      LAYER via ;
        RECT 18.960 1600.420 19.220 1600.680 ;
        RECT 393.400 1600.420 393.660 1600.680 ;
      LAYER met2 ;
        RECT 18.950 2189.755 19.230 2190.125 ;
        RECT 19.020 1600.710 19.160 2189.755 ;
        RECT 18.960 1600.390 19.220 1600.710 ;
        RECT 393.400 1600.390 393.660 1600.710 ;
        RECT 393.460 1597.165 393.600 1600.390 ;
        RECT 393.390 1596.795 393.670 1597.165 ;
      LAYER via2 ;
        RECT 18.950 2189.800 19.230 2190.080 ;
        RECT 393.390 1596.840 393.670 1597.120 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.925 2190.090 19.255 2190.105 ;
        RECT -4.800 2189.790 19.255 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.925 2189.775 19.255 2189.790 ;
        RECT 393.365 1597.130 393.695 1597.145 ;
        RECT 410.000 1597.130 414.000 1597.280 ;
        RECT 393.365 1596.830 414.000 1597.130 ;
        RECT 393.365 1596.815 393.695 1596.830 ;
        RECT 410.000 1596.680 414.000 1596.830 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1483.320 17.410 1483.380 ;
        RECT 393.370 1483.320 393.690 1483.380 ;
        RECT 17.090 1483.180 393.690 1483.320 ;
        RECT 17.090 1483.120 17.410 1483.180 ;
        RECT 393.370 1483.120 393.690 1483.180 ;
      LAYER via ;
        RECT 17.120 1483.120 17.380 1483.380 ;
        RECT 393.400 1483.120 393.660 1483.380 ;
      LAYER met2 ;
        RECT 17.110 1902.795 17.390 1903.165 ;
        RECT 17.180 1483.410 17.320 1902.795 ;
        RECT 17.120 1483.090 17.380 1483.410 ;
        RECT 393.400 1483.090 393.660 1483.410 ;
        RECT 393.460 1482.925 393.600 1483.090 ;
        RECT 393.390 1482.555 393.670 1482.925 ;
      LAYER via2 ;
        RECT 17.110 1902.840 17.390 1903.120 ;
        RECT 393.390 1482.600 393.670 1482.880 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.085 1903.130 17.415 1903.145 ;
        RECT -4.800 1902.830 17.415 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.085 1902.815 17.415 1902.830 ;
        RECT 393.365 1482.890 393.695 1482.905 ;
        RECT 410.000 1482.890 414.000 1483.040 ;
        RECT 393.365 1482.590 414.000 1482.890 ;
        RECT 393.365 1482.575 393.695 1482.590 ;
        RECT 410.000 1482.440 414.000 1482.590 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.190 620.740 2011.510 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2011.190 620.600 2901.150 620.740 ;
        RECT 2011.190 620.540 2011.510 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2011.220 620.540 2011.480 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2011.210 776.715 2011.490 777.085 ;
        RECT 2011.280 620.830 2011.420 776.715 ;
        RECT 2011.220 620.510 2011.480 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2011.210 776.760 2011.490 777.040 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 1997.465 777.050 2001.465 777.200 ;
        RECT 2011.185 777.050 2011.515 777.065 ;
        RECT 1997.465 776.750 2011.515 777.050 ;
        RECT 1997.465 776.600 2001.465 776.750 ;
        RECT 2011.185 776.735 2011.515 776.750 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 1373.160 18.330 1373.220 ;
        RECT 393.370 1373.160 393.690 1373.220 ;
        RECT 18.010 1373.020 393.690 1373.160 ;
        RECT 18.010 1372.960 18.330 1373.020 ;
        RECT 393.370 1372.960 393.690 1373.020 ;
      LAYER via ;
        RECT 18.040 1372.960 18.300 1373.220 ;
        RECT 393.400 1372.960 393.660 1373.220 ;
      LAYER met2 ;
        RECT 18.030 1615.155 18.310 1615.525 ;
        RECT 18.100 1373.250 18.240 1615.155 ;
        RECT 18.040 1372.930 18.300 1373.250 ;
        RECT 393.400 1372.930 393.660 1373.250 ;
        RECT 393.460 1368.685 393.600 1372.930 ;
        RECT 393.390 1368.315 393.670 1368.685 ;
      LAYER via2 ;
        RECT 18.030 1615.200 18.310 1615.480 ;
        RECT 393.390 1368.360 393.670 1368.640 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 18.005 1615.490 18.335 1615.505 ;
        RECT -4.800 1615.190 18.335 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 18.005 1615.175 18.335 1615.190 ;
        RECT 393.365 1368.650 393.695 1368.665 ;
        RECT 410.000 1368.650 414.000 1368.800 ;
        RECT 393.365 1368.350 414.000 1368.650 ;
        RECT 393.365 1368.335 393.695 1368.350 ;
        RECT 410.000 1368.200 414.000 1368.350 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1255.860 17.870 1255.920 ;
        RECT 393.370 1255.860 393.690 1255.920 ;
        RECT 17.550 1255.720 393.690 1255.860 ;
        RECT 17.550 1255.660 17.870 1255.720 ;
        RECT 393.370 1255.660 393.690 1255.720 ;
      LAYER via ;
        RECT 17.580 1255.660 17.840 1255.920 ;
        RECT 393.400 1255.660 393.660 1255.920 ;
      LAYER met2 ;
        RECT 17.570 1400.275 17.850 1400.645 ;
        RECT 17.640 1255.950 17.780 1400.275 ;
        RECT 17.580 1255.630 17.840 1255.950 ;
        RECT 393.400 1255.630 393.660 1255.950 ;
        RECT 393.460 1253.765 393.600 1255.630 ;
        RECT 393.390 1253.395 393.670 1253.765 ;
      LAYER via2 ;
        RECT 17.570 1400.320 17.850 1400.600 ;
        RECT 393.390 1253.440 393.670 1253.720 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.545 1400.610 17.875 1400.625 ;
        RECT -4.800 1400.310 17.875 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.545 1400.295 17.875 1400.310 ;
        RECT 393.365 1253.730 393.695 1253.745 ;
        RECT 410.000 1253.730 414.000 1253.880 ;
        RECT 393.365 1253.430 414.000 1253.730 ;
        RECT 393.365 1253.415 393.695 1253.430 ;
        RECT 410.000 1253.280 414.000 1253.430 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1145.360 17.870 1145.420 ;
        RECT 393.370 1145.360 393.690 1145.420 ;
        RECT 17.550 1145.220 393.690 1145.360 ;
        RECT 17.550 1145.160 17.870 1145.220 ;
        RECT 393.370 1145.160 393.690 1145.220 ;
      LAYER via ;
        RECT 17.580 1145.160 17.840 1145.420 ;
        RECT 393.400 1145.160 393.660 1145.420 ;
      LAYER met2 ;
        RECT 17.570 1184.715 17.850 1185.085 ;
        RECT 17.640 1145.450 17.780 1184.715 ;
        RECT 17.580 1145.130 17.840 1145.450 ;
        RECT 393.400 1145.130 393.660 1145.450 ;
        RECT 393.460 1139.525 393.600 1145.130 ;
        RECT 393.390 1139.155 393.670 1139.525 ;
      LAYER via2 ;
        RECT 17.570 1184.760 17.850 1185.040 ;
        RECT 393.390 1139.200 393.670 1139.480 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.545 1185.050 17.875 1185.065 ;
        RECT -4.800 1184.750 17.875 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.545 1184.735 17.875 1184.750 ;
        RECT 393.365 1139.490 393.695 1139.505 ;
        RECT 410.000 1139.490 414.000 1139.640 ;
        RECT 393.365 1139.190 414.000 1139.490 ;
        RECT 393.365 1139.175 393.695 1139.190 ;
        RECT 410.000 1139.040 414.000 1139.190 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 396.590 972.640 396.910 972.700 ;
        RECT 15.710 972.500 396.910 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 396.590 972.440 396.910 972.500 ;
      LAYER via ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 396.620 972.440 396.880 972.700 ;
      LAYER met2 ;
        RECT 396.610 1024.915 396.890 1025.285 ;
        RECT 396.680 972.730 396.820 1024.915 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 396.620 972.410 396.880 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 396.610 1024.960 396.890 1025.240 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 396.585 1025.250 396.915 1025.265 ;
        RECT 410.000 1025.250 414.000 1025.400 ;
        RECT 396.585 1024.950 414.000 1025.250 ;
        RECT 396.585 1024.935 396.915 1024.950 ;
        RECT 410.000 1024.800 414.000 1024.950 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 397.510 758.780 397.830 758.840 ;
        RECT 15.710 758.640 397.830 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 397.510 758.580 397.830 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 397.540 758.580 397.800 758.840 ;
      LAYER met2 ;
        RECT 397.530 909.995 397.810 910.365 ;
        RECT 397.600 758.870 397.740 909.995 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 397.540 758.550 397.800 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 397.530 910.040 397.810 910.320 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 397.505 910.330 397.835 910.345 ;
        RECT 410.000 910.330 414.000 910.480 ;
        RECT 397.505 910.030 414.000 910.330 ;
        RECT 397.505 910.015 397.835 910.030 ;
        RECT 410.000 909.880 414.000 910.030 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 396.590 544.920 396.910 544.980 ;
        RECT 16.170 544.780 396.910 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 396.590 544.720 396.910 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 396.620 544.720 396.880 544.980 ;
      LAYER met2 ;
        RECT 396.610 795.755 396.890 796.125 ;
        RECT 396.680 545.010 396.820 795.755 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 396.620 544.690 396.880 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 396.610 795.800 396.890 796.080 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 396.585 796.090 396.915 796.105 ;
        RECT 410.000 796.090 414.000 796.240 ;
        RECT 396.585 795.790 414.000 796.090 ;
        RECT 396.585 795.775 396.915 795.790 ;
        RECT 410.000 795.640 414.000 795.790 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 397.970 324.260 398.290 324.320 ;
        RECT 16.630 324.120 398.290 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 397.970 324.060 398.290 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 398.000 324.060 398.260 324.320 ;
      LAYER met2 ;
        RECT 397.990 681.515 398.270 681.885 ;
        RECT 398.060 324.350 398.200 681.515 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 398.000 324.030 398.260 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 397.990 681.560 398.270 681.840 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 397.965 681.850 398.295 681.865 ;
        RECT 410.000 681.850 414.000 682.000 ;
        RECT 397.965 681.550 414.000 681.850 ;
        RECT 397.965 681.535 398.295 681.550 ;
        RECT 410.000 681.400 414.000 681.550 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 397.050 110.400 397.370 110.460 ;
        RECT 15.710 110.260 397.370 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 397.050 110.200 397.370 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 397.080 110.200 397.340 110.460 ;
      LAYER met2 ;
        RECT 397.070 567.275 397.350 567.645 ;
        RECT 397.140 110.490 397.280 567.275 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 397.080 110.170 397.340 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 397.070 567.320 397.350 567.600 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 397.045 567.610 397.375 567.625 ;
        RECT 410.000 567.610 414.000 567.760 ;
        RECT 397.045 567.310 414.000 567.610 ;
        RECT 397.045 567.295 397.375 567.310 ;
        RECT 410.000 567.160 414.000 567.310 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2011.190 855.340 2011.510 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2011.190 855.200 2901.150 855.340 ;
        RECT 2011.190 855.140 2011.510 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2011.220 855.140 2011.480 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2011.210 883.475 2011.490 883.845 ;
        RECT 2011.280 855.430 2011.420 883.475 ;
        RECT 2011.220 855.110 2011.480 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2011.210 883.520 2011.490 883.800 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 1997.465 883.810 2001.465 883.960 ;
        RECT 2011.185 883.810 2011.515 883.825 ;
        RECT 1997.465 883.510 2011.515 883.810 ;
        RECT 1997.465 883.360 2001.465 883.510 ;
        RECT 2011.185 883.495 2011.515 883.510 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 993.380 2008.290 993.440 ;
        RECT 2901.290 993.380 2901.610 993.440 ;
        RECT 2007.970 993.240 2901.610 993.380 ;
        RECT 2007.970 993.180 2008.290 993.240 ;
        RECT 2901.290 993.180 2901.610 993.240 ;
      LAYER via ;
        RECT 2008.000 993.180 2008.260 993.440 ;
        RECT 2901.320 993.180 2901.580 993.440 ;
      LAYER met2 ;
        RECT 2901.310 1084.755 2901.590 1085.125 ;
        RECT 2901.380 993.470 2901.520 1084.755 ;
        RECT 2008.000 993.150 2008.260 993.470 ;
        RECT 2901.320 993.150 2901.580 993.470 ;
        RECT 2008.060 990.605 2008.200 993.150 ;
        RECT 2007.990 990.235 2008.270 990.605 ;
      LAYER via2 ;
        RECT 2901.310 1084.800 2901.590 1085.080 ;
        RECT 2007.990 990.280 2008.270 990.560 ;
      LAYER met3 ;
        RECT 2901.285 1085.090 2901.615 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2901.285 1084.790 2924.800 1085.090 ;
        RECT 2901.285 1084.775 2901.615 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 1997.465 990.570 2001.465 990.720 ;
        RECT 2007.965 990.570 2008.295 990.585 ;
        RECT 1997.465 990.270 2008.295 990.570 ;
        RECT 1997.465 990.120 2001.465 990.270 ;
        RECT 2007.965 990.255 2008.295 990.270 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2038.790 1318.080 2039.110 1318.140 ;
        RECT 2898.990 1318.080 2899.310 1318.140 ;
        RECT 2038.790 1317.940 2899.310 1318.080 ;
        RECT 2038.790 1317.880 2039.110 1317.940 ;
        RECT 2898.990 1317.880 2899.310 1317.940 ;
        RECT 2007.970 1103.880 2008.290 1103.940 ;
        RECT 2038.790 1103.880 2039.110 1103.940 ;
        RECT 2007.970 1103.740 2039.110 1103.880 ;
        RECT 2007.970 1103.680 2008.290 1103.740 ;
        RECT 2038.790 1103.680 2039.110 1103.740 ;
      LAYER via ;
        RECT 2038.820 1317.880 2039.080 1318.140 ;
        RECT 2899.020 1317.880 2899.280 1318.140 ;
        RECT 2008.000 1103.680 2008.260 1103.940 ;
        RECT 2038.820 1103.680 2039.080 1103.940 ;
      LAYER met2 ;
        RECT 2899.010 1319.355 2899.290 1319.725 ;
        RECT 2899.080 1318.170 2899.220 1319.355 ;
        RECT 2038.820 1317.850 2039.080 1318.170 ;
        RECT 2899.020 1317.850 2899.280 1318.170 ;
        RECT 2038.880 1103.970 2039.020 1317.850 ;
        RECT 2008.000 1103.650 2008.260 1103.970 ;
        RECT 2038.820 1103.650 2039.080 1103.970 ;
        RECT 2008.060 1097.365 2008.200 1103.650 ;
        RECT 2007.990 1096.995 2008.270 1097.365 ;
      LAYER via2 ;
        RECT 2899.010 1319.400 2899.290 1319.680 ;
        RECT 2007.990 1097.040 2008.270 1097.320 ;
      LAYER met3 ;
        RECT 2898.985 1319.690 2899.315 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2898.985 1319.390 2924.800 1319.690 ;
        RECT 2898.985 1319.375 2899.315 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 1997.465 1097.330 2001.465 1097.480 ;
        RECT 2007.965 1097.330 2008.295 1097.345 ;
        RECT 1997.465 1097.030 2008.295 1097.330 ;
        RECT 1997.465 1096.880 2001.465 1097.030 ;
        RECT 2007.965 1097.015 2008.295 1097.030 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2045.690 1552.680 2046.010 1552.740 ;
        RECT 2898.070 1552.680 2898.390 1552.740 ;
        RECT 2045.690 1552.540 2898.390 1552.680 ;
        RECT 2045.690 1552.480 2046.010 1552.540 ;
        RECT 2898.070 1552.480 2898.390 1552.540 ;
        RECT 2007.970 1207.240 2008.290 1207.300 ;
        RECT 2045.690 1207.240 2046.010 1207.300 ;
        RECT 2007.970 1207.100 2046.010 1207.240 ;
        RECT 2007.970 1207.040 2008.290 1207.100 ;
        RECT 2045.690 1207.040 2046.010 1207.100 ;
      LAYER via ;
        RECT 2045.720 1552.480 2045.980 1552.740 ;
        RECT 2898.100 1552.480 2898.360 1552.740 ;
        RECT 2008.000 1207.040 2008.260 1207.300 ;
        RECT 2045.720 1207.040 2045.980 1207.300 ;
      LAYER met2 ;
        RECT 2898.090 1553.955 2898.370 1554.325 ;
        RECT 2898.160 1552.770 2898.300 1553.955 ;
        RECT 2045.720 1552.450 2045.980 1552.770 ;
        RECT 2898.100 1552.450 2898.360 1552.770 ;
        RECT 2045.780 1207.330 2045.920 1552.450 ;
        RECT 2008.000 1207.010 2008.260 1207.330 ;
        RECT 2045.720 1207.010 2045.980 1207.330 ;
        RECT 2008.060 1204.125 2008.200 1207.010 ;
        RECT 2007.990 1203.755 2008.270 1204.125 ;
      LAYER via2 ;
        RECT 2898.090 1554.000 2898.370 1554.280 ;
        RECT 2007.990 1203.800 2008.270 1204.080 ;
      LAYER met3 ;
        RECT 2898.065 1554.290 2898.395 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2898.065 1553.990 2924.800 1554.290 ;
        RECT 2898.065 1553.975 2898.395 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 1997.465 1204.090 2001.465 1204.240 ;
        RECT 2007.965 1204.090 2008.295 1204.105 ;
        RECT 1997.465 1203.790 2008.295 1204.090 ;
        RECT 1997.465 1203.640 2001.465 1203.790 ;
        RECT 2007.965 1203.775 2008.295 1203.790 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2024.990 1787.280 2025.310 1787.340 ;
        RECT 2899.450 1787.280 2899.770 1787.340 ;
        RECT 2024.990 1787.140 2899.770 1787.280 ;
        RECT 2024.990 1787.080 2025.310 1787.140 ;
        RECT 2899.450 1787.080 2899.770 1787.140 ;
        RECT 2007.970 1310.940 2008.290 1311.000 ;
        RECT 2024.990 1310.940 2025.310 1311.000 ;
        RECT 2007.970 1310.800 2025.310 1310.940 ;
        RECT 2007.970 1310.740 2008.290 1310.800 ;
        RECT 2024.990 1310.740 2025.310 1310.800 ;
      LAYER via ;
        RECT 2025.020 1787.080 2025.280 1787.340 ;
        RECT 2899.480 1787.080 2899.740 1787.340 ;
        RECT 2008.000 1310.740 2008.260 1311.000 ;
        RECT 2025.020 1310.740 2025.280 1311.000 ;
      LAYER met2 ;
        RECT 2899.470 1789.235 2899.750 1789.605 ;
        RECT 2899.540 1787.370 2899.680 1789.235 ;
        RECT 2025.020 1787.050 2025.280 1787.370 ;
        RECT 2899.480 1787.050 2899.740 1787.370 ;
        RECT 2025.080 1311.030 2025.220 1787.050 ;
        RECT 2008.000 1310.885 2008.260 1311.030 ;
        RECT 2007.990 1310.515 2008.270 1310.885 ;
        RECT 2025.020 1310.710 2025.280 1311.030 ;
      LAYER via2 ;
        RECT 2899.470 1789.280 2899.750 1789.560 ;
        RECT 2007.990 1310.560 2008.270 1310.840 ;
      LAYER met3 ;
        RECT 2899.445 1789.570 2899.775 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2899.445 1789.270 2924.800 1789.570 ;
        RECT 2899.445 1789.255 2899.775 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 1997.465 1310.850 2001.465 1311.000 ;
        RECT 2007.965 1310.850 2008.295 1310.865 ;
        RECT 1997.465 1310.550 2008.295 1310.850 ;
        RECT 1997.465 1310.400 2001.465 1310.550 ;
        RECT 2007.965 1310.535 2008.295 1310.550 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 1421.440 2008.290 1421.500 ;
        RECT 2901.290 1421.440 2901.610 1421.500 ;
        RECT 2007.970 1421.300 2901.610 1421.440 ;
        RECT 2007.970 1421.240 2008.290 1421.300 ;
        RECT 2901.290 1421.240 2901.610 1421.300 ;
      LAYER via ;
        RECT 2008.000 1421.240 2008.260 1421.500 ;
        RECT 2901.320 1421.240 2901.580 1421.500 ;
      LAYER met2 ;
        RECT 2901.310 2023.835 2901.590 2024.205 ;
        RECT 2901.380 1421.530 2901.520 2023.835 ;
        RECT 2008.000 1421.210 2008.260 1421.530 ;
        RECT 2901.320 1421.210 2901.580 1421.530 ;
        RECT 2008.060 1417.645 2008.200 1421.210 ;
        RECT 2007.990 1417.275 2008.270 1417.645 ;
      LAYER via2 ;
        RECT 2901.310 2023.880 2901.590 2024.160 ;
        RECT 2007.990 1417.320 2008.270 1417.600 ;
      LAYER met3 ;
        RECT 2901.285 2024.170 2901.615 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.285 2023.870 2924.800 2024.170 ;
        RECT 2901.285 2023.855 2901.615 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 1997.465 1417.610 2001.465 1417.760 ;
        RECT 2007.965 1417.610 2008.295 1417.625 ;
        RECT 1997.465 1417.310 2008.295 1417.610 ;
        RECT 1997.465 1417.160 2001.465 1417.310 ;
        RECT 2007.965 1417.295 2008.295 1417.310 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 1524.800 2008.290 1524.860 ;
        RECT 2901.750 1524.800 2902.070 1524.860 ;
        RECT 2007.970 1524.660 2902.070 1524.800 ;
        RECT 2007.970 1524.600 2008.290 1524.660 ;
        RECT 2901.750 1524.600 2902.070 1524.660 ;
      LAYER via ;
        RECT 2008.000 1524.600 2008.260 1524.860 ;
        RECT 2901.780 1524.600 2902.040 1524.860 ;
      LAYER met2 ;
        RECT 2901.770 2258.435 2902.050 2258.805 ;
        RECT 2901.840 1524.890 2901.980 2258.435 ;
        RECT 2008.000 1524.570 2008.260 1524.890 ;
        RECT 2901.780 1524.570 2902.040 1524.890 ;
        RECT 2008.060 1524.405 2008.200 1524.570 ;
        RECT 2007.990 1524.035 2008.270 1524.405 ;
      LAYER via2 ;
        RECT 2901.770 2258.480 2902.050 2258.760 ;
        RECT 2007.990 1524.080 2008.270 1524.360 ;
      LAYER met3 ;
        RECT 2901.745 2258.770 2902.075 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2901.745 2258.470 2924.800 2258.770 ;
        RECT 2901.745 2258.455 2902.075 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 1997.465 1524.370 2001.465 1524.520 ;
        RECT 2007.965 1524.370 2008.295 1524.385 ;
        RECT 1997.465 1524.070 2008.295 1524.370 ;
        RECT 1997.465 1523.920 2001.465 1524.070 ;
        RECT 2007.965 1524.055 2008.295 1524.070 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 24.380 420.830 24.440 ;
        RECT 633.030 24.380 633.350 24.440 ;
        RECT 420.510 24.240 633.350 24.380 ;
        RECT 420.510 24.180 420.830 24.240 ;
        RECT 633.030 24.180 633.350 24.240 ;
      LAYER via ;
        RECT 420.540 24.180 420.800 24.440 ;
        RECT 633.060 24.180 633.320 24.440 ;
      LAYER met2 ;
        RECT 419.750 510.410 420.030 514.000 ;
        RECT 419.750 510.270 420.740 510.410 ;
        RECT 419.750 510.000 420.030 510.270 ;
        RECT 420.600 24.470 420.740 510.270 ;
        RECT 420.540 24.150 420.800 24.470 ;
        RECT 633.060 24.150 633.320 24.470 ;
        RECT 633.120 2.400 633.260 24.150 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1656.990 500.380 1657.310 500.440 ;
        RECT 2100.890 500.380 2101.210 500.440 ;
        RECT 1656.990 500.240 2101.210 500.380 ;
        RECT 1656.990 500.180 1657.310 500.240 ;
        RECT 2100.890 500.180 2101.210 500.240 ;
        RECT 2100.890 24.380 2101.210 24.440 ;
        RECT 2417.370 24.380 2417.690 24.440 ;
        RECT 2100.890 24.240 2417.690 24.380 ;
        RECT 2100.890 24.180 2101.210 24.240 ;
        RECT 2417.370 24.180 2417.690 24.240 ;
      LAYER via ;
        RECT 1657.020 500.180 1657.280 500.440 ;
        RECT 2100.920 500.180 2101.180 500.440 ;
        RECT 2100.920 24.180 2101.180 24.440 ;
        RECT 2417.400 24.180 2417.660 24.440 ;
      LAYER met2 ;
        RECT 1657.150 510.340 1657.430 514.000 ;
        RECT 1657.080 510.000 1657.430 510.340 ;
        RECT 1657.080 500.470 1657.220 510.000 ;
        RECT 1657.020 500.150 1657.280 500.470 ;
        RECT 2100.920 500.150 2101.180 500.470 ;
        RECT 2100.980 24.470 2101.120 500.150 ;
        RECT 2100.920 24.150 2101.180 24.470 ;
        RECT 2417.400 24.150 2417.660 24.470 ;
        RECT 2417.460 2.400 2417.600 24.150 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.490 493.240 1668.810 493.300 ;
        RECT 2428.870 493.240 2429.190 493.300 ;
        RECT 1668.490 493.100 2429.190 493.240 ;
        RECT 1668.490 493.040 1668.810 493.100 ;
        RECT 2428.870 493.040 2429.190 493.100 ;
        RECT 2428.870 37.640 2429.190 37.700 ;
        RECT 2434.850 37.640 2435.170 37.700 ;
        RECT 2428.870 37.500 2435.170 37.640 ;
        RECT 2428.870 37.440 2429.190 37.500 ;
        RECT 2434.850 37.440 2435.170 37.500 ;
      LAYER via ;
        RECT 1668.520 493.040 1668.780 493.300 ;
        RECT 2428.900 493.040 2429.160 493.300 ;
        RECT 2428.900 37.440 2429.160 37.700 ;
        RECT 2434.880 37.440 2435.140 37.700 ;
      LAYER met2 ;
        RECT 1669.110 510.410 1669.390 514.000 ;
        RECT 1668.580 510.270 1669.390 510.410 ;
        RECT 1668.580 493.330 1668.720 510.270 ;
        RECT 1669.110 510.000 1669.390 510.270 ;
        RECT 1668.520 493.010 1668.780 493.330 ;
        RECT 2428.900 493.010 2429.160 493.330 ;
        RECT 2428.960 37.730 2429.100 493.010 ;
        RECT 2428.900 37.410 2429.160 37.730 ;
        RECT 2434.880 37.410 2435.140 37.730 ;
        RECT 2434.940 2.400 2435.080 37.410 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 31.180 1683.530 31.240 ;
        RECT 2452.790 31.180 2453.110 31.240 ;
        RECT 1683.210 31.040 2453.110 31.180 ;
        RECT 1683.210 30.980 1683.530 31.040 ;
        RECT 2452.790 30.980 2453.110 31.040 ;
      LAYER via ;
        RECT 1683.240 30.980 1683.500 31.240 ;
        RECT 2452.820 30.980 2453.080 31.240 ;
      LAYER met2 ;
        RECT 1681.530 510.410 1681.810 514.000 ;
        RECT 1681.530 510.270 1683.440 510.410 ;
        RECT 1681.530 510.000 1681.810 510.270 ;
        RECT 1683.300 31.270 1683.440 510.270 ;
        RECT 1683.240 30.950 1683.500 31.270 ;
        RECT 2452.820 30.950 2453.080 31.270 ;
        RECT 2452.880 2.400 2453.020 30.950 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2470.730 38.660 2471.050 38.720 ;
        RECT 2449.660 38.520 2471.050 38.660 ;
        RECT 1697.010 38.320 1697.330 38.380 ;
        RECT 2449.660 38.320 2449.800 38.520 ;
        RECT 2470.730 38.460 2471.050 38.520 ;
        RECT 1697.010 38.180 2449.800 38.320 ;
        RECT 1697.010 38.120 1697.330 38.180 ;
      LAYER via ;
        RECT 1697.040 38.120 1697.300 38.380 ;
        RECT 2470.760 38.460 2471.020 38.720 ;
      LAYER met2 ;
        RECT 1693.950 510.410 1694.230 514.000 ;
        RECT 1693.950 510.270 1697.240 510.410 ;
        RECT 1693.950 510.000 1694.230 510.270 ;
        RECT 1697.100 38.410 1697.240 510.270 ;
        RECT 2470.760 38.430 2471.020 38.750 ;
        RECT 1697.040 38.090 1697.300 38.410 ;
        RECT 2470.820 2.400 2470.960 38.430 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1706.210 486.440 1706.530 486.500 ;
        RECT 2484.070 486.440 2484.390 486.500 ;
        RECT 1706.210 486.300 2484.390 486.440 ;
        RECT 1706.210 486.240 1706.530 486.300 ;
        RECT 2484.070 486.240 2484.390 486.300 ;
      LAYER via ;
        RECT 1706.240 486.240 1706.500 486.500 ;
        RECT 2484.100 486.240 2484.360 486.500 ;
      LAYER met2 ;
        RECT 1706.370 510.340 1706.650 514.000 ;
        RECT 1706.300 510.000 1706.650 510.340 ;
        RECT 1706.300 486.530 1706.440 510.000 ;
        RECT 1706.240 486.210 1706.500 486.530 ;
        RECT 2484.100 486.210 2484.360 486.530 ;
        RECT 2484.160 17.410 2484.300 486.210 ;
        RECT 2484.160 17.270 2488.900 17.410 ;
        RECT 2488.760 2.400 2488.900 17.270 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.630 479.640 1718.950 479.700 ;
        RECT 2504.770 479.640 2505.090 479.700 ;
        RECT 1718.630 479.500 2505.090 479.640 ;
        RECT 1718.630 479.440 1718.950 479.500 ;
        RECT 2504.770 479.440 2505.090 479.500 ;
      LAYER via ;
        RECT 1718.660 479.440 1718.920 479.700 ;
        RECT 2504.800 479.440 2505.060 479.700 ;
      LAYER met2 ;
        RECT 1718.790 510.340 1719.070 514.000 ;
        RECT 1718.720 510.000 1719.070 510.340 ;
        RECT 1718.720 479.730 1718.860 510.000 ;
        RECT 1718.660 479.410 1718.920 479.730 ;
        RECT 2504.800 479.410 2505.060 479.730 ;
        RECT 2504.860 17.410 2505.000 479.410 ;
        RECT 2504.860 17.270 2506.380 17.410 ;
        RECT 2506.240 2.400 2506.380 17.270 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.050 472.840 1731.370 472.900 ;
        RECT 2518.570 472.840 2518.890 472.900 ;
        RECT 1731.050 472.700 2518.890 472.840 ;
        RECT 1731.050 472.640 1731.370 472.700 ;
        RECT 2518.570 472.640 2518.890 472.700 ;
      LAYER via ;
        RECT 1731.080 472.640 1731.340 472.900 ;
        RECT 2518.600 472.640 2518.860 472.900 ;
      LAYER met2 ;
        RECT 1731.210 510.340 1731.490 514.000 ;
        RECT 1731.140 510.000 1731.490 510.340 ;
        RECT 1731.140 472.930 1731.280 510.000 ;
        RECT 1731.080 472.610 1731.340 472.930 ;
        RECT 2518.600 472.610 2518.860 472.930 ;
        RECT 2518.660 17.410 2518.800 472.610 ;
        RECT 2518.660 17.270 2524.320 17.410 ;
        RECT 2524.180 2.400 2524.320 17.270 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.310 45.120 1745.630 45.180 ;
        RECT 2542.030 45.120 2542.350 45.180 ;
        RECT 1745.310 44.980 2542.350 45.120 ;
        RECT 1745.310 44.920 1745.630 44.980 ;
        RECT 2542.030 44.920 2542.350 44.980 ;
      LAYER via ;
        RECT 1745.340 44.920 1745.600 45.180 ;
        RECT 2542.060 44.920 2542.320 45.180 ;
      LAYER met2 ;
        RECT 1743.630 510.410 1743.910 514.000 ;
        RECT 1743.630 510.270 1745.540 510.410 ;
        RECT 1743.630 510.000 1743.910 510.270 ;
        RECT 1745.400 45.210 1745.540 510.270 ;
        RECT 1745.340 44.890 1745.600 45.210 ;
        RECT 2542.060 44.890 2542.320 45.210 ;
        RECT 2542.120 2.400 2542.260 44.890 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 51.920 1759.430 51.980 ;
        RECT 2560.430 51.920 2560.750 51.980 ;
        RECT 1759.110 51.780 2560.750 51.920 ;
        RECT 1759.110 51.720 1759.430 51.780 ;
        RECT 2560.430 51.720 2560.750 51.780 ;
      LAYER via ;
        RECT 1759.140 51.720 1759.400 51.980 ;
        RECT 2560.460 51.720 2560.720 51.980 ;
      LAYER met2 ;
        RECT 1756.050 510.410 1756.330 514.000 ;
        RECT 1756.050 510.270 1759.340 510.410 ;
        RECT 1756.050 510.000 1756.330 510.270 ;
        RECT 1759.200 52.010 1759.340 510.270 ;
        RECT 1759.140 51.690 1759.400 52.010 ;
        RECT 2560.460 51.690 2560.720 52.010 ;
        RECT 2560.520 7.210 2560.660 51.690 ;
        RECT 2560.060 7.070 2560.660 7.210 ;
        RECT 2560.060 2.400 2560.200 7.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.310 496.980 1768.630 497.040 ;
        RECT 1772.450 496.980 1772.770 497.040 ;
        RECT 1768.310 496.840 1772.770 496.980 ;
        RECT 1768.310 496.780 1768.630 496.840 ;
        RECT 1772.450 496.780 1772.770 496.840 ;
        RECT 1772.450 465.700 1772.770 465.760 ;
        RECT 2573.770 465.700 2574.090 465.760 ;
        RECT 1772.450 465.560 2574.090 465.700 ;
        RECT 1772.450 465.500 1772.770 465.560 ;
        RECT 2573.770 465.500 2574.090 465.560 ;
        RECT 2573.770 62.120 2574.090 62.180 ;
        RECT 2577.910 62.120 2578.230 62.180 ;
        RECT 2573.770 61.980 2578.230 62.120 ;
        RECT 2573.770 61.920 2574.090 61.980 ;
        RECT 2577.910 61.920 2578.230 61.980 ;
      LAYER via ;
        RECT 1768.340 496.780 1768.600 497.040 ;
        RECT 1772.480 496.780 1772.740 497.040 ;
        RECT 1772.480 465.500 1772.740 465.760 ;
        RECT 2573.800 465.500 2574.060 465.760 ;
        RECT 2573.800 61.920 2574.060 62.180 ;
        RECT 2577.940 61.920 2578.200 62.180 ;
      LAYER met2 ;
        RECT 1768.470 510.340 1768.750 514.000 ;
        RECT 1768.400 510.000 1768.750 510.340 ;
        RECT 1768.400 497.070 1768.540 510.000 ;
        RECT 1768.340 496.750 1768.600 497.070 ;
        RECT 1772.480 496.750 1772.740 497.070 ;
        RECT 1772.540 465.790 1772.680 496.750 ;
        RECT 1772.480 465.470 1772.740 465.790 ;
        RECT 2573.800 465.470 2574.060 465.790 ;
        RECT 2573.860 62.210 2574.000 465.470 ;
        RECT 2573.800 61.890 2574.060 62.210 ;
        RECT 2577.940 61.890 2578.200 62.210 ;
        RECT 2578.000 2.400 2578.140 61.890 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 724.185 24.225 724.355 43.435 ;
        RECT 772.945 19.465 773.115 24.395 ;
      LAYER mcon ;
        RECT 724.185 43.265 724.355 43.435 ;
        RECT 772.945 24.225 773.115 24.395 ;
      LAYER met1 ;
        RECT 543.330 500.380 543.650 500.440 ;
        RECT 679.490 500.380 679.810 500.440 ;
        RECT 543.330 500.240 679.810 500.380 ;
        RECT 543.330 500.180 543.650 500.240 ;
        RECT 679.490 500.180 679.810 500.240 ;
        RECT 679.490 43.420 679.810 43.480 ;
        RECT 724.125 43.420 724.415 43.465 ;
        RECT 679.490 43.280 724.415 43.420 ;
        RECT 679.490 43.220 679.810 43.280 ;
        RECT 724.125 43.235 724.415 43.280 ;
        RECT 724.125 24.380 724.415 24.425 ;
        RECT 772.885 24.380 773.175 24.425 ;
        RECT 724.125 24.240 773.175 24.380 ;
        RECT 724.125 24.195 724.415 24.240 ;
        RECT 772.885 24.195 773.175 24.240 ;
        RECT 772.885 19.620 773.175 19.665 ;
        RECT 811.510 19.620 811.830 19.680 ;
        RECT 772.885 19.480 811.830 19.620 ;
        RECT 772.885 19.435 773.175 19.480 ;
        RECT 811.510 19.420 811.830 19.480 ;
      LAYER via ;
        RECT 543.360 500.180 543.620 500.440 ;
        RECT 679.520 500.180 679.780 500.440 ;
        RECT 679.520 43.220 679.780 43.480 ;
        RECT 811.540 19.420 811.800 19.680 ;
      LAYER met2 ;
        RECT 543.490 510.340 543.770 514.000 ;
        RECT 543.420 510.000 543.770 510.340 ;
        RECT 543.420 500.470 543.560 510.000 ;
        RECT 543.360 500.150 543.620 500.470 ;
        RECT 679.520 500.150 679.780 500.470 ;
        RECT 679.580 43.510 679.720 500.150 ;
        RECT 679.520 43.190 679.780 43.510 ;
        RECT 811.540 19.390 811.800 19.710 ;
        RECT 811.600 2.400 811.740 19.390 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2594.545 379.525 2594.715 427.635 ;
        RECT 2594.545 282.965 2594.715 331.075 ;
        RECT 2594.545 186.405 2594.715 234.515 ;
        RECT 2594.545 89.845 2594.715 137.955 ;
        RECT 2595.465 2.805 2595.635 48.195 ;
      LAYER mcon ;
        RECT 2594.545 427.465 2594.715 427.635 ;
        RECT 2594.545 330.905 2594.715 331.075 ;
        RECT 2594.545 234.345 2594.715 234.515 ;
        RECT 2594.545 137.785 2594.715 137.955 ;
        RECT 2595.465 48.025 2595.635 48.195 ;
      LAYER met1 ;
        RECT 1780.270 496.980 1780.590 497.040 ;
        RECT 1786.250 496.980 1786.570 497.040 ;
        RECT 1780.270 496.840 1786.570 496.980 ;
        RECT 1780.270 496.780 1780.590 496.840 ;
        RECT 1786.250 496.780 1786.570 496.840 ;
        RECT 1786.250 458.900 1786.570 458.960 ;
        RECT 2594.470 458.900 2594.790 458.960 ;
        RECT 1786.250 458.760 2594.790 458.900 ;
        RECT 1786.250 458.700 1786.570 458.760 ;
        RECT 2594.470 458.700 2594.790 458.760 ;
        RECT 2594.470 427.620 2594.790 427.680 ;
        RECT 2594.275 427.480 2594.790 427.620 ;
        RECT 2594.470 427.420 2594.790 427.480 ;
        RECT 2594.470 379.680 2594.790 379.740 ;
        RECT 2594.275 379.540 2594.790 379.680 ;
        RECT 2594.470 379.480 2594.790 379.540 ;
        RECT 2594.470 331.060 2594.790 331.120 ;
        RECT 2594.275 330.920 2594.790 331.060 ;
        RECT 2594.470 330.860 2594.790 330.920 ;
        RECT 2594.470 283.120 2594.790 283.180 ;
        RECT 2594.275 282.980 2594.790 283.120 ;
        RECT 2594.470 282.920 2594.790 282.980 ;
        RECT 2594.470 234.500 2594.790 234.560 ;
        RECT 2594.275 234.360 2594.790 234.500 ;
        RECT 2594.470 234.300 2594.790 234.360 ;
        RECT 2594.470 186.560 2594.790 186.620 ;
        RECT 2594.275 186.420 2594.790 186.560 ;
        RECT 2594.470 186.360 2594.790 186.420 ;
        RECT 2594.470 137.940 2594.790 138.000 ;
        RECT 2594.275 137.800 2594.790 137.940 ;
        RECT 2594.470 137.740 2594.790 137.800 ;
        RECT 2594.470 90.000 2594.790 90.060 ;
        RECT 2594.275 89.860 2594.790 90.000 ;
        RECT 2594.470 89.800 2594.790 89.860 ;
        RECT 2594.470 62.260 2594.790 62.520 ;
        RECT 2594.560 61.780 2594.700 62.260 ;
        RECT 2595.390 61.780 2595.710 61.840 ;
        RECT 2594.560 61.640 2595.710 61.780 ;
        RECT 2595.390 61.580 2595.710 61.640 ;
        RECT 2595.390 48.180 2595.710 48.240 ;
        RECT 2595.195 48.040 2595.710 48.180 ;
        RECT 2595.390 47.980 2595.710 48.040 ;
        RECT 2595.390 2.960 2595.710 3.020 ;
        RECT 2595.195 2.820 2595.710 2.960 ;
        RECT 2595.390 2.760 2595.710 2.820 ;
      LAYER via ;
        RECT 1780.300 496.780 1780.560 497.040 ;
        RECT 1786.280 496.780 1786.540 497.040 ;
        RECT 1786.280 458.700 1786.540 458.960 ;
        RECT 2594.500 458.700 2594.760 458.960 ;
        RECT 2594.500 427.420 2594.760 427.680 ;
        RECT 2594.500 379.480 2594.760 379.740 ;
        RECT 2594.500 330.860 2594.760 331.120 ;
        RECT 2594.500 282.920 2594.760 283.180 ;
        RECT 2594.500 234.300 2594.760 234.560 ;
        RECT 2594.500 186.360 2594.760 186.620 ;
        RECT 2594.500 137.740 2594.760 138.000 ;
        RECT 2594.500 89.800 2594.760 90.060 ;
        RECT 2594.500 62.260 2594.760 62.520 ;
        RECT 2595.420 61.580 2595.680 61.840 ;
        RECT 2595.420 47.980 2595.680 48.240 ;
        RECT 2595.420 2.760 2595.680 3.020 ;
      LAYER met2 ;
        RECT 1780.430 510.340 1780.710 514.000 ;
        RECT 1780.360 510.000 1780.710 510.340 ;
        RECT 1780.360 497.070 1780.500 510.000 ;
        RECT 1780.300 496.750 1780.560 497.070 ;
        RECT 1786.280 496.750 1786.540 497.070 ;
        RECT 1786.340 458.990 1786.480 496.750 ;
        RECT 1786.280 458.670 1786.540 458.990 ;
        RECT 2594.500 458.670 2594.760 458.990 ;
        RECT 2594.560 427.710 2594.700 458.670 ;
        RECT 2594.500 427.390 2594.760 427.710 ;
        RECT 2594.500 379.450 2594.760 379.770 ;
        RECT 2594.560 331.150 2594.700 379.450 ;
        RECT 2594.500 330.830 2594.760 331.150 ;
        RECT 2594.500 282.890 2594.760 283.210 ;
        RECT 2594.560 234.590 2594.700 282.890 ;
        RECT 2594.500 234.270 2594.760 234.590 ;
        RECT 2594.500 186.330 2594.760 186.650 ;
        RECT 2594.560 138.030 2594.700 186.330 ;
        RECT 2594.500 137.710 2594.760 138.030 ;
        RECT 2594.500 89.770 2594.760 90.090 ;
        RECT 2594.560 62.550 2594.700 89.770 ;
        RECT 2594.500 62.230 2594.760 62.550 ;
        RECT 2595.420 61.550 2595.680 61.870 ;
        RECT 2595.480 48.270 2595.620 61.550 ;
        RECT 2595.420 47.950 2595.680 48.270 ;
        RECT 2595.420 2.730 2595.680 3.050 ;
        RECT 2595.480 2.400 2595.620 2.730 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1792.690 451.760 1793.010 451.820 ;
        RECT 2608.270 451.760 2608.590 451.820 ;
        RECT 1792.690 451.620 2608.590 451.760 ;
        RECT 1792.690 451.560 1793.010 451.620 ;
        RECT 2608.270 451.560 2608.590 451.620 ;
        RECT 2608.270 62.120 2608.590 62.180 ;
        RECT 2613.330 62.120 2613.650 62.180 ;
        RECT 2608.270 61.980 2613.650 62.120 ;
        RECT 2608.270 61.920 2608.590 61.980 ;
        RECT 2613.330 61.920 2613.650 61.980 ;
      LAYER via ;
        RECT 1792.720 451.560 1792.980 451.820 ;
        RECT 2608.300 451.560 2608.560 451.820 ;
        RECT 2608.300 61.920 2608.560 62.180 ;
        RECT 2613.360 61.920 2613.620 62.180 ;
      LAYER met2 ;
        RECT 1792.850 510.340 1793.130 514.000 ;
        RECT 1792.780 510.000 1793.130 510.340 ;
        RECT 1792.780 451.850 1792.920 510.000 ;
        RECT 1792.720 451.530 1792.980 451.850 ;
        RECT 2608.300 451.530 2608.560 451.850 ;
        RECT 2608.360 62.210 2608.500 451.530 ;
        RECT 2608.300 61.890 2608.560 62.210 ;
        RECT 2613.360 61.890 2613.620 62.210 ;
        RECT 2613.420 2.400 2613.560 61.890 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1805.110 497.320 1805.430 497.380 ;
        RECT 1817.990 497.320 1818.310 497.380 ;
        RECT 1805.110 497.180 1818.310 497.320 ;
        RECT 1805.110 497.120 1805.430 497.180 ;
        RECT 1817.990 497.120 1818.310 497.180 ;
        RECT 1817.990 59.060 1818.310 59.120 ;
        RECT 2631.270 59.060 2631.590 59.120 ;
        RECT 1817.990 58.920 2631.590 59.060 ;
        RECT 1817.990 58.860 1818.310 58.920 ;
        RECT 2631.270 58.860 2631.590 58.920 ;
      LAYER via ;
        RECT 1805.140 497.120 1805.400 497.380 ;
        RECT 1818.020 497.120 1818.280 497.380 ;
        RECT 1818.020 58.860 1818.280 59.120 ;
        RECT 2631.300 58.860 2631.560 59.120 ;
      LAYER met2 ;
        RECT 1805.270 510.340 1805.550 514.000 ;
        RECT 1805.200 510.000 1805.550 510.340 ;
        RECT 1805.200 497.410 1805.340 510.000 ;
        RECT 1805.140 497.090 1805.400 497.410 ;
        RECT 1818.020 497.090 1818.280 497.410 ;
        RECT 1818.080 59.150 1818.220 497.090 ;
        RECT 1818.020 58.830 1818.280 59.150 ;
        RECT 2631.300 58.830 2631.560 59.150 ;
        RECT 2631.360 2.400 2631.500 58.830 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 444.960 1821.530 445.020 ;
        RECT 2642.770 444.960 2643.090 445.020 ;
        RECT 1821.210 444.820 2643.090 444.960 ;
        RECT 1821.210 444.760 1821.530 444.820 ;
        RECT 2642.770 444.760 2643.090 444.820 ;
        RECT 2642.770 37.980 2643.090 38.040 ;
        RECT 2649.210 37.980 2649.530 38.040 ;
        RECT 2642.770 37.840 2649.530 37.980 ;
        RECT 2642.770 37.780 2643.090 37.840 ;
        RECT 2649.210 37.780 2649.530 37.840 ;
      LAYER via ;
        RECT 1821.240 444.760 1821.500 445.020 ;
        RECT 2642.800 444.760 2643.060 445.020 ;
        RECT 2642.800 37.780 2643.060 38.040 ;
        RECT 2649.240 37.780 2649.500 38.040 ;
      LAYER met2 ;
        RECT 1817.690 510.410 1817.970 514.000 ;
        RECT 1817.690 510.270 1821.440 510.410 ;
        RECT 1817.690 510.000 1817.970 510.270 ;
        RECT 1821.300 445.050 1821.440 510.270 ;
        RECT 1821.240 444.730 1821.500 445.050 ;
        RECT 2642.800 444.730 2643.060 445.050 ;
        RECT 2642.860 38.070 2643.000 444.730 ;
        RECT 2642.800 37.750 2643.060 38.070 ;
        RECT 2649.240 37.750 2649.500 38.070 ;
        RECT 2649.300 2.400 2649.440 37.750 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2663.545 379.525 2663.715 427.635 ;
        RECT 2663.545 282.965 2663.715 331.075 ;
        RECT 2663.545 186.405 2663.715 234.515 ;
        RECT 2663.545 48.365 2663.715 137.955 ;
      LAYER mcon ;
        RECT 2663.545 427.465 2663.715 427.635 ;
        RECT 2663.545 330.905 2663.715 331.075 ;
        RECT 2663.545 234.345 2663.715 234.515 ;
        RECT 2663.545 137.785 2663.715 137.955 ;
      LAYER met1 ;
        RECT 1829.950 496.980 1830.270 497.040 ;
        RECT 1834.550 496.980 1834.870 497.040 ;
        RECT 1829.950 496.840 1834.870 496.980 ;
        RECT 1829.950 496.780 1830.270 496.840 ;
        RECT 1834.550 496.780 1834.870 496.840 ;
        RECT 1834.550 431.360 1834.870 431.420 ;
        RECT 2663.470 431.360 2663.790 431.420 ;
        RECT 1834.550 431.220 2663.790 431.360 ;
        RECT 1834.550 431.160 1834.870 431.220 ;
        RECT 2663.470 431.160 2663.790 431.220 ;
        RECT 2663.470 427.620 2663.790 427.680 ;
        RECT 2663.275 427.480 2663.790 427.620 ;
        RECT 2663.470 427.420 2663.790 427.480 ;
        RECT 2663.470 379.680 2663.790 379.740 ;
        RECT 2663.275 379.540 2663.790 379.680 ;
        RECT 2663.470 379.480 2663.790 379.540 ;
        RECT 2663.470 331.060 2663.790 331.120 ;
        RECT 2663.275 330.920 2663.790 331.060 ;
        RECT 2663.470 330.860 2663.790 330.920 ;
        RECT 2663.470 283.120 2663.790 283.180 ;
        RECT 2663.275 282.980 2663.790 283.120 ;
        RECT 2663.470 282.920 2663.790 282.980 ;
        RECT 2663.470 234.500 2663.790 234.560 ;
        RECT 2663.275 234.360 2663.790 234.500 ;
        RECT 2663.470 234.300 2663.790 234.360 ;
        RECT 2663.470 186.560 2663.790 186.620 ;
        RECT 2663.275 186.420 2663.790 186.560 ;
        RECT 2663.470 186.360 2663.790 186.420 ;
        RECT 2663.470 137.940 2663.790 138.000 ;
        RECT 2663.275 137.800 2663.790 137.940 ;
        RECT 2663.470 137.740 2663.790 137.800 ;
        RECT 2663.485 48.520 2663.775 48.565 ;
        RECT 2667.150 48.520 2667.470 48.580 ;
        RECT 2663.485 48.380 2667.470 48.520 ;
        RECT 2663.485 48.335 2663.775 48.380 ;
        RECT 2667.150 48.320 2667.470 48.380 ;
      LAYER via ;
        RECT 1829.980 496.780 1830.240 497.040 ;
        RECT 1834.580 496.780 1834.840 497.040 ;
        RECT 1834.580 431.160 1834.840 431.420 ;
        RECT 2663.500 431.160 2663.760 431.420 ;
        RECT 2663.500 427.420 2663.760 427.680 ;
        RECT 2663.500 379.480 2663.760 379.740 ;
        RECT 2663.500 330.860 2663.760 331.120 ;
        RECT 2663.500 282.920 2663.760 283.180 ;
        RECT 2663.500 234.300 2663.760 234.560 ;
        RECT 2663.500 186.360 2663.760 186.620 ;
        RECT 2663.500 137.740 2663.760 138.000 ;
        RECT 2667.180 48.320 2667.440 48.580 ;
      LAYER met2 ;
        RECT 1830.110 510.340 1830.390 514.000 ;
        RECT 1830.040 510.000 1830.390 510.340 ;
        RECT 1830.040 497.070 1830.180 510.000 ;
        RECT 1829.980 496.750 1830.240 497.070 ;
        RECT 1834.580 496.750 1834.840 497.070 ;
        RECT 1834.640 431.450 1834.780 496.750 ;
        RECT 1834.580 431.130 1834.840 431.450 ;
        RECT 2663.500 431.130 2663.760 431.450 ;
        RECT 2663.560 427.710 2663.700 431.130 ;
        RECT 2663.500 427.390 2663.760 427.710 ;
        RECT 2663.500 379.450 2663.760 379.770 ;
        RECT 2663.560 331.150 2663.700 379.450 ;
        RECT 2663.500 330.830 2663.760 331.150 ;
        RECT 2663.500 282.890 2663.760 283.210 ;
        RECT 2663.560 234.590 2663.700 282.890 ;
        RECT 2663.500 234.270 2663.760 234.590 ;
        RECT 2663.500 186.330 2663.760 186.650 ;
        RECT 2663.560 138.030 2663.700 186.330 ;
        RECT 2663.500 137.710 2663.760 138.030 ;
        RECT 2667.180 48.290 2667.440 48.610 ;
        RECT 2667.240 2.400 2667.380 48.290 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1842.370 496.980 1842.690 497.040 ;
        RECT 1848.350 496.980 1848.670 497.040 ;
        RECT 1842.370 496.840 1848.670 496.980 ;
        RECT 1842.370 496.780 1842.690 496.840 ;
        RECT 1848.350 496.780 1848.670 496.840 ;
        RECT 1848.350 424.220 1848.670 424.280 ;
        RECT 2684.170 424.220 2684.490 424.280 ;
        RECT 1848.350 424.080 2684.490 424.220 ;
        RECT 1848.350 424.020 1848.670 424.080 ;
        RECT 2684.170 424.020 2684.490 424.080 ;
      LAYER via ;
        RECT 1842.400 496.780 1842.660 497.040 ;
        RECT 1848.380 496.780 1848.640 497.040 ;
        RECT 1848.380 424.020 1848.640 424.280 ;
        RECT 2684.200 424.020 2684.460 424.280 ;
      LAYER met2 ;
        RECT 1842.530 510.340 1842.810 514.000 ;
        RECT 1842.460 510.000 1842.810 510.340 ;
        RECT 1842.460 497.070 1842.600 510.000 ;
        RECT 1842.400 496.750 1842.660 497.070 ;
        RECT 1848.380 496.750 1848.640 497.070 ;
        RECT 1848.440 424.310 1848.580 496.750 ;
        RECT 1848.380 423.990 1848.640 424.310 ;
        RECT 2684.200 423.990 2684.460 424.310 ;
        RECT 2684.260 17.410 2684.400 423.990 ;
        RECT 2684.260 17.270 2684.860 17.410 ;
        RECT 2684.720 2.400 2684.860 17.270 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1854.405 496.485 1854.575 510.595 ;
      LAYER mcon ;
        RECT 1854.405 510.425 1854.575 510.595 ;
      LAYER met1 ;
        RECT 1854.330 510.580 1854.650 510.640 ;
        RECT 1854.135 510.440 1854.650 510.580 ;
        RECT 1854.330 510.380 1854.650 510.440 ;
        RECT 1854.330 496.640 1854.650 496.700 ;
        RECT 1854.135 496.500 1854.650 496.640 ;
        RECT 1854.330 496.440 1854.650 496.500 ;
        RECT 1853.410 417.420 1853.730 417.480 ;
        RECT 2697.970 417.420 2698.290 417.480 ;
        RECT 1853.410 417.280 2698.290 417.420 ;
        RECT 1853.410 417.220 1853.730 417.280 ;
        RECT 2697.970 417.220 2698.290 417.280 ;
      LAYER via ;
        RECT 1854.360 510.380 1854.620 510.640 ;
        RECT 1854.360 496.440 1854.620 496.700 ;
        RECT 1853.440 417.220 1853.700 417.480 ;
        RECT 2698.000 417.220 2698.260 417.480 ;
      LAYER met2 ;
        RECT 1854.950 511.090 1855.230 514.000 ;
        RECT 1854.420 510.950 1855.230 511.090 ;
        RECT 1854.420 510.670 1854.560 510.950 ;
        RECT 1854.360 510.350 1854.620 510.670 ;
        RECT 1854.950 510.000 1855.230 510.950 ;
        RECT 1854.360 496.410 1854.620 496.730 ;
        RECT 1854.420 435.045 1854.560 496.410 ;
        RECT 1853.430 434.675 1853.710 435.045 ;
        RECT 1854.350 434.675 1854.630 435.045 ;
        RECT 1853.500 417.510 1853.640 434.675 ;
        RECT 1853.440 417.190 1853.700 417.510 ;
        RECT 2698.000 417.190 2698.260 417.510 ;
        RECT 2698.060 16.730 2698.200 417.190 ;
        RECT 2698.060 16.590 2702.800 16.730 ;
        RECT 2702.660 2.400 2702.800 16.590 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
      LAYER via2 ;
        RECT 1853.430 434.720 1853.710 435.000 ;
        RECT 1854.350 434.720 1854.630 435.000 ;
      LAYER met3 ;
        RECT 1853.405 435.010 1853.735 435.025 ;
        RECT 1854.325 435.010 1854.655 435.025 ;
        RECT 1853.405 434.710 1854.655 435.010 ;
        RECT 1853.405 434.695 1853.735 434.710 ;
        RECT 1854.325 434.695 1854.655 434.710 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.510 65.520 1869.830 65.580 ;
        RECT 2720.510 65.520 2720.830 65.580 ;
        RECT 1869.510 65.380 2720.830 65.520 ;
        RECT 1869.510 65.320 1869.830 65.380 ;
        RECT 2720.510 65.320 2720.830 65.380 ;
      LAYER via ;
        RECT 1869.540 65.320 1869.800 65.580 ;
        RECT 2720.540 65.320 2720.800 65.580 ;
      LAYER met2 ;
        RECT 1867.370 510.410 1867.650 514.000 ;
        RECT 1867.370 510.270 1869.740 510.410 ;
        RECT 1867.370 510.000 1867.650 510.270 ;
        RECT 1869.600 65.610 1869.740 510.270 ;
        RECT 1869.540 65.290 1869.800 65.610 ;
        RECT 2720.540 65.290 2720.800 65.610 ;
        RECT 2720.600 2.400 2720.740 65.290 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1879.630 503.440 1879.950 503.500 ;
        RECT 1883.310 503.440 1883.630 503.500 ;
        RECT 1879.630 503.300 1883.630 503.440 ;
        RECT 1879.630 503.240 1879.950 503.300 ;
        RECT 1883.310 503.240 1883.630 503.300 ;
        RECT 1883.310 86.260 1883.630 86.320 ;
        RECT 2732.470 86.260 2732.790 86.320 ;
        RECT 1883.310 86.120 2732.790 86.260 ;
        RECT 1883.310 86.060 1883.630 86.120 ;
        RECT 2732.470 86.060 2732.790 86.120 ;
        RECT 2732.470 37.980 2732.790 38.040 ;
        RECT 2738.450 37.980 2738.770 38.040 ;
        RECT 2732.470 37.840 2738.770 37.980 ;
        RECT 2732.470 37.780 2732.790 37.840 ;
        RECT 2738.450 37.780 2738.770 37.840 ;
      LAYER via ;
        RECT 1879.660 503.240 1879.920 503.500 ;
        RECT 1883.340 503.240 1883.600 503.500 ;
        RECT 1883.340 86.060 1883.600 86.320 ;
        RECT 2732.500 86.060 2732.760 86.320 ;
        RECT 2732.500 37.780 2732.760 38.040 ;
        RECT 2738.480 37.780 2738.740 38.040 ;
      LAYER met2 ;
        RECT 1879.790 510.340 1880.070 514.000 ;
        RECT 1879.720 510.000 1880.070 510.340 ;
        RECT 1879.720 503.530 1879.860 510.000 ;
        RECT 1879.660 503.210 1879.920 503.530 ;
        RECT 1883.340 503.210 1883.600 503.530 ;
        RECT 1883.400 86.350 1883.540 503.210 ;
        RECT 1883.340 86.030 1883.600 86.350 ;
        RECT 2732.500 86.030 2732.760 86.350 ;
        RECT 2732.560 38.070 2732.700 86.030 ;
        RECT 2732.500 37.750 2732.760 38.070 ;
        RECT 2738.480 37.750 2738.740 38.070 ;
        RECT 2738.540 2.400 2738.680 37.750 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2753.245 61.625 2753.415 96.475 ;
      LAYER mcon ;
        RECT 2753.245 96.305 2753.415 96.475 ;
      LAYER met1 ;
        RECT 1891.590 497.320 1891.910 497.380 ;
        RECT 1907.690 497.320 1908.010 497.380 ;
        RECT 1891.590 497.180 1908.010 497.320 ;
        RECT 1891.590 497.120 1891.910 497.180 ;
        RECT 1907.690 497.120 1908.010 497.180 ;
        RECT 1907.690 410.620 1908.010 410.680 ;
        RECT 2753.170 410.620 2753.490 410.680 ;
        RECT 1907.690 410.480 2753.490 410.620 ;
        RECT 1907.690 410.420 1908.010 410.480 ;
        RECT 2753.170 410.420 2753.490 410.480 ;
        RECT 2753.170 338.200 2753.490 338.260 ;
        RECT 2754.550 338.200 2754.870 338.260 ;
        RECT 2753.170 338.060 2754.870 338.200 ;
        RECT 2753.170 338.000 2753.490 338.060 ;
        RECT 2754.550 338.000 2754.870 338.060 ;
        RECT 2753.170 96.460 2753.490 96.520 ;
        RECT 2753.170 96.320 2753.685 96.460 ;
        RECT 2753.170 96.260 2753.490 96.320 ;
        RECT 2753.185 61.780 2753.475 61.825 ;
        RECT 2755.930 61.780 2756.250 61.840 ;
        RECT 2753.185 61.640 2756.250 61.780 ;
        RECT 2753.185 61.595 2753.475 61.640 ;
        RECT 2755.930 61.580 2756.250 61.640 ;
      LAYER via ;
        RECT 1891.620 497.120 1891.880 497.380 ;
        RECT 1907.720 497.120 1907.980 497.380 ;
        RECT 1907.720 410.420 1907.980 410.680 ;
        RECT 2753.200 410.420 2753.460 410.680 ;
        RECT 2753.200 338.000 2753.460 338.260 ;
        RECT 2754.580 338.000 2754.840 338.260 ;
        RECT 2753.200 96.260 2753.460 96.520 ;
        RECT 2755.960 61.580 2756.220 61.840 ;
      LAYER met2 ;
        RECT 1891.750 510.340 1892.030 514.000 ;
        RECT 1891.680 510.000 1892.030 510.340 ;
        RECT 1891.680 497.410 1891.820 510.000 ;
        RECT 1891.620 497.090 1891.880 497.410 ;
        RECT 1907.720 497.090 1907.980 497.410 ;
        RECT 1907.780 410.710 1907.920 497.090 ;
        RECT 1907.720 410.390 1907.980 410.710 ;
        RECT 2753.200 410.390 2753.460 410.710 ;
        RECT 2753.260 386.085 2753.400 410.390 ;
        RECT 2753.190 385.715 2753.470 386.085 ;
        RECT 2754.570 385.715 2754.850 386.085 ;
        RECT 2754.640 338.290 2754.780 385.715 ;
        RECT 2753.200 337.970 2753.460 338.290 ;
        RECT 2754.580 337.970 2754.840 338.290 ;
        RECT 2753.260 290.885 2753.400 337.970 ;
        RECT 2753.190 290.515 2753.470 290.885 ;
        RECT 2753.190 289.835 2753.470 290.205 ;
        RECT 2753.260 96.550 2753.400 289.835 ;
        RECT 2753.200 96.230 2753.460 96.550 ;
        RECT 2755.960 61.550 2756.220 61.870 ;
        RECT 2756.020 2.400 2756.160 61.550 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
      LAYER via2 ;
        RECT 2753.190 385.760 2753.470 386.040 ;
        RECT 2754.570 385.760 2754.850 386.040 ;
        RECT 2753.190 290.560 2753.470 290.840 ;
        RECT 2753.190 289.880 2753.470 290.160 ;
      LAYER met3 ;
        RECT 2753.165 386.050 2753.495 386.065 ;
        RECT 2754.545 386.050 2754.875 386.065 ;
        RECT 2753.165 385.750 2754.875 386.050 ;
        RECT 2753.165 385.735 2753.495 385.750 ;
        RECT 2754.545 385.735 2754.875 385.750 ;
        RECT 2753.165 290.850 2753.495 290.865 ;
        RECT 2752.950 290.535 2753.495 290.850 ;
        RECT 2752.950 290.185 2753.250 290.535 ;
        RECT 2752.950 289.870 2753.495 290.185 ;
        RECT 2753.165 289.855 2753.495 289.870 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.510 30.840 558.830 30.900 ;
        RECT 829.450 30.840 829.770 30.900 ;
        RECT 558.510 30.700 829.770 30.840 ;
        RECT 558.510 30.640 558.830 30.700 ;
        RECT 829.450 30.640 829.770 30.700 ;
      LAYER via ;
        RECT 558.540 30.640 558.800 30.900 ;
        RECT 829.480 30.640 829.740 30.900 ;
      LAYER met2 ;
        RECT 555.910 510.410 556.190 514.000 ;
        RECT 555.910 510.270 558.740 510.410 ;
        RECT 555.910 510.000 556.190 510.270 ;
        RECT 558.600 30.930 558.740 510.270 ;
        RECT 558.540 30.610 558.800 30.930 ;
        RECT 829.480 30.610 829.740 30.930 ;
        RECT 829.540 2.400 829.680 30.610 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 93.060 1904.330 93.120 ;
        RECT 2774.330 93.060 2774.650 93.120 ;
        RECT 1904.010 92.920 2774.650 93.060 ;
        RECT 1904.010 92.860 1904.330 92.920 ;
        RECT 2774.330 92.860 2774.650 92.920 ;
      LAYER via ;
        RECT 1904.040 92.860 1904.300 93.120 ;
        RECT 2774.360 92.860 2774.620 93.120 ;
      LAYER met2 ;
        RECT 1904.170 510.340 1904.450 514.000 ;
        RECT 1904.100 510.000 1904.450 510.340 ;
        RECT 1904.100 93.150 1904.240 510.000 ;
        RECT 1904.040 92.830 1904.300 93.150 ;
        RECT 2774.360 92.830 2774.620 93.150 ;
        RECT 2774.420 37.130 2774.560 92.830 ;
        RECT 2773.960 36.990 2774.560 37.130 ;
        RECT 2773.960 2.400 2774.100 36.990 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1916.430 497.320 1916.750 497.380 ;
        RECT 1928.390 497.320 1928.710 497.380 ;
        RECT 1916.430 497.180 1928.710 497.320 ;
        RECT 1916.430 497.120 1916.750 497.180 ;
        RECT 1928.390 497.120 1928.710 497.180 ;
        RECT 1928.390 403.480 1928.710 403.540 ;
        RECT 2787.670 403.480 2787.990 403.540 ;
        RECT 1928.390 403.340 2787.990 403.480 ;
        RECT 1928.390 403.280 1928.710 403.340 ;
        RECT 2787.670 403.280 2787.990 403.340 ;
        RECT 2787.670 62.120 2787.990 62.180 ;
        RECT 2791.810 62.120 2792.130 62.180 ;
        RECT 2787.670 61.980 2792.130 62.120 ;
        RECT 2787.670 61.920 2787.990 61.980 ;
        RECT 2791.810 61.920 2792.130 61.980 ;
      LAYER via ;
        RECT 1916.460 497.120 1916.720 497.380 ;
        RECT 1928.420 497.120 1928.680 497.380 ;
        RECT 1928.420 403.280 1928.680 403.540 ;
        RECT 2787.700 403.280 2787.960 403.540 ;
        RECT 2787.700 61.920 2787.960 62.180 ;
        RECT 2791.840 61.920 2792.100 62.180 ;
      LAYER met2 ;
        RECT 1916.590 510.340 1916.870 514.000 ;
        RECT 1916.520 510.000 1916.870 510.340 ;
        RECT 1916.520 497.410 1916.660 510.000 ;
        RECT 1916.460 497.090 1916.720 497.410 ;
        RECT 1928.420 497.090 1928.680 497.410 ;
        RECT 1928.480 403.570 1928.620 497.090 ;
        RECT 1928.420 403.250 1928.680 403.570 ;
        RECT 2787.700 403.250 2787.960 403.570 ;
        RECT 2787.760 62.210 2787.900 403.250 ;
        RECT 2787.700 61.890 2787.960 62.210 ;
        RECT 2791.840 61.890 2792.100 62.210 ;
        RECT 2791.900 2.400 2792.040 61.890 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.610 72.320 1931.930 72.380 ;
        RECT 2809.750 72.320 2810.070 72.380 ;
        RECT 1931.610 72.180 2810.070 72.320 ;
        RECT 1931.610 72.120 1931.930 72.180 ;
        RECT 2809.750 72.120 2810.070 72.180 ;
      LAYER via ;
        RECT 1931.640 72.120 1931.900 72.380 ;
        RECT 2809.780 72.120 2810.040 72.380 ;
      LAYER met2 ;
        RECT 1929.010 510.410 1929.290 514.000 ;
        RECT 1929.010 510.270 1931.840 510.410 ;
        RECT 1929.010 510.000 1929.290 510.270 ;
        RECT 1931.700 72.410 1931.840 510.270 ;
        RECT 1931.640 72.090 1931.900 72.410 ;
        RECT 2809.780 72.090 2810.040 72.410 ;
        RECT 2809.840 2.400 2809.980 72.090 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1941.270 496.980 1941.590 497.040 ;
        RECT 1944.950 496.980 1945.270 497.040 ;
        RECT 1941.270 496.840 1945.270 496.980 ;
        RECT 1941.270 496.780 1941.590 496.840 ;
        RECT 1944.950 496.780 1945.270 496.840 ;
        RECT 1944.950 396.680 1945.270 396.740 ;
        RECT 2822.170 396.680 2822.490 396.740 ;
        RECT 1944.950 396.540 2822.490 396.680 ;
        RECT 1944.950 396.480 1945.270 396.540 ;
        RECT 2822.170 396.480 2822.490 396.540 ;
        RECT 2822.170 62.120 2822.490 62.180 ;
        RECT 2827.690 62.120 2828.010 62.180 ;
        RECT 2822.170 61.980 2828.010 62.120 ;
        RECT 2822.170 61.920 2822.490 61.980 ;
        RECT 2827.690 61.920 2828.010 61.980 ;
      LAYER via ;
        RECT 1941.300 496.780 1941.560 497.040 ;
        RECT 1944.980 496.780 1945.240 497.040 ;
        RECT 1944.980 396.480 1945.240 396.740 ;
        RECT 2822.200 396.480 2822.460 396.740 ;
        RECT 2822.200 61.920 2822.460 62.180 ;
        RECT 2827.720 61.920 2827.980 62.180 ;
      LAYER met2 ;
        RECT 1941.430 510.340 1941.710 514.000 ;
        RECT 1941.360 510.000 1941.710 510.340 ;
        RECT 1941.360 497.070 1941.500 510.000 ;
        RECT 1941.300 496.750 1941.560 497.070 ;
        RECT 1944.980 496.750 1945.240 497.070 ;
        RECT 1945.040 396.770 1945.180 496.750 ;
        RECT 1944.980 396.450 1945.240 396.770 ;
        RECT 2822.200 396.450 2822.460 396.770 ;
        RECT 2822.260 62.210 2822.400 396.450 ;
        RECT 2822.200 61.890 2822.460 62.210 ;
        RECT 2827.720 61.890 2827.980 62.210 ;
        RECT 2827.780 2.400 2827.920 61.890 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.690 496.980 1954.010 497.040 ;
        RECT 1958.750 496.980 1959.070 497.040 ;
        RECT 1953.690 496.840 1959.070 496.980 ;
        RECT 1953.690 496.780 1954.010 496.840 ;
        RECT 1958.750 496.780 1959.070 496.840 ;
        RECT 1958.750 389.880 1959.070 389.940 ;
        RECT 2842.870 389.880 2843.190 389.940 ;
        RECT 1958.750 389.740 2843.190 389.880 ;
        RECT 1958.750 389.680 1959.070 389.740 ;
        RECT 2842.870 389.680 2843.190 389.740 ;
        RECT 2842.870 62.260 2843.190 62.520 ;
        RECT 2842.960 62.120 2843.100 62.260 ;
        RECT 2845.170 62.120 2845.490 62.180 ;
        RECT 2842.960 61.980 2845.490 62.120 ;
        RECT 2845.170 61.920 2845.490 61.980 ;
      LAYER via ;
        RECT 1953.720 496.780 1953.980 497.040 ;
        RECT 1958.780 496.780 1959.040 497.040 ;
        RECT 1958.780 389.680 1959.040 389.940 ;
        RECT 2842.900 389.680 2843.160 389.940 ;
        RECT 2842.900 62.260 2843.160 62.520 ;
        RECT 2845.200 61.920 2845.460 62.180 ;
      LAYER met2 ;
        RECT 1953.850 510.340 1954.130 514.000 ;
        RECT 1953.780 510.000 1954.130 510.340 ;
        RECT 1953.780 497.070 1953.920 510.000 ;
        RECT 1953.720 496.750 1953.980 497.070 ;
        RECT 1958.780 496.750 1959.040 497.070 ;
        RECT 1958.840 389.970 1958.980 496.750 ;
        RECT 1958.780 389.650 1959.040 389.970 ;
        RECT 2842.900 389.650 2843.160 389.970 ;
        RECT 2842.960 242.605 2843.100 389.650 ;
        RECT 2842.890 242.235 2843.170 242.605 ;
        RECT 2842.890 241.555 2843.170 241.925 ;
        RECT 2842.960 62.550 2843.100 241.555 ;
        RECT 2842.900 62.230 2843.160 62.550 ;
        RECT 2845.200 61.890 2845.460 62.210 ;
        RECT 2845.260 2.400 2845.400 61.890 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 2842.890 242.280 2843.170 242.560 ;
        RECT 2842.890 241.600 2843.170 241.880 ;
      LAYER met3 ;
        RECT 2842.865 242.570 2843.195 242.585 ;
        RECT 2842.190 242.270 2843.195 242.570 ;
        RECT 2842.190 241.890 2842.490 242.270 ;
        RECT 2842.865 242.255 2843.195 242.270 ;
        RECT 2842.865 241.890 2843.195 241.905 ;
        RECT 2842.190 241.590 2843.195 241.890 ;
        RECT 2842.865 241.575 2843.195 241.590 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 375.940 1966.430 376.000 ;
        RECT 2856.670 375.940 2856.990 376.000 ;
        RECT 1966.110 375.800 2856.990 375.940 ;
        RECT 1966.110 375.740 1966.430 375.800 ;
        RECT 2856.670 375.740 2856.990 375.800 ;
        RECT 2856.670 37.980 2856.990 38.040 ;
        RECT 2863.110 37.980 2863.430 38.040 ;
        RECT 2856.670 37.840 2863.430 37.980 ;
        RECT 2856.670 37.780 2856.990 37.840 ;
        RECT 2863.110 37.780 2863.430 37.840 ;
      LAYER via ;
        RECT 1966.140 375.740 1966.400 376.000 ;
        RECT 2856.700 375.740 2856.960 376.000 ;
        RECT 2856.700 37.780 2856.960 38.040 ;
        RECT 2863.140 37.780 2863.400 38.040 ;
      LAYER met2 ;
        RECT 1966.270 510.340 1966.550 514.000 ;
        RECT 1966.200 510.000 1966.550 510.340 ;
        RECT 1966.200 376.030 1966.340 510.000 ;
        RECT 1966.140 375.710 1966.400 376.030 ;
        RECT 2856.700 375.710 2856.960 376.030 ;
        RECT 2856.760 38.070 2856.900 375.710 ;
        RECT 2856.700 37.750 2856.960 38.070 ;
        RECT 2863.140 37.750 2863.400 38.070 ;
        RECT 2863.200 2.400 2863.340 37.750 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 369.140 1980.230 369.200 ;
        RECT 2877.370 369.140 2877.690 369.200 ;
        RECT 1979.910 369.000 2877.690 369.140 ;
        RECT 1979.910 368.940 1980.230 369.000 ;
        RECT 2877.370 368.940 2877.690 369.000 ;
      LAYER via ;
        RECT 1979.940 368.940 1980.200 369.200 ;
        RECT 2877.400 368.940 2877.660 369.200 ;
      LAYER met2 ;
        RECT 1978.690 510.410 1978.970 514.000 ;
        RECT 1978.690 510.270 1980.140 510.410 ;
        RECT 1978.690 510.000 1978.970 510.270 ;
        RECT 1980.000 369.230 1980.140 510.270 ;
        RECT 1979.940 368.910 1980.200 369.230 ;
        RECT 2877.400 368.910 2877.660 369.230 ;
        RECT 2877.460 18.090 2877.600 368.910 ;
        RECT 2877.460 17.950 2881.280 18.090 ;
        RECT 2881.140 2.400 2881.280 17.950 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 79.460 1994.030 79.520 ;
        RECT 2894.850 79.460 2895.170 79.520 ;
        RECT 1993.710 79.320 2895.170 79.460 ;
        RECT 1993.710 79.260 1994.030 79.320 ;
        RECT 2894.850 79.260 2895.170 79.320 ;
        RECT 2894.850 17.580 2895.170 17.640 ;
        RECT 2898.990 17.580 2899.310 17.640 ;
        RECT 2894.850 17.440 2899.310 17.580 ;
        RECT 2894.850 17.380 2895.170 17.440 ;
        RECT 2898.990 17.380 2899.310 17.440 ;
      LAYER via ;
        RECT 1993.740 79.260 1994.000 79.520 ;
        RECT 2894.880 79.260 2895.140 79.520 ;
        RECT 2894.880 17.380 2895.140 17.640 ;
        RECT 2899.020 17.380 2899.280 17.640 ;
      LAYER met2 ;
        RECT 1991.110 510.410 1991.390 514.000 ;
        RECT 1991.110 510.270 1993.940 510.410 ;
        RECT 1991.110 510.000 1991.390 510.270 ;
        RECT 1993.800 79.550 1993.940 510.270 ;
        RECT 1993.740 79.230 1994.000 79.550 ;
        RECT 2894.880 79.230 2895.140 79.550 ;
        RECT 2894.940 17.670 2895.080 79.230 ;
        RECT 2894.880 17.350 2895.140 17.670 ;
        RECT 2899.020 17.350 2899.280 17.670 ;
        RECT 2899.080 2.400 2899.220 17.350 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 571.850 224.640 572.170 224.700 ;
        RECT 841.870 224.640 842.190 224.700 ;
        RECT 571.850 224.500 842.190 224.640 ;
        RECT 571.850 224.440 572.170 224.500 ;
        RECT 841.870 224.440 842.190 224.500 ;
      LAYER via ;
        RECT 571.880 224.440 572.140 224.700 ;
        RECT 841.900 224.440 842.160 224.700 ;
      LAYER met2 ;
        RECT 568.330 510.410 568.610 514.000 ;
        RECT 568.330 510.270 572.080 510.410 ;
        RECT 568.330 510.000 568.610 510.270 ;
        RECT 571.940 224.730 572.080 510.270 ;
        RECT 571.880 224.410 572.140 224.730 ;
        RECT 841.900 224.410 842.160 224.730 ;
        RECT 841.960 17.410 842.100 224.410 ;
        RECT 841.960 17.270 847.160 17.410 ;
        RECT 847.020 2.400 847.160 17.270 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.590 496.980 580.910 497.040 ;
        RECT 586.110 496.980 586.430 497.040 ;
        RECT 580.590 496.840 586.430 496.980 ;
        RECT 580.590 496.780 580.910 496.840 ;
        RECT 586.110 496.780 586.430 496.840 ;
        RECT 586.110 37.980 586.430 38.040 ;
        RECT 864.870 37.980 865.190 38.040 ;
        RECT 586.110 37.840 865.190 37.980 ;
        RECT 586.110 37.780 586.430 37.840 ;
        RECT 864.870 37.780 865.190 37.840 ;
      LAYER via ;
        RECT 580.620 496.780 580.880 497.040 ;
        RECT 586.140 496.780 586.400 497.040 ;
        RECT 586.140 37.780 586.400 38.040 ;
        RECT 864.900 37.780 865.160 38.040 ;
      LAYER met2 ;
        RECT 580.750 510.340 581.030 514.000 ;
        RECT 580.680 510.000 581.030 510.340 ;
        RECT 580.680 497.070 580.820 510.000 ;
        RECT 580.620 496.750 580.880 497.070 ;
        RECT 586.140 496.750 586.400 497.070 ;
        RECT 586.200 38.070 586.340 496.750 ;
        RECT 586.140 37.750 586.400 38.070 ;
        RECT 864.900 37.750 865.160 38.070 ;
        RECT 864.960 2.400 865.100 37.750 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 44.780 593.330 44.840 ;
        RECT 882.810 44.780 883.130 44.840 ;
        RECT 593.010 44.640 883.130 44.780 ;
        RECT 593.010 44.580 593.330 44.640 ;
        RECT 882.810 44.580 883.130 44.640 ;
      LAYER via ;
        RECT 593.040 44.580 593.300 44.840 ;
        RECT 882.840 44.580 883.100 44.840 ;
      LAYER met2 ;
        RECT 593.170 510.340 593.450 514.000 ;
        RECT 593.100 510.000 593.450 510.340 ;
        RECT 593.100 44.870 593.240 510.000 ;
        RECT 593.040 44.550 593.300 44.870 ;
        RECT 882.840 44.550 883.100 44.870 ;
        RECT 882.900 2.400 883.040 44.550 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 51.580 607.130 51.640 ;
        RECT 897.070 51.580 897.390 51.640 ;
        RECT 606.810 51.440 897.390 51.580 ;
        RECT 606.810 51.380 607.130 51.440 ;
        RECT 897.070 51.380 897.390 51.440 ;
      LAYER via ;
        RECT 606.840 51.380 607.100 51.640 ;
        RECT 897.100 51.380 897.360 51.640 ;
      LAYER met2 ;
        RECT 605.590 510.410 605.870 514.000 ;
        RECT 605.590 510.270 607.040 510.410 ;
        RECT 605.590 510.000 605.870 510.270 ;
        RECT 606.900 51.670 607.040 510.270 ;
        RECT 606.840 51.350 607.100 51.670 ;
        RECT 897.100 51.350 897.360 51.670 ;
        RECT 897.160 17.410 897.300 51.350 ;
        RECT 897.160 17.270 900.980 17.410 ;
        RECT 900.840 2.400 900.980 17.270 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 58.720 620.930 58.780 ;
        RECT 917.770 58.720 918.090 58.780 ;
        RECT 620.610 58.580 918.090 58.720 ;
        RECT 620.610 58.520 620.930 58.580 ;
        RECT 917.770 58.520 918.090 58.580 ;
      LAYER via ;
        RECT 620.640 58.520 620.900 58.780 ;
        RECT 917.800 58.520 918.060 58.780 ;
      LAYER met2 ;
        RECT 618.010 510.410 618.290 514.000 ;
        RECT 618.010 510.270 620.840 510.410 ;
        RECT 618.010 510.000 618.290 510.270 ;
        RECT 620.700 58.810 620.840 510.270 ;
        RECT 620.640 58.490 620.900 58.810 ;
        RECT 917.800 58.490 918.060 58.810 ;
        RECT 917.860 17.410 918.000 58.490 ;
        RECT 917.860 17.270 918.920 17.410 ;
        RECT 918.780 2.400 918.920 17.270 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 630.270 496.980 630.590 497.040 ;
        RECT 634.410 496.980 634.730 497.040 ;
        RECT 630.270 496.840 634.730 496.980 ;
        RECT 630.270 496.780 630.590 496.840 ;
        RECT 634.410 496.780 634.730 496.840 ;
        RECT 634.410 65.520 634.730 65.580 ;
        RECT 931.570 65.520 931.890 65.580 ;
        RECT 634.410 65.380 931.890 65.520 ;
        RECT 634.410 65.320 634.730 65.380 ;
        RECT 931.570 65.320 931.890 65.380 ;
      LAYER via ;
        RECT 630.300 496.780 630.560 497.040 ;
        RECT 634.440 496.780 634.700 497.040 ;
        RECT 634.440 65.320 634.700 65.580 ;
        RECT 931.600 65.320 931.860 65.580 ;
      LAYER met2 ;
        RECT 630.430 510.340 630.710 514.000 ;
        RECT 630.360 510.000 630.710 510.340 ;
        RECT 630.360 497.070 630.500 510.000 ;
        RECT 630.300 496.750 630.560 497.070 ;
        RECT 634.440 496.750 634.700 497.070 ;
        RECT 634.500 65.610 634.640 496.750 ;
        RECT 634.440 65.290 634.700 65.610 ;
        RECT 931.600 65.290 931.860 65.610 ;
        RECT 931.660 17.410 931.800 65.290 ;
        RECT 931.660 17.270 936.400 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 642.230 496.980 642.550 497.040 ;
        RECT 648.210 496.980 648.530 497.040 ;
        RECT 642.230 496.840 648.530 496.980 ;
        RECT 642.230 496.780 642.550 496.840 ;
        RECT 648.210 496.780 648.530 496.840 ;
        RECT 648.210 72.320 648.530 72.380 ;
        RECT 952.270 72.320 952.590 72.380 ;
        RECT 648.210 72.180 952.590 72.320 ;
        RECT 648.210 72.120 648.530 72.180 ;
        RECT 952.270 72.120 952.590 72.180 ;
      LAYER via ;
        RECT 642.260 496.780 642.520 497.040 ;
        RECT 648.240 496.780 648.500 497.040 ;
        RECT 648.240 72.120 648.500 72.380 ;
        RECT 952.300 72.120 952.560 72.380 ;
      LAYER met2 ;
        RECT 642.390 510.340 642.670 514.000 ;
        RECT 642.320 510.000 642.670 510.340 ;
        RECT 642.320 497.070 642.460 510.000 ;
        RECT 642.260 496.750 642.520 497.070 ;
        RECT 648.240 496.750 648.500 497.070 ;
        RECT 648.300 72.410 648.440 496.750 ;
        RECT 648.240 72.090 648.500 72.410 ;
        RECT 952.300 72.090 952.560 72.410 ;
        RECT 952.360 17.410 952.500 72.090 ;
        RECT 952.360 17.270 954.340 17.410 ;
        RECT 954.200 2.400 954.340 17.270 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 654.650 497.320 654.970 497.380 ;
        RECT 658.790 497.320 659.110 497.380 ;
        RECT 654.650 497.180 659.110 497.320 ;
        RECT 654.650 497.120 654.970 497.180 ;
        RECT 658.790 497.120 659.110 497.180 ;
        RECT 658.790 79.460 659.110 79.520 ;
        RECT 966.530 79.460 966.850 79.520 ;
        RECT 658.790 79.320 966.850 79.460 ;
        RECT 658.790 79.260 659.110 79.320 ;
        RECT 966.530 79.260 966.850 79.320 ;
      LAYER via ;
        RECT 654.680 497.120 654.940 497.380 ;
        RECT 658.820 497.120 659.080 497.380 ;
        RECT 658.820 79.260 659.080 79.520 ;
        RECT 966.560 79.260 966.820 79.520 ;
      LAYER met2 ;
        RECT 654.810 510.340 655.090 514.000 ;
        RECT 654.740 510.000 655.090 510.340 ;
        RECT 654.740 497.410 654.880 510.000 ;
        RECT 654.680 497.090 654.940 497.410 ;
        RECT 658.820 497.090 659.080 497.410 ;
        RECT 658.880 79.550 659.020 497.090 ;
        RECT 658.820 79.230 659.080 79.550 ;
        RECT 966.560 79.230 966.820 79.550 ;
        RECT 966.620 17.410 966.760 79.230 ;
        RECT 966.620 17.270 972.280 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 434.310 79.460 434.630 79.520 ;
        RECT 648.670 79.460 648.990 79.520 ;
        RECT 434.310 79.320 648.990 79.460 ;
        RECT 434.310 79.260 434.630 79.320 ;
        RECT 648.670 79.260 648.990 79.320 ;
      LAYER via ;
        RECT 434.340 79.260 434.600 79.520 ;
        RECT 648.700 79.260 648.960 79.520 ;
      LAYER met2 ;
        RECT 432.170 510.410 432.450 514.000 ;
        RECT 432.170 510.270 434.540 510.410 ;
        RECT 432.170 510.000 432.450 510.270 ;
        RECT 434.400 79.550 434.540 510.270 ;
        RECT 434.340 79.230 434.600 79.550 ;
        RECT 648.700 79.230 648.960 79.550 ;
        RECT 648.760 3.130 648.900 79.230 ;
        RECT 648.760 2.990 651.200 3.130 ;
        RECT 651.060 2.400 651.200 2.990 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 667.070 500.040 667.390 500.100 ;
        RECT 893.390 500.040 893.710 500.100 ;
        RECT 667.070 499.900 893.710 500.040 ;
        RECT 667.070 499.840 667.390 499.900 ;
        RECT 893.390 499.840 893.710 499.900 ;
        RECT 893.390 24.380 893.710 24.440 ;
        RECT 989.990 24.380 990.310 24.440 ;
        RECT 893.390 24.240 990.310 24.380 ;
        RECT 893.390 24.180 893.710 24.240 ;
        RECT 989.990 24.180 990.310 24.240 ;
      LAYER via ;
        RECT 667.100 499.840 667.360 500.100 ;
        RECT 893.420 499.840 893.680 500.100 ;
        RECT 893.420 24.180 893.680 24.440 ;
        RECT 990.020 24.180 990.280 24.440 ;
      LAYER met2 ;
        RECT 667.230 510.340 667.510 514.000 ;
        RECT 667.160 510.000 667.510 510.340 ;
        RECT 667.160 500.130 667.300 510.000 ;
        RECT 667.100 499.810 667.360 500.130 ;
        RECT 893.420 499.810 893.680 500.130 ;
        RECT 893.480 24.470 893.620 499.810 ;
        RECT 893.420 24.150 893.680 24.470 ;
        RECT 990.020 24.150 990.280 24.470 ;
        RECT 990.080 2.400 990.220 24.150 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 86.600 683.030 86.660 ;
        RECT 1007.930 86.600 1008.250 86.660 ;
        RECT 682.710 86.460 1008.250 86.600 ;
        RECT 682.710 86.400 683.030 86.460 ;
        RECT 1007.930 86.400 1008.250 86.460 ;
      LAYER via ;
        RECT 682.740 86.400 683.000 86.660 ;
        RECT 1007.960 86.400 1008.220 86.660 ;
      LAYER met2 ;
        RECT 679.650 510.410 679.930 514.000 ;
        RECT 679.650 510.270 682.940 510.410 ;
        RECT 679.650 510.000 679.930 510.270 ;
        RECT 682.800 86.690 682.940 510.270 ;
        RECT 682.740 86.370 683.000 86.690 ;
        RECT 1007.960 86.370 1008.220 86.690 ;
        RECT 1008.020 37.130 1008.160 86.370 ;
        RECT 1007.560 36.990 1008.160 37.130 ;
        RECT 1007.560 2.400 1007.700 36.990 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 691.910 496.980 692.230 497.040 ;
        RECT 696.510 496.980 696.830 497.040 ;
        RECT 691.910 496.840 696.830 496.980 ;
        RECT 691.910 496.780 692.230 496.840 ;
        RECT 696.510 496.780 696.830 496.840 ;
        RECT 696.510 93.060 696.830 93.120 ;
        RECT 1021.270 93.060 1021.590 93.120 ;
        RECT 696.510 92.920 1021.590 93.060 ;
        RECT 696.510 92.860 696.830 92.920 ;
        RECT 1021.270 92.860 1021.590 92.920 ;
        RECT 1021.270 62.120 1021.590 62.180 ;
        RECT 1025.410 62.120 1025.730 62.180 ;
        RECT 1021.270 61.980 1025.730 62.120 ;
        RECT 1021.270 61.920 1021.590 61.980 ;
        RECT 1025.410 61.920 1025.730 61.980 ;
      LAYER via ;
        RECT 691.940 496.780 692.200 497.040 ;
        RECT 696.540 496.780 696.800 497.040 ;
        RECT 696.540 92.860 696.800 93.120 ;
        RECT 1021.300 92.860 1021.560 93.120 ;
        RECT 1021.300 61.920 1021.560 62.180 ;
        RECT 1025.440 61.920 1025.700 62.180 ;
      LAYER met2 ;
        RECT 692.070 510.340 692.350 514.000 ;
        RECT 692.000 510.000 692.350 510.340 ;
        RECT 692.000 497.070 692.140 510.000 ;
        RECT 691.940 496.750 692.200 497.070 ;
        RECT 696.540 496.750 696.800 497.070 ;
        RECT 696.600 93.150 696.740 496.750 ;
        RECT 696.540 92.830 696.800 93.150 ;
        RECT 1021.300 92.830 1021.560 93.150 ;
        RECT 1021.360 62.210 1021.500 92.830 ;
        RECT 1021.300 61.890 1021.560 62.210 ;
        RECT 1025.440 61.890 1025.700 62.210 ;
        RECT 1025.500 2.400 1025.640 61.890 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 496.980 704.650 497.040 ;
        RECT 710.310 496.980 710.630 497.040 ;
        RECT 704.330 496.840 710.630 496.980 ;
        RECT 704.330 496.780 704.650 496.840 ;
        RECT 710.310 496.780 710.630 496.840 ;
        RECT 710.310 100.200 710.630 100.260 ;
        RECT 1041.970 100.200 1042.290 100.260 ;
        RECT 710.310 100.060 1042.290 100.200 ;
        RECT 710.310 100.000 710.630 100.060 ;
        RECT 1041.970 100.000 1042.290 100.060 ;
      LAYER via ;
        RECT 704.360 496.780 704.620 497.040 ;
        RECT 710.340 496.780 710.600 497.040 ;
        RECT 710.340 100.000 710.600 100.260 ;
        RECT 1042.000 100.000 1042.260 100.260 ;
      LAYER met2 ;
        RECT 704.490 510.340 704.770 514.000 ;
        RECT 704.420 510.000 704.770 510.340 ;
        RECT 704.420 497.070 704.560 510.000 ;
        RECT 704.360 496.750 704.620 497.070 ;
        RECT 710.340 496.750 710.600 497.070 ;
        RECT 710.400 100.290 710.540 496.750 ;
        RECT 710.340 99.970 710.600 100.290 ;
        RECT 1042.000 99.970 1042.260 100.290 ;
        RECT 1042.060 16.730 1042.200 99.970 ;
        RECT 1042.060 16.590 1043.580 16.730 ;
        RECT 1043.440 2.400 1043.580 16.590 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 107.000 717.530 107.060 ;
        RECT 1055.770 107.000 1056.090 107.060 ;
        RECT 717.210 106.860 1056.090 107.000 ;
        RECT 717.210 106.800 717.530 106.860 ;
        RECT 1055.770 106.800 1056.090 106.860 ;
      LAYER via ;
        RECT 717.240 106.800 717.500 107.060 ;
        RECT 1055.800 106.800 1056.060 107.060 ;
      LAYER met2 ;
        RECT 716.910 510.340 717.190 514.000 ;
        RECT 716.840 510.000 717.190 510.340 ;
        RECT 716.840 497.490 716.980 510.000 ;
        RECT 716.840 497.350 717.440 497.490 ;
        RECT 717.300 107.090 717.440 497.350 ;
        RECT 717.240 106.770 717.500 107.090 ;
        RECT 1055.800 106.770 1056.060 107.090 ;
        RECT 1055.860 17.410 1056.000 106.770 ;
        RECT 1055.860 17.270 1061.520 17.410 ;
        RECT 1061.380 2.400 1061.520 17.270 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 729.170 493.240 729.490 493.300 ;
        RECT 1076.470 493.240 1076.790 493.300 ;
        RECT 729.170 493.100 1076.790 493.240 ;
        RECT 729.170 493.040 729.490 493.100 ;
        RECT 1076.470 493.040 1076.790 493.100 ;
      LAYER via ;
        RECT 729.200 493.040 729.460 493.300 ;
        RECT 1076.500 493.040 1076.760 493.300 ;
      LAYER met2 ;
        RECT 729.330 510.340 729.610 514.000 ;
        RECT 729.260 510.000 729.610 510.340 ;
        RECT 729.260 493.330 729.400 510.000 ;
        RECT 729.200 493.010 729.460 493.330 ;
        RECT 1076.500 493.010 1076.760 493.330 ;
        RECT 1076.560 17.410 1076.700 493.010 ;
        RECT 1076.560 17.270 1079.460 17.410 ;
        RECT 1079.320 2.400 1079.460 17.270 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 744.810 113.800 745.130 113.860 ;
        RECT 1090.730 113.800 1091.050 113.860 ;
        RECT 744.810 113.660 1091.050 113.800 ;
        RECT 744.810 113.600 745.130 113.660 ;
        RECT 1090.730 113.600 1091.050 113.660 ;
        RECT 1090.730 17.920 1091.050 17.980 ;
        RECT 1096.710 17.920 1097.030 17.980 ;
        RECT 1090.730 17.780 1097.030 17.920 ;
        RECT 1090.730 17.720 1091.050 17.780 ;
        RECT 1096.710 17.720 1097.030 17.780 ;
      LAYER via ;
        RECT 744.840 113.600 745.100 113.860 ;
        RECT 1090.760 113.600 1091.020 113.860 ;
        RECT 1090.760 17.720 1091.020 17.980 ;
        RECT 1096.740 17.720 1097.000 17.980 ;
      LAYER met2 ;
        RECT 741.750 510.410 742.030 514.000 ;
        RECT 741.750 510.270 745.040 510.410 ;
        RECT 741.750 510.000 742.030 510.270 ;
        RECT 744.900 113.890 745.040 510.270 ;
        RECT 744.840 113.570 745.100 113.890 ;
        RECT 1090.760 113.570 1091.020 113.890 ;
        RECT 1090.820 18.010 1090.960 113.570 ;
        RECT 1090.760 17.690 1091.020 18.010 ;
        RECT 1096.740 17.690 1097.000 18.010 ;
        RECT 1096.800 2.400 1096.940 17.690 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.550 498.680 753.870 498.740 ;
        RECT 758.610 498.680 758.930 498.740 ;
        RECT 753.550 498.540 758.930 498.680 ;
        RECT 753.550 498.480 753.870 498.540 ;
        RECT 758.610 498.480 758.930 498.540 ;
        RECT 758.610 120.600 758.930 120.660 ;
        RECT 1110.970 120.600 1111.290 120.660 ;
        RECT 758.610 120.460 1111.290 120.600 ;
        RECT 758.610 120.400 758.930 120.460 ;
        RECT 1110.970 120.400 1111.290 120.460 ;
      LAYER via ;
        RECT 753.580 498.480 753.840 498.740 ;
        RECT 758.640 498.480 758.900 498.740 ;
        RECT 758.640 120.400 758.900 120.660 ;
        RECT 1111.000 120.400 1111.260 120.660 ;
      LAYER met2 ;
        RECT 753.710 510.340 753.990 514.000 ;
        RECT 753.640 510.000 753.990 510.340 ;
        RECT 753.640 498.770 753.780 510.000 ;
        RECT 753.580 498.450 753.840 498.770 ;
        RECT 758.640 498.450 758.900 498.770 ;
        RECT 758.700 120.690 758.840 498.450 ;
        RECT 758.640 120.370 758.900 120.690 ;
        RECT 1111.000 120.370 1111.260 120.690 ;
        RECT 1111.060 17.410 1111.200 120.370 ;
        RECT 1111.060 17.270 1114.880 17.410 ;
        RECT 1114.740 2.400 1114.880 17.270 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.970 503.440 766.290 503.500 ;
        RECT 772.410 503.440 772.730 503.500 ;
        RECT 765.970 503.300 772.730 503.440 ;
        RECT 765.970 503.240 766.290 503.300 ;
        RECT 772.410 503.240 772.730 503.300 ;
        RECT 772.410 127.740 772.730 127.800 ;
        RECT 1131.670 127.740 1131.990 127.800 ;
        RECT 772.410 127.600 1131.990 127.740 ;
        RECT 772.410 127.540 772.730 127.600 ;
        RECT 1131.670 127.540 1131.990 127.600 ;
      LAYER via ;
        RECT 766.000 503.240 766.260 503.500 ;
        RECT 772.440 503.240 772.700 503.500 ;
        RECT 772.440 127.540 772.700 127.800 ;
        RECT 1131.700 127.540 1131.960 127.800 ;
      LAYER met2 ;
        RECT 766.130 510.340 766.410 514.000 ;
        RECT 766.060 510.000 766.410 510.340 ;
        RECT 766.060 503.530 766.200 510.000 ;
        RECT 766.000 503.210 766.260 503.530 ;
        RECT 772.440 503.210 772.700 503.530 ;
        RECT 772.500 127.830 772.640 503.210 ;
        RECT 772.440 127.510 772.700 127.830 ;
        RECT 1131.700 127.510 1131.960 127.830 ;
        RECT 1131.760 17.410 1131.900 127.510 ;
        RECT 1131.760 17.270 1132.820 17.410 ;
        RECT 1132.680 2.400 1132.820 17.270 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 134.540 779.630 134.600 ;
        RECT 1145.470 134.540 1145.790 134.600 ;
        RECT 779.310 134.400 1145.790 134.540 ;
        RECT 779.310 134.340 779.630 134.400 ;
        RECT 1145.470 134.340 1145.790 134.400 ;
      LAYER via ;
        RECT 779.340 134.340 779.600 134.600 ;
        RECT 1145.500 134.340 1145.760 134.600 ;
      LAYER met2 ;
        RECT 778.550 510.410 778.830 514.000 ;
        RECT 778.550 510.270 779.540 510.410 ;
        RECT 778.550 510.000 778.830 510.270 ;
        RECT 779.400 134.630 779.540 510.270 ;
        RECT 779.340 134.310 779.600 134.630 ;
        RECT 1145.500 134.310 1145.760 134.630 ;
        RECT 1145.560 17.410 1145.700 134.310 ;
        RECT 1145.560 17.270 1150.760 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 444.430 496.980 444.750 497.040 ;
        RECT 448.110 496.980 448.430 497.040 ;
        RECT 444.430 496.840 448.430 496.980 ;
        RECT 444.430 496.780 444.750 496.840 ;
        RECT 448.110 496.780 448.430 496.840 ;
        RECT 448.110 86.260 448.430 86.320 ;
        RECT 662.930 86.260 663.250 86.320 ;
        RECT 448.110 86.120 663.250 86.260 ;
        RECT 448.110 86.060 448.430 86.120 ;
        RECT 662.930 86.060 663.250 86.120 ;
        RECT 662.930 38.320 663.250 38.380 ;
        RECT 668.910 38.320 669.230 38.380 ;
        RECT 662.930 38.180 669.230 38.320 ;
        RECT 662.930 38.120 663.250 38.180 ;
        RECT 668.910 38.120 669.230 38.180 ;
      LAYER via ;
        RECT 444.460 496.780 444.720 497.040 ;
        RECT 448.140 496.780 448.400 497.040 ;
        RECT 448.140 86.060 448.400 86.320 ;
        RECT 662.960 86.060 663.220 86.320 ;
        RECT 662.960 38.120 663.220 38.380 ;
        RECT 668.940 38.120 669.200 38.380 ;
      LAYER met2 ;
        RECT 444.590 510.340 444.870 514.000 ;
        RECT 444.520 510.000 444.870 510.340 ;
        RECT 444.520 497.070 444.660 510.000 ;
        RECT 444.460 496.750 444.720 497.070 ;
        RECT 448.140 496.750 448.400 497.070 ;
        RECT 448.200 86.350 448.340 496.750 ;
        RECT 448.140 86.030 448.400 86.350 ;
        RECT 662.960 86.030 663.220 86.350 ;
        RECT 663.020 38.410 663.160 86.030 ;
        RECT 662.960 38.090 663.220 38.410 ;
        RECT 668.940 38.090 669.200 38.410 ;
        RECT 669.000 2.400 669.140 38.090 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 141.340 793.430 141.400 ;
        RECT 1166.170 141.340 1166.490 141.400 ;
        RECT 793.110 141.200 1166.490 141.340 ;
        RECT 793.110 141.140 793.430 141.200 ;
        RECT 1166.170 141.140 1166.490 141.200 ;
      LAYER via ;
        RECT 793.140 141.140 793.400 141.400 ;
        RECT 1166.200 141.140 1166.460 141.400 ;
      LAYER met2 ;
        RECT 790.970 510.410 791.250 514.000 ;
        RECT 790.970 510.270 793.340 510.410 ;
        RECT 790.970 510.000 791.250 510.270 ;
        RECT 793.200 141.430 793.340 510.270 ;
        RECT 793.140 141.110 793.400 141.430 ;
        RECT 1166.200 141.110 1166.460 141.430 ;
        RECT 1166.260 17.410 1166.400 141.110 ;
        RECT 1166.260 17.270 1168.700 17.410 ;
        RECT 1168.560 2.400 1168.700 17.270 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 803.230 496.980 803.550 497.040 ;
        RECT 806.910 496.980 807.230 497.040 ;
        RECT 803.230 496.840 807.230 496.980 ;
        RECT 803.230 496.780 803.550 496.840 ;
        RECT 806.910 496.780 807.230 496.840 ;
        RECT 806.910 31.180 807.230 31.240 ;
        RECT 1185.950 31.180 1186.270 31.240 ;
        RECT 806.910 31.040 1186.270 31.180 ;
        RECT 806.910 30.980 807.230 31.040 ;
        RECT 1185.950 30.980 1186.270 31.040 ;
      LAYER via ;
        RECT 803.260 496.780 803.520 497.040 ;
        RECT 806.940 496.780 807.200 497.040 ;
        RECT 806.940 30.980 807.200 31.240 ;
        RECT 1185.980 30.980 1186.240 31.240 ;
      LAYER met2 ;
        RECT 803.390 510.340 803.670 514.000 ;
        RECT 803.320 510.000 803.670 510.340 ;
        RECT 803.320 497.070 803.460 510.000 ;
        RECT 803.260 496.750 803.520 497.070 ;
        RECT 806.940 496.750 807.200 497.070 ;
        RECT 807.000 31.270 807.140 496.750 ;
        RECT 806.940 30.950 807.200 31.270 ;
        RECT 1185.980 30.950 1186.240 31.270 ;
        RECT 1186.040 2.400 1186.180 30.950 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 815.650 486.780 815.970 486.840 ;
        RECT 1200.670 486.780 1200.990 486.840 ;
        RECT 815.650 486.640 1200.990 486.780 ;
        RECT 815.650 486.580 815.970 486.640 ;
        RECT 1200.670 486.580 1200.990 486.640 ;
      LAYER via ;
        RECT 815.680 486.580 815.940 486.840 ;
        RECT 1200.700 486.580 1200.960 486.840 ;
      LAYER met2 ;
        RECT 815.810 510.340 816.090 514.000 ;
        RECT 815.740 510.000 816.090 510.340 ;
        RECT 815.740 486.870 815.880 510.000 ;
        RECT 815.680 486.550 815.940 486.870 ;
        RECT 1200.700 486.550 1200.960 486.870 ;
        RECT 1200.760 17.410 1200.900 486.550 ;
        RECT 1200.760 17.270 1204.120 17.410 ;
        RECT 1203.980 2.400 1204.120 17.270 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 828.070 500.720 828.390 500.780 ;
        RECT 872.690 500.720 873.010 500.780 ;
        RECT 828.070 500.580 873.010 500.720 ;
        RECT 828.070 500.520 828.390 500.580 ;
        RECT 872.690 500.520 873.010 500.580 ;
        RECT 872.690 38.660 873.010 38.720 ;
        RECT 1221.830 38.660 1222.150 38.720 ;
        RECT 872.690 38.520 1222.150 38.660 ;
        RECT 872.690 38.460 873.010 38.520 ;
        RECT 1221.830 38.460 1222.150 38.520 ;
      LAYER via ;
        RECT 828.100 500.520 828.360 500.780 ;
        RECT 872.720 500.520 872.980 500.780 ;
        RECT 872.720 38.460 872.980 38.720 ;
        RECT 1221.860 38.460 1222.120 38.720 ;
      LAYER met2 ;
        RECT 828.230 510.340 828.510 514.000 ;
        RECT 828.160 510.000 828.510 510.340 ;
        RECT 828.160 500.810 828.300 510.000 ;
        RECT 828.100 500.490 828.360 500.810 ;
        RECT 872.720 500.490 872.980 500.810 ;
        RECT 872.780 38.750 872.920 500.490 ;
        RECT 872.720 38.430 872.980 38.750 ;
        RECT 1221.860 38.430 1222.120 38.750 ;
        RECT 1221.920 2.400 1222.060 38.430 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 148.140 841.730 148.200 ;
        RECT 1235.170 148.140 1235.490 148.200 ;
        RECT 841.410 148.000 1235.490 148.140 ;
        RECT 841.410 147.940 841.730 148.000 ;
        RECT 1235.170 147.940 1235.490 148.000 ;
      LAYER via ;
        RECT 841.440 147.940 841.700 148.200 ;
        RECT 1235.200 147.940 1235.460 148.200 ;
      LAYER met2 ;
        RECT 840.650 510.410 840.930 514.000 ;
        RECT 840.650 510.270 841.640 510.410 ;
        RECT 840.650 510.000 840.930 510.270 ;
        RECT 841.500 148.230 841.640 510.270 ;
        RECT 841.440 147.910 841.700 148.230 ;
        RECT 1235.200 147.910 1235.460 148.230 ;
        RECT 1235.260 17.410 1235.400 147.910 ;
        RECT 1235.260 17.270 1240.000 17.410 ;
        RECT 1239.860 2.400 1240.000 17.270 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.210 45.460 855.530 45.520 ;
        RECT 1257.250 45.460 1257.570 45.520 ;
        RECT 855.210 45.320 1257.570 45.460 ;
        RECT 855.210 45.260 855.530 45.320 ;
        RECT 1257.250 45.260 1257.570 45.320 ;
      LAYER via ;
        RECT 855.240 45.260 855.500 45.520 ;
        RECT 1257.280 45.260 1257.540 45.520 ;
      LAYER met2 ;
        RECT 853.070 510.410 853.350 514.000 ;
        RECT 853.070 510.270 855.440 510.410 ;
        RECT 853.070 510.000 853.350 510.270 ;
        RECT 855.300 45.550 855.440 510.270 ;
        RECT 855.240 45.230 855.500 45.550 ;
        RECT 1257.280 45.230 1257.540 45.550 ;
        RECT 1257.340 2.400 1257.480 45.230 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 865.330 496.980 865.650 497.040 ;
        RECT 869.010 496.980 869.330 497.040 ;
        RECT 865.330 496.840 869.330 496.980 ;
        RECT 865.330 496.780 865.650 496.840 ;
        RECT 869.010 496.780 869.330 496.840 ;
        RECT 869.010 155.280 869.330 155.340 ;
        RECT 1269.670 155.280 1269.990 155.340 ;
        RECT 869.010 155.140 1269.990 155.280 ;
        RECT 869.010 155.080 869.330 155.140 ;
        RECT 1269.670 155.080 1269.990 155.140 ;
      LAYER via ;
        RECT 865.360 496.780 865.620 497.040 ;
        RECT 869.040 496.780 869.300 497.040 ;
        RECT 869.040 155.080 869.300 155.340 ;
        RECT 1269.700 155.080 1269.960 155.340 ;
      LAYER met2 ;
        RECT 865.490 510.340 865.770 514.000 ;
        RECT 865.420 510.000 865.770 510.340 ;
        RECT 865.420 497.070 865.560 510.000 ;
        RECT 865.360 496.750 865.620 497.070 ;
        RECT 869.040 496.750 869.300 497.070 ;
        RECT 869.100 155.370 869.240 496.750 ;
        RECT 869.040 155.050 869.300 155.370 ;
        RECT 1269.700 155.050 1269.960 155.370 ;
        RECT 1269.760 17.410 1269.900 155.050 ;
        RECT 1269.760 17.270 1275.420 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 877.290 496.980 877.610 497.040 ;
        RECT 882.810 496.980 883.130 497.040 ;
        RECT 877.290 496.840 883.130 496.980 ;
        RECT 877.290 496.780 877.610 496.840 ;
        RECT 882.810 496.780 883.130 496.840 ;
        RECT 882.810 162.080 883.130 162.140 ;
        RECT 1290.370 162.080 1290.690 162.140 ;
        RECT 882.810 161.940 1290.690 162.080 ;
        RECT 882.810 161.880 883.130 161.940 ;
        RECT 1290.370 161.880 1290.690 161.940 ;
      LAYER via ;
        RECT 877.320 496.780 877.580 497.040 ;
        RECT 882.840 496.780 883.100 497.040 ;
        RECT 882.840 161.880 883.100 162.140 ;
        RECT 1290.400 161.880 1290.660 162.140 ;
      LAYER met2 ;
        RECT 877.450 510.340 877.730 514.000 ;
        RECT 877.380 510.000 877.730 510.340 ;
        RECT 877.380 497.070 877.520 510.000 ;
        RECT 877.320 496.750 877.580 497.070 ;
        RECT 882.840 496.750 883.100 497.070 ;
        RECT 882.900 162.170 883.040 496.750 ;
        RECT 882.840 161.850 883.100 162.170 ;
        RECT 1290.400 161.850 1290.660 162.170 ;
        RECT 1290.460 17.410 1290.600 161.850 ;
        RECT 1290.460 17.270 1293.360 17.410 ;
        RECT 1293.220 2.400 1293.360 17.270 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 889.710 168.880 890.030 168.940 ;
        RECT 1311.530 168.880 1311.850 168.940 ;
        RECT 889.710 168.740 1311.850 168.880 ;
        RECT 889.710 168.680 890.030 168.740 ;
        RECT 1311.530 168.680 1311.850 168.740 ;
      LAYER via ;
        RECT 889.740 168.680 890.000 168.940 ;
        RECT 1311.560 168.680 1311.820 168.940 ;
      LAYER met2 ;
        RECT 889.870 510.340 890.150 514.000 ;
        RECT 889.800 510.000 890.150 510.340 ;
        RECT 889.800 168.970 889.940 510.000 ;
        RECT 889.740 168.650 890.000 168.970 ;
        RECT 1311.560 168.650 1311.820 168.970 ;
        RECT 1311.620 17.410 1311.760 168.650 ;
        RECT 1311.160 17.270 1311.760 17.410 ;
        RECT 1311.160 2.400 1311.300 17.270 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 902.130 500.720 902.450 500.780 ;
        RECT 1017.590 500.720 1017.910 500.780 ;
        RECT 902.130 500.580 1017.910 500.720 ;
        RECT 902.130 500.520 902.450 500.580 ;
        RECT 1017.590 500.520 1017.910 500.580 ;
        RECT 1017.590 24.040 1017.910 24.100 ;
        RECT 1329.010 24.040 1329.330 24.100 ;
        RECT 1017.590 23.900 1329.330 24.040 ;
        RECT 1017.590 23.840 1017.910 23.900 ;
        RECT 1329.010 23.840 1329.330 23.900 ;
      LAYER via ;
        RECT 902.160 500.520 902.420 500.780 ;
        RECT 1017.620 500.520 1017.880 500.780 ;
        RECT 1017.620 23.840 1017.880 24.100 ;
        RECT 1329.040 23.840 1329.300 24.100 ;
      LAYER met2 ;
        RECT 902.290 510.340 902.570 514.000 ;
        RECT 902.220 510.000 902.570 510.340 ;
        RECT 902.220 500.810 902.360 510.000 ;
        RECT 902.160 500.490 902.420 500.810 ;
        RECT 1017.620 500.490 1017.880 500.810 ;
        RECT 1017.680 24.130 1017.820 500.490 ;
        RECT 1017.620 23.810 1017.880 24.130 ;
        RECT 1329.040 23.810 1329.300 24.130 ;
        RECT 1329.100 2.400 1329.240 23.810 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 456.850 493.240 457.170 493.300 ;
        RECT 461.910 493.240 462.230 493.300 ;
        RECT 456.850 493.100 462.230 493.240 ;
        RECT 456.850 493.040 457.170 493.100 ;
        RECT 461.910 493.040 462.230 493.100 ;
        RECT 461.910 93.060 462.230 93.120 ;
        RECT 683.170 93.060 683.490 93.120 ;
        RECT 461.910 92.920 683.490 93.060 ;
        RECT 461.910 92.860 462.230 92.920 ;
        RECT 683.170 92.860 683.490 92.920 ;
        RECT 683.170 62.120 683.490 62.180 ;
        RECT 685.930 62.120 686.250 62.180 ;
        RECT 683.170 61.980 686.250 62.120 ;
        RECT 683.170 61.920 683.490 61.980 ;
        RECT 685.930 61.920 686.250 61.980 ;
      LAYER via ;
        RECT 456.880 493.040 457.140 493.300 ;
        RECT 461.940 493.040 462.200 493.300 ;
        RECT 461.940 92.860 462.200 93.120 ;
        RECT 683.200 92.860 683.460 93.120 ;
        RECT 683.200 61.920 683.460 62.180 ;
        RECT 685.960 61.920 686.220 62.180 ;
      LAYER met2 ;
        RECT 457.010 510.340 457.290 514.000 ;
        RECT 456.940 510.000 457.290 510.340 ;
        RECT 456.940 493.330 457.080 510.000 ;
        RECT 456.880 493.010 457.140 493.330 ;
        RECT 461.940 493.010 462.200 493.330 ;
        RECT 462.000 93.150 462.140 493.010 ;
        RECT 461.940 92.830 462.200 93.150 ;
        RECT 683.200 92.830 683.460 93.150 ;
        RECT 683.260 62.210 683.400 92.830 ;
        RECT 683.200 61.890 683.460 62.210 ;
        RECT 685.960 61.890 686.220 62.210 ;
        RECT 686.020 61.610 686.160 61.890 ;
        RECT 686.020 61.470 686.620 61.610 ;
        RECT 686.480 2.400 686.620 61.470 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 51.920 917.630 51.980 ;
        RECT 1346.490 51.920 1346.810 51.980 ;
        RECT 917.310 51.780 1346.810 51.920 ;
        RECT 917.310 51.720 917.630 51.780 ;
        RECT 1346.490 51.720 1346.810 51.780 ;
      LAYER via ;
        RECT 917.340 51.720 917.600 51.980 ;
        RECT 1346.520 51.720 1346.780 51.980 ;
      LAYER met2 ;
        RECT 914.710 510.410 914.990 514.000 ;
        RECT 914.710 510.270 917.540 510.410 ;
        RECT 914.710 510.000 914.990 510.270 ;
        RECT 917.400 52.010 917.540 510.270 ;
        RECT 917.340 51.690 917.600 52.010 ;
        RECT 1346.520 51.690 1346.780 52.010 ;
        RECT 1346.580 2.400 1346.720 51.690 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 926.970 496.980 927.290 497.040 ;
        RECT 931.110 496.980 931.430 497.040 ;
        RECT 926.970 496.840 931.430 496.980 ;
        RECT 926.970 496.780 927.290 496.840 ;
        RECT 931.110 496.780 931.430 496.840 ;
        RECT 931.110 59.400 931.430 59.460 ;
        RECT 1364.430 59.400 1364.750 59.460 ;
        RECT 931.110 59.260 1364.750 59.400 ;
        RECT 931.110 59.200 931.430 59.260 ;
        RECT 1364.430 59.200 1364.750 59.260 ;
      LAYER via ;
        RECT 927.000 496.780 927.260 497.040 ;
        RECT 931.140 496.780 931.400 497.040 ;
        RECT 931.140 59.200 931.400 59.460 ;
        RECT 1364.460 59.200 1364.720 59.460 ;
      LAYER met2 ;
        RECT 927.130 510.340 927.410 514.000 ;
        RECT 927.060 510.000 927.410 510.340 ;
        RECT 927.060 497.070 927.200 510.000 ;
        RECT 927.000 496.750 927.260 497.070 ;
        RECT 931.140 496.750 931.400 497.070 ;
        RECT 931.200 59.490 931.340 496.750 ;
        RECT 931.140 59.170 931.400 59.490 ;
        RECT 1364.460 59.170 1364.720 59.490 ;
        RECT 1364.520 2.400 1364.660 59.170 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 939.390 496.980 939.710 497.040 ;
        RECT 944.910 496.980 945.230 497.040 ;
        RECT 939.390 496.840 945.230 496.980 ;
        RECT 939.390 496.780 939.710 496.840 ;
        RECT 944.910 496.780 945.230 496.840 ;
        RECT 944.910 65.860 945.230 65.920 ;
        RECT 1380.070 65.860 1380.390 65.920 ;
        RECT 944.910 65.720 1380.390 65.860 ;
        RECT 944.910 65.660 945.230 65.720 ;
        RECT 1380.070 65.660 1380.390 65.720 ;
      LAYER via ;
        RECT 939.420 496.780 939.680 497.040 ;
        RECT 944.940 496.780 945.200 497.040 ;
        RECT 944.940 65.660 945.200 65.920 ;
        RECT 1380.100 65.660 1380.360 65.920 ;
      LAYER met2 ;
        RECT 939.550 510.340 939.830 514.000 ;
        RECT 939.480 510.000 939.830 510.340 ;
        RECT 939.480 497.070 939.620 510.000 ;
        RECT 939.420 496.750 939.680 497.070 ;
        RECT 944.940 496.750 945.200 497.070 ;
        RECT 945.000 65.950 945.140 496.750 ;
        RECT 944.940 65.630 945.200 65.950 ;
        RECT 1380.100 65.630 1380.360 65.950 ;
        RECT 1380.160 17.410 1380.300 65.630 ;
        RECT 1380.160 17.270 1382.600 17.410 ;
        RECT 1382.460 2.400 1382.600 17.270 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 176.360 952.130 176.420 ;
        RECT 1394.330 176.360 1394.650 176.420 ;
        RECT 951.810 176.220 1394.650 176.360 ;
        RECT 951.810 176.160 952.130 176.220 ;
        RECT 1394.330 176.160 1394.650 176.220 ;
        RECT 1394.330 17.920 1394.650 17.980 ;
        RECT 1400.310 17.920 1400.630 17.980 ;
        RECT 1394.330 17.780 1400.630 17.920 ;
        RECT 1394.330 17.720 1394.650 17.780 ;
        RECT 1400.310 17.720 1400.630 17.780 ;
      LAYER via ;
        RECT 951.840 176.160 952.100 176.420 ;
        RECT 1394.360 176.160 1394.620 176.420 ;
        RECT 1394.360 17.720 1394.620 17.980 ;
        RECT 1400.340 17.720 1400.600 17.980 ;
      LAYER met2 ;
        RECT 951.970 510.340 952.250 514.000 ;
        RECT 951.900 510.000 952.250 510.340 ;
        RECT 951.900 176.450 952.040 510.000 ;
        RECT 951.840 176.130 952.100 176.450 ;
        RECT 1394.360 176.130 1394.620 176.450 ;
        RECT 1394.420 18.010 1394.560 176.130 ;
        RECT 1394.360 17.690 1394.620 18.010 ;
        RECT 1400.340 17.690 1400.600 18.010 ;
        RECT 1400.400 2.400 1400.540 17.690 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 965.610 72.660 965.930 72.720 ;
        RECT 1414.570 72.660 1414.890 72.720 ;
        RECT 965.610 72.520 1414.890 72.660 ;
        RECT 965.610 72.460 965.930 72.520 ;
        RECT 1414.570 72.460 1414.890 72.520 ;
      LAYER via ;
        RECT 965.640 72.460 965.900 72.720 ;
        RECT 1414.600 72.460 1414.860 72.720 ;
      LAYER met2 ;
        RECT 964.390 510.410 964.670 514.000 ;
        RECT 964.390 510.270 965.840 510.410 ;
        RECT 964.390 510.000 964.670 510.270 ;
        RECT 965.700 72.750 965.840 510.270 ;
        RECT 965.640 72.430 965.900 72.750 ;
        RECT 1414.600 72.430 1414.860 72.750 ;
        RECT 1414.660 17.410 1414.800 72.430 ;
        RECT 1414.660 17.270 1418.480 17.410 ;
        RECT 1418.340 2.400 1418.480 17.270 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.410 79.800 979.730 79.860 ;
        RECT 1435.730 79.800 1436.050 79.860 ;
        RECT 979.410 79.660 1436.050 79.800 ;
        RECT 979.410 79.600 979.730 79.660 ;
        RECT 1435.730 79.600 1436.050 79.660 ;
      LAYER via ;
        RECT 979.440 79.600 979.700 79.860 ;
        RECT 1435.760 79.600 1436.020 79.860 ;
      LAYER met2 ;
        RECT 976.810 510.410 977.090 514.000 ;
        RECT 976.810 510.270 979.640 510.410 ;
        RECT 976.810 510.000 977.090 510.270 ;
        RECT 979.500 79.890 979.640 510.270 ;
        RECT 979.440 79.570 979.700 79.890 ;
        RECT 1435.760 79.570 1436.020 79.890 ;
        RECT 1435.820 2.400 1435.960 79.570 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1335.065 448.205 1335.235 483.055 ;
        RECT 1335.525 386.325 1335.695 400.775 ;
        RECT 1335.525 338.045 1335.695 352.155 ;
        RECT 1335.525 289.765 1335.695 313.735 ;
        RECT 1335.525 241.485 1335.695 255.595 ;
        RECT 1335.065 193.205 1335.235 207.655 ;
        RECT 1335.525 96.645 1335.695 144.755 ;
      LAYER mcon ;
        RECT 1335.065 482.885 1335.235 483.055 ;
        RECT 1335.525 400.605 1335.695 400.775 ;
        RECT 1335.525 351.985 1335.695 352.155 ;
        RECT 1335.525 313.565 1335.695 313.735 ;
        RECT 1335.525 255.425 1335.695 255.595 ;
        RECT 1335.065 207.485 1335.235 207.655 ;
        RECT 1335.525 144.585 1335.695 144.755 ;
      LAYER met1 ;
        RECT 988.610 500.040 988.930 500.100 ;
        RECT 1334.990 500.040 1335.310 500.100 ;
        RECT 988.610 499.900 1335.310 500.040 ;
        RECT 988.610 499.840 988.930 499.900 ;
        RECT 1334.990 499.840 1335.310 499.900 ;
        RECT 1334.990 483.040 1335.310 483.100 ;
        RECT 1334.795 482.900 1335.310 483.040 ;
        RECT 1334.990 482.840 1335.310 482.900 ;
        RECT 1334.990 448.360 1335.310 448.420 ;
        RECT 1334.795 448.220 1335.310 448.360 ;
        RECT 1334.990 448.160 1335.310 448.220 ;
        RECT 1335.450 400.760 1335.770 400.820 ;
        RECT 1335.255 400.620 1335.770 400.760 ;
        RECT 1335.450 400.560 1335.770 400.620 ;
        RECT 1335.450 386.480 1335.770 386.540 ;
        RECT 1335.255 386.340 1335.770 386.480 ;
        RECT 1335.450 386.280 1335.770 386.340 ;
        RECT 1335.450 352.140 1335.770 352.200 ;
        RECT 1335.255 352.000 1335.770 352.140 ;
        RECT 1335.450 351.940 1335.770 352.000 ;
        RECT 1335.450 338.200 1335.770 338.260 ;
        RECT 1335.255 338.060 1335.770 338.200 ;
        RECT 1335.450 338.000 1335.770 338.060 ;
        RECT 1335.450 313.720 1335.770 313.780 ;
        RECT 1335.255 313.580 1335.770 313.720 ;
        RECT 1335.450 313.520 1335.770 313.580 ;
        RECT 1335.450 289.920 1335.770 289.980 ;
        RECT 1335.255 289.780 1335.770 289.920 ;
        RECT 1335.450 289.720 1335.770 289.780 ;
        RECT 1335.450 255.580 1335.770 255.640 ;
        RECT 1335.255 255.440 1335.770 255.580 ;
        RECT 1335.450 255.380 1335.770 255.440 ;
        RECT 1335.450 241.640 1335.770 241.700 ;
        RECT 1335.255 241.500 1335.770 241.640 ;
        RECT 1335.450 241.440 1335.770 241.500 ;
        RECT 1335.005 207.640 1335.295 207.685 ;
        RECT 1335.450 207.640 1335.770 207.700 ;
        RECT 1335.005 207.500 1335.770 207.640 ;
        RECT 1335.005 207.455 1335.295 207.500 ;
        RECT 1335.450 207.440 1335.770 207.500 ;
        RECT 1334.990 193.360 1335.310 193.420 ;
        RECT 1334.795 193.220 1335.310 193.360 ;
        RECT 1334.990 193.160 1335.310 193.220 ;
        RECT 1334.990 158.680 1335.310 158.740 ;
        RECT 1335.910 158.680 1336.230 158.740 ;
        RECT 1334.990 158.540 1336.230 158.680 ;
        RECT 1334.990 158.480 1335.310 158.540 ;
        RECT 1335.910 158.480 1336.230 158.540 ;
        RECT 1335.465 144.740 1335.755 144.785 ;
        RECT 1335.910 144.740 1336.230 144.800 ;
        RECT 1335.465 144.600 1336.230 144.740 ;
        RECT 1335.465 144.555 1335.755 144.600 ;
        RECT 1335.910 144.540 1336.230 144.600 ;
        RECT 1335.450 96.800 1335.770 96.860 ;
        RECT 1335.255 96.660 1335.770 96.800 ;
        RECT 1335.450 96.600 1335.770 96.660 ;
        RECT 1335.910 24.040 1336.230 24.100 ;
        RECT 1453.670 24.040 1453.990 24.100 ;
        RECT 1335.910 23.900 1453.990 24.040 ;
        RECT 1335.910 23.840 1336.230 23.900 ;
        RECT 1453.670 23.840 1453.990 23.900 ;
      LAYER via ;
        RECT 988.640 499.840 988.900 500.100 ;
        RECT 1335.020 499.840 1335.280 500.100 ;
        RECT 1335.020 482.840 1335.280 483.100 ;
        RECT 1335.020 448.160 1335.280 448.420 ;
        RECT 1335.480 400.560 1335.740 400.820 ;
        RECT 1335.480 386.280 1335.740 386.540 ;
        RECT 1335.480 351.940 1335.740 352.200 ;
        RECT 1335.480 338.000 1335.740 338.260 ;
        RECT 1335.480 313.520 1335.740 313.780 ;
        RECT 1335.480 289.720 1335.740 289.980 ;
        RECT 1335.480 255.380 1335.740 255.640 ;
        RECT 1335.480 241.440 1335.740 241.700 ;
        RECT 1335.480 207.440 1335.740 207.700 ;
        RECT 1335.020 193.160 1335.280 193.420 ;
        RECT 1335.020 158.480 1335.280 158.740 ;
        RECT 1335.940 158.480 1336.200 158.740 ;
        RECT 1335.940 144.540 1336.200 144.800 ;
        RECT 1335.480 96.600 1335.740 96.860 ;
        RECT 1335.940 23.840 1336.200 24.100 ;
        RECT 1453.700 23.840 1453.960 24.100 ;
      LAYER met2 ;
        RECT 988.770 510.340 989.050 514.000 ;
        RECT 988.700 510.000 989.050 510.340 ;
        RECT 988.700 500.130 988.840 510.000 ;
        RECT 988.640 499.810 988.900 500.130 ;
        RECT 1335.020 499.810 1335.280 500.130 ;
        RECT 1335.080 483.130 1335.220 499.810 ;
        RECT 1335.020 482.810 1335.280 483.130 ;
        RECT 1335.020 448.130 1335.280 448.450 ;
        RECT 1335.080 434.930 1335.220 448.130 ;
        RECT 1335.080 434.790 1335.680 434.930 ;
        RECT 1335.540 400.850 1335.680 434.790 ;
        RECT 1335.480 400.530 1335.740 400.850 ;
        RECT 1335.480 386.250 1335.740 386.570 ;
        RECT 1335.540 352.230 1335.680 386.250 ;
        RECT 1335.480 351.910 1335.740 352.230 ;
        RECT 1335.480 337.970 1335.740 338.290 ;
        RECT 1335.540 313.810 1335.680 337.970 ;
        RECT 1335.480 313.490 1335.740 313.810 ;
        RECT 1335.480 289.690 1335.740 290.010 ;
        RECT 1335.540 255.670 1335.680 289.690 ;
        RECT 1335.480 255.350 1335.740 255.670 ;
        RECT 1335.480 241.410 1335.740 241.730 ;
        RECT 1335.540 207.730 1335.680 241.410 ;
        RECT 1335.480 207.410 1335.740 207.730 ;
        RECT 1335.020 193.130 1335.280 193.450 ;
        RECT 1335.080 158.770 1335.220 193.130 ;
        RECT 1335.020 158.450 1335.280 158.770 ;
        RECT 1335.940 158.450 1336.200 158.770 ;
        RECT 1336.000 144.830 1336.140 158.450 ;
        RECT 1335.940 144.510 1336.200 144.830 ;
        RECT 1335.480 96.570 1335.740 96.890 ;
        RECT 1335.540 62.290 1335.680 96.570 ;
        RECT 1335.540 62.150 1336.140 62.290 ;
        RECT 1336.000 24.130 1336.140 62.150 ;
        RECT 1335.940 23.810 1336.200 24.130 ;
        RECT 1453.700 23.810 1453.960 24.130 ;
        RECT 1453.760 2.400 1453.900 23.810 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.030 498.680 1001.350 498.740 ;
        RECT 1007.010 498.680 1007.330 498.740 ;
        RECT 1001.030 498.540 1007.330 498.680 ;
        RECT 1001.030 498.480 1001.350 498.540 ;
        RECT 1007.010 498.480 1007.330 498.540 ;
        RECT 1007.010 86.260 1007.330 86.320 ;
        RECT 1469.770 86.260 1470.090 86.320 ;
        RECT 1007.010 86.120 1470.090 86.260 ;
        RECT 1007.010 86.060 1007.330 86.120 ;
        RECT 1469.770 86.060 1470.090 86.120 ;
      LAYER via ;
        RECT 1001.060 498.480 1001.320 498.740 ;
        RECT 1007.040 498.480 1007.300 498.740 ;
        RECT 1007.040 86.060 1007.300 86.320 ;
        RECT 1469.800 86.060 1470.060 86.320 ;
      LAYER met2 ;
        RECT 1001.190 510.340 1001.470 514.000 ;
        RECT 1001.120 510.000 1001.470 510.340 ;
        RECT 1001.120 498.770 1001.260 510.000 ;
        RECT 1001.060 498.450 1001.320 498.770 ;
        RECT 1007.040 498.450 1007.300 498.770 ;
        RECT 1007.100 86.350 1007.240 498.450 ;
        RECT 1007.040 86.030 1007.300 86.350 ;
        RECT 1469.800 86.030 1470.060 86.350 ;
        RECT 1469.860 17.410 1470.000 86.030 ;
        RECT 1469.860 17.270 1471.840 17.410 ;
        RECT 1471.700 2.400 1471.840 17.270 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1013.450 497.320 1013.770 497.380 ;
        RECT 1038.290 497.320 1038.610 497.380 ;
        RECT 1013.450 497.180 1038.610 497.320 ;
        RECT 1013.450 497.120 1013.770 497.180 ;
        RECT 1038.290 497.120 1038.610 497.180 ;
        RECT 1038.290 93.060 1038.610 93.120 ;
        RECT 1484.030 93.060 1484.350 93.120 ;
        RECT 1038.290 92.920 1484.350 93.060 ;
        RECT 1038.290 92.860 1038.610 92.920 ;
        RECT 1484.030 92.860 1484.350 92.920 ;
      LAYER via ;
        RECT 1013.480 497.120 1013.740 497.380 ;
        RECT 1038.320 497.120 1038.580 497.380 ;
        RECT 1038.320 92.860 1038.580 93.120 ;
        RECT 1484.060 92.860 1484.320 93.120 ;
      LAYER met2 ;
        RECT 1013.610 510.340 1013.890 514.000 ;
        RECT 1013.540 510.000 1013.890 510.340 ;
        RECT 1013.540 497.410 1013.680 510.000 ;
        RECT 1013.480 497.090 1013.740 497.410 ;
        RECT 1038.320 497.090 1038.580 497.410 ;
        RECT 1038.380 93.150 1038.520 497.090 ;
        RECT 1038.320 92.830 1038.580 93.150 ;
        RECT 1484.060 92.830 1484.320 93.150 ;
        RECT 1484.120 16.730 1484.260 92.830 ;
        RECT 1484.120 16.590 1489.780 16.730 ;
        RECT 1489.640 2.400 1489.780 16.590 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 99.860 1028.030 99.920 ;
        RECT 1504.270 99.860 1504.590 99.920 ;
        RECT 1027.710 99.720 1504.590 99.860 ;
        RECT 1027.710 99.660 1028.030 99.720 ;
        RECT 1504.270 99.660 1504.590 99.720 ;
      LAYER via ;
        RECT 1027.740 99.660 1028.000 99.920 ;
        RECT 1504.300 99.660 1504.560 99.920 ;
      LAYER met2 ;
        RECT 1026.030 510.410 1026.310 514.000 ;
        RECT 1026.030 510.270 1027.940 510.410 ;
        RECT 1026.030 510.000 1026.310 510.270 ;
        RECT 1027.800 99.950 1027.940 510.270 ;
        RECT 1027.740 99.630 1028.000 99.950 ;
        RECT 1504.300 99.630 1504.560 99.950 ;
        RECT 1504.360 16.730 1504.500 99.630 ;
        RECT 1504.360 16.590 1507.260 16.730 ;
        RECT 1507.120 2.400 1507.260 16.590 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 469.270 503.100 469.590 503.160 ;
        RECT 486.290 503.100 486.610 503.160 ;
        RECT 469.270 502.960 486.610 503.100 ;
        RECT 469.270 502.900 469.590 502.960 ;
        RECT 486.290 502.900 486.610 502.960 ;
        RECT 486.290 99.860 486.610 99.920 ;
        RECT 704.330 99.860 704.650 99.920 ;
        RECT 486.290 99.720 704.650 99.860 ;
        RECT 486.290 99.660 486.610 99.720 ;
        RECT 704.330 99.660 704.650 99.720 ;
      LAYER via ;
        RECT 469.300 502.900 469.560 503.160 ;
        RECT 486.320 502.900 486.580 503.160 ;
        RECT 486.320 99.660 486.580 99.920 ;
        RECT 704.360 99.660 704.620 99.920 ;
      LAYER met2 ;
        RECT 469.430 510.340 469.710 514.000 ;
        RECT 469.360 510.000 469.710 510.340 ;
        RECT 469.360 503.190 469.500 510.000 ;
        RECT 469.300 502.870 469.560 503.190 ;
        RECT 486.320 502.870 486.580 503.190 ;
        RECT 486.380 99.950 486.520 502.870 ;
        RECT 486.320 99.630 486.580 99.950 ;
        RECT 704.360 99.630 704.620 99.950 ;
        RECT 704.420 2.400 704.560 99.630 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 107.340 1041.830 107.400 ;
        RECT 1525.430 107.340 1525.750 107.400 ;
        RECT 1041.510 107.200 1525.750 107.340 ;
        RECT 1041.510 107.140 1041.830 107.200 ;
        RECT 1525.430 107.140 1525.750 107.200 ;
      LAYER via ;
        RECT 1041.540 107.140 1041.800 107.400 ;
        RECT 1525.460 107.140 1525.720 107.400 ;
      LAYER met2 ;
        RECT 1038.450 510.410 1038.730 514.000 ;
        RECT 1038.450 510.270 1041.740 510.410 ;
        RECT 1038.450 510.000 1038.730 510.270 ;
        RECT 1041.600 107.430 1041.740 510.270 ;
        RECT 1041.540 107.110 1041.800 107.430 ;
        RECT 1525.460 107.110 1525.720 107.430 ;
        RECT 1525.520 17.410 1525.660 107.110 ;
        RECT 1525.060 17.270 1525.660 17.410 ;
        RECT 1525.060 2.400 1525.200 17.270 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1050.710 496.980 1051.030 497.040 ;
        RECT 1054.850 496.980 1055.170 497.040 ;
        RECT 1050.710 496.840 1055.170 496.980 ;
        RECT 1050.710 496.780 1051.030 496.840 ;
        RECT 1054.850 496.780 1055.170 496.840 ;
        RECT 1054.850 444.960 1055.170 445.020 ;
        RECT 1538.770 444.960 1539.090 445.020 ;
        RECT 1054.850 444.820 1539.090 444.960 ;
        RECT 1054.850 444.760 1055.170 444.820 ;
        RECT 1538.770 444.760 1539.090 444.820 ;
        RECT 1538.770 2.960 1539.090 3.020 ;
        RECT 1542.910 2.960 1543.230 3.020 ;
        RECT 1538.770 2.820 1543.230 2.960 ;
        RECT 1538.770 2.760 1539.090 2.820 ;
        RECT 1542.910 2.760 1543.230 2.820 ;
      LAYER via ;
        RECT 1050.740 496.780 1051.000 497.040 ;
        RECT 1054.880 496.780 1055.140 497.040 ;
        RECT 1054.880 444.760 1055.140 445.020 ;
        RECT 1538.800 444.760 1539.060 445.020 ;
        RECT 1538.800 2.760 1539.060 3.020 ;
        RECT 1542.940 2.760 1543.200 3.020 ;
      LAYER met2 ;
        RECT 1050.870 510.340 1051.150 514.000 ;
        RECT 1050.800 510.000 1051.150 510.340 ;
        RECT 1050.800 497.070 1050.940 510.000 ;
        RECT 1050.740 496.750 1051.000 497.070 ;
        RECT 1054.880 496.750 1055.140 497.070 ;
        RECT 1054.940 445.050 1055.080 496.750 ;
        RECT 1054.880 444.730 1055.140 445.050 ;
        RECT 1538.800 444.730 1539.060 445.050 ;
        RECT 1538.860 3.050 1539.000 444.730 ;
        RECT 1538.800 2.730 1539.060 3.050 ;
        RECT 1542.940 2.730 1543.200 3.050 ;
        RECT 1543.000 2.400 1543.140 2.730 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1063.130 496.980 1063.450 497.040 ;
        RECT 1069.110 496.980 1069.430 497.040 ;
        RECT 1063.130 496.840 1069.430 496.980 ;
        RECT 1063.130 496.780 1063.450 496.840 ;
        RECT 1069.110 496.780 1069.430 496.840 ;
        RECT 1069.110 182.820 1069.430 182.880 ;
        RECT 1559.470 182.820 1559.790 182.880 ;
        RECT 1069.110 182.680 1559.790 182.820 ;
        RECT 1069.110 182.620 1069.430 182.680 ;
        RECT 1559.470 182.620 1559.790 182.680 ;
      LAYER via ;
        RECT 1063.160 496.780 1063.420 497.040 ;
        RECT 1069.140 496.780 1069.400 497.040 ;
        RECT 1069.140 182.620 1069.400 182.880 ;
        RECT 1559.500 182.620 1559.760 182.880 ;
      LAYER met2 ;
        RECT 1063.290 510.340 1063.570 514.000 ;
        RECT 1063.220 510.000 1063.570 510.340 ;
        RECT 1063.220 497.070 1063.360 510.000 ;
        RECT 1063.160 496.750 1063.420 497.070 ;
        RECT 1069.140 496.750 1069.400 497.070 ;
        RECT 1069.200 182.910 1069.340 496.750 ;
        RECT 1069.140 182.590 1069.400 182.910 ;
        RECT 1559.500 182.590 1559.760 182.910 ;
        RECT 1559.560 3.130 1559.700 182.590 ;
        RECT 1559.560 2.990 1561.080 3.130 ;
        RECT 1560.940 2.400 1561.080 2.990 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1075.165 138.125 1075.335 186.235 ;
      LAYER mcon ;
        RECT 1075.165 186.065 1075.335 186.235 ;
      LAYER met1 ;
        RECT 1075.090 372.540 1075.410 372.600 ;
        RECT 1076.010 372.540 1076.330 372.600 ;
        RECT 1075.090 372.400 1076.330 372.540 ;
        RECT 1075.090 372.340 1075.410 372.400 ;
        RECT 1076.010 372.340 1076.330 372.400 ;
        RECT 1074.630 317.460 1074.950 317.520 ;
        RECT 1075.090 317.460 1075.410 317.520 ;
        RECT 1074.630 317.320 1075.410 317.460 ;
        RECT 1074.630 317.260 1074.950 317.320 ;
        RECT 1075.090 317.260 1075.410 317.320 ;
        RECT 1074.630 207.100 1074.950 207.360 ;
        RECT 1074.720 206.620 1074.860 207.100 ;
        RECT 1075.090 206.620 1075.410 206.680 ;
        RECT 1074.720 206.480 1075.410 206.620 ;
        RECT 1075.090 206.420 1075.410 206.480 ;
        RECT 1075.090 186.220 1075.410 186.280 ;
        RECT 1074.895 186.080 1075.410 186.220 ;
        RECT 1075.090 186.020 1075.410 186.080 ;
        RECT 1075.105 138.280 1075.395 138.325 ;
        RECT 1075.550 138.280 1075.870 138.340 ;
        RECT 1075.105 138.140 1075.870 138.280 ;
        RECT 1075.105 138.095 1075.395 138.140 ;
        RECT 1075.550 138.080 1075.870 138.140 ;
        RECT 1075.550 114.140 1075.870 114.200 ;
        RECT 1573.270 114.140 1573.590 114.200 ;
        RECT 1075.550 114.000 1573.590 114.140 ;
        RECT 1075.550 113.940 1075.870 114.000 ;
        RECT 1573.270 113.940 1573.590 114.000 ;
        RECT 1573.270 2.960 1573.590 3.020 ;
        RECT 1578.790 2.960 1579.110 3.020 ;
        RECT 1573.270 2.820 1579.110 2.960 ;
        RECT 1573.270 2.760 1573.590 2.820 ;
        RECT 1578.790 2.760 1579.110 2.820 ;
      LAYER via ;
        RECT 1075.120 372.340 1075.380 372.600 ;
        RECT 1076.040 372.340 1076.300 372.600 ;
        RECT 1074.660 317.260 1074.920 317.520 ;
        RECT 1075.120 317.260 1075.380 317.520 ;
        RECT 1074.660 207.100 1074.920 207.360 ;
        RECT 1075.120 206.420 1075.380 206.680 ;
        RECT 1075.120 186.020 1075.380 186.280 ;
        RECT 1075.580 138.080 1075.840 138.340 ;
        RECT 1075.580 113.940 1075.840 114.200 ;
        RECT 1573.300 113.940 1573.560 114.200 ;
        RECT 1573.300 2.760 1573.560 3.020 ;
        RECT 1578.820 2.760 1579.080 3.020 ;
      LAYER met2 ;
        RECT 1075.710 510.340 1075.990 514.000 ;
        RECT 1075.640 510.000 1075.990 510.340 ;
        RECT 1075.640 468.930 1075.780 510.000 ;
        RECT 1075.640 468.790 1076.240 468.930 ;
        RECT 1076.100 400.250 1076.240 468.790 ;
        RECT 1075.180 400.110 1076.240 400.250 ;
        RECT 1075.180 372.630 1075.320 400.110 ;
        RECT 1075.120 372.310 1075.380 372.630 ;
        RECT 1076.040 372.310 1076.300 372.630 ;
        RECT 1076.100 324.885 1076.240 372.310 ;
        RECT 1075.110 324.770 1075.390 324.885 ;
        RECT 1074.720 324.630 1075.390 324.770 ;
        RECT 1074.720 317.550 1074.860 324.630 ;
        RECT 1075.110 324.515 1075.390 324.630 ;
        RECT 1076.030 324.515 1076.310 324.885 ;
        RECT 1074.660 317.230 1074.920 317.550 ;
        RECT 1075.120 317.230 1075.380 317.550 ;
        RECT 1075.180 303.805 1075.320 317.230 ;
        RECT 1075.110 303.435 1075.390 303.805 ;
        RECT 1075.110 241.810 1075.390 241.925 ;
        RECT 1074.720 241.670 1075.390 241.810 ;
        RECT 1074.720 207.390 1074.860 241.670 ;
        RECT 1075.110 241.555 1075.390 241.670 ;
        RECT 1074.660 207.070 1074.920 207.390 ;
        RECT 1075.120 206.390 1075.380 206.710 ;
        RECT 1075.180 186.310 1075.320 206.390 ;
        RECT 1075.120 185.990 1075.380 186.310 ;
        RECT 1075.580 138.050 1075.840 138.370 ;
        RECT 1075.640 114.230 1075.780 138.050 ;
        RECT 1075.580 113.910 1075.840 114.230 ;
        RECT 1573.300 113.910 1573.560 114.230 ;
        RECT 1573.360 3.050 1573.500 113.910 ;
        RECT 1573.300 2.730 1573.560 3.050 ;
        RECT 1578.820 2.730 1579.080 3.050 ;
        RECT 1578.880 2.400 1579.020 2.730 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
      LAYER via2 ;
        RECT 1075.110 324.560 1075.390 324.840 ;
        RECT 1076.030 324.560 1076.310 324.840 ;
        RECT 1075.110 303.480 1075.390 303.760 ;
        RECT 1075.110 241.600 1075.390 241.880 ;
      LAYER met3 ;
        RECT 1075.085 324.850 1075.415 324.865 ;
        RECT 1076.005 324.850 1076.335 324.865 ;
        RECT 1075.085 324.550 1076.335 324.850 ;
        RECT 1075.085 324.535 1075.415 324.550 ;
        RECT 1076.005 324.535 1076.335 324.550 ;
        RECT 1075.085 303.770 1075.415 303.785 ;
        RECT 1075.750 303.770 1076.130 303.780 ;
        RECT 1075.085 303.470 1076.130 303.770 ;
        RECT 1075.085 303.455 1075.415 303.470 ;
        RECT 1075.750 303.460 1076.130 303.470 ;
        RECT 1075.085 241.890 1075.415 241.905 ;
        RECT 1075.750 241.890 1076.130 241.900 ;
        RECT 1075.085 241.590 1076.130 241.890 ;
        RECT 1075.085 241.575 1075.415 241.590 ;
        RECT 1075.750 241.580 1076.130 241.590 ;
      LAYER via3 ;
        RECT 1075.780 303.460 1076.100 303.780 ;
        RECT 1075.780 241.580 1076.100 241.900 ;
      LAYER met4 ;
        RECT 1075.775 303.455 1076.105 303.785 ;
        RECT 1075.790 241.905 1076.090 303.455 ;
        RECT 1075.775 241.575 1076.105 241.905 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1087.970 500.720 1088.290 500.780 ;
        RECT 1121.090 500.720 1121.410 500.780 ;
        RECT 1087.970 500.580 1121.410 500.720 ;
        RECT 1087.970 500.520 1088.290 500.580 ;
        RECT 1121.090 500.520 1121.410 500.580 ;
        RECT 1121.090 120.940 1121.410 121.000 ;
        RECT 1593.970 120.940 1594.290 121.000 ;
        RECT 1121.090 120.800 1594.290 120.940 ;
        RECT 1121.090 120.740 1121.410 120.800 ;
        RECT 1593.970 120.740 1594.290 120.800 ;
      LAYER via ;
        RECT 1088.000 500.520 1088.260 500.780 ;
        RECT 1121.120 500.520 1121.380 500.780 ;
        RECT 1121.120 120.740 1121.380 121.000 ;
        RECT 1594.000 120.740 1594.260 121.000 ;
      LAYER met2 ;
        RECT 1088.130 510.340 1088.410 514.000 ;
        RECT 1088.060 510.000 1088.410 510.340 ;
        RECT 1088.060 500.810 1088.200 510.000 ;
        RECT 1088.000 500.490 1088.260 500.810 ;
        RECT 1121.120 500.490 1121.380 500.810 ;
        RECT 1121.180 121.030 1121.320 500.490 ;
        RECT 1121.120 120.710 1121.380 121.030 ;
        RECT 1594.000 120.710 1594.260 121.030 ;
        RECT 1594.060 16.730 1594.200 120.710 ;
        RECT 1594.060 16.590 1596.500 16.730 ;
        RECT 1596.360 2.400 1596.500 16.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1103.610 189.960 1103.930 190.020 ;
        RECT 1608.230 189.960 1608.550 190.020 ;
        RECT 1103.610 189.820 1608.550 189.960 ;
        RECT 1103.610 189.760 1103.930 189.820 ;
        RECT 1608.230 189.760 1608.550 189.820 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1608.230 17.780 1614.530 17.920 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
      LAYER via ;
        RECT 1103.640 189.760 1103.900 190.020 ;
        RECT 1608.260 189.760 1608.520 190.020 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
      LAYER met2 ;
        RECT 1100.090 510.410 1100.370 514.000 ;
        RECT 1100.090 510.270 1103.840 510.410 ;
        RECT 1100.090 510.000 1100.370 510.270 ;
        RECT 1103.700 190.050 1103.840 510.270 ;
        RECT 1103.640 189.730 1103.900 190.050 ;
        RECT 1608.260 189.730 1608.520 190.050 ;
        RECT 1608.320 18.010 1608.460 189.730 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1614.300 2.400 1614.440 17.690 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1112.350 496.980 1112.670 497.040 ;
        RECT 1116.950 496.980 1117.270 497.040 ;
        RECT 1112.350 496.840 1117.270 496.980 ;
        RECT 1112.350 496.780 1112.670 496.840 ;
        RECT 1116.950 496.780 1117.270 496.840 ;
        RECT 1116.950 196.760 1117.270 196.820 ;
        RECT 1628.470 196.760 1628.790 196.820 ;
        RECT 1116.950 196.620 1628.790 196.760 ;
        RECT 1116.950 196.560 1117.270 196.620 ;
        RECT 1628.470 196.560 1628.790 196.620 ;
      LAYER via ;
        RECT 1112.380 496.780 1112.640 497.040 ;
        RECT 1116.980 496.780 1117.240 497.040 ;
        RECT 1116.980 196.560 1117.240 196.820 ;
        RECT 1628.500 196.560 1628.760 196.820 ;
      LAYER met2 ;
        RECT 1112.510 510.340 1112.790 514.000 ;
        RECT 1112.440 510.000 1112.790 510.340 ;
        RECT 1112.440 497.070 1112.580 510.000 ;
        RECT 1112.380 496.750 1112.640 497.070 ;
        RECT 1116.980 496.750 1117.240 497.070 ;
        RECT 1117.040 196.850 1117.180 496.750 ;
        RECT 1116.980 196.530 1117.240 196.850 ;
        RECT 1628.500 196.530 1628.760 196.850 ;
        RECT 1628.560 17.410 1628.700 196.530 ;
        RECT 1628.560 17.270 1632.380 17.410 ;
        RECT 1632.240 2.400 1632.380 17.270 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1124.770 496.980 1125.090 497.040 ;
        RECT 1131.210 496.980 1131.530 497.040 ;
        RECT 1124.770 496.840 1131.530 496.980 ;
        RECT 1124.770 496.780 1125.090 496.840 ;
        RECT 1131.210 496.780 1131.530 496.840 ;
        RECT 1131.210 204.240 1131.530 204.300 ;
        RECT 1649.170 204.240 1649.490 204.300 ;
        RECT 1131.210 204.100 1649.490 204.240 ;
        RECT 1131.210 204.040 1131.530 204.100 ;
        RECT 1649.170 204.040 1649.490 204.100 ;
      LAYER via ;
        RECT 1124.800 496.780 1125.060 497.040 ;
        RECT 1131.240 496.780 1131.500 497.040 ;
        RECT 1131.240 204.040 1131.500 204.300 ;
        RECT 1649.200 204.040 1649.460 204.300 ;
      LAYER met2 ;
        RECT 1124.930 510.340 1125.210 514.000 ;
        RECT 1124.860 510.000 1125.210 510.340 ;
        RECT 1124.860 497.070 1125.000 510.000 ;
        RECT 1124.800 496.750 1125.060 497.070 ;
        RECT 1131.240 496.750 1131.500 497.070 ;
        RECT 1131.300 204.330 1131.440 496.750 ;
        RECT 1131.240 204.010 1131.500 204.330 ;
        RECT 1649.200 204.010 1649.460 204.330 ;
        RECT 1649.260 17.410 1649.400 204.010 ;
        RECT 1649.260 17.270 1650.320 17.410 ;
        RECT 1650.180 2.400 1650.320 17.270 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1137.265 434.945 1137.435 448.715 ;
        RECT 1136.805 138.125 1136.975 186.235 ;
      LAYER mcon ;
        RECT 1137.265 448.545 1137.435 448.715 ;
        RECT 1136.805 186.065 1136.975 186.235 ;
      LAYER met1 ;
        RECT 1137.190 448.700 1137.510 448.760 ;
        RECT 1136.995 448.560 1137.510 448.700 ;
        RECT 1137.190 448.500 1137.510 448.560 ;
        RECT 1137.190 435.100 1137.510 435.160 ;
        RECT 1136.995 434.960 1137.510 435.100 ;
        RECT 1137.190 434.900 1137.510 434.960 ;
        RECT 1135.350 410.280 1135.670 410.340 ;
        RECT 1137.190 410.280 1137.510 410.340 ;
        RECT 1135.350 410.140 1137.510 410.280 ;
        RECT 1135.350 410.080 1135.670 410.140 ;
        RECT 1137.190 410.080 1137.510 410.140 ;
        RECT 1136.730 352.480 1137.050 352.540 ;
        RECT 1136.360 352.340 1137.050 352.480 ;
        RECT 1136.360 351.860 1136.500 352.340 ;
        RECT 1136.730 352.280 1137.050 352.340 ;
        RECT 1136.270 351.600 1136.590 351.860 ;
        RECT 1136.270 331.060 1136.590 331.120 ;
        RECT 1137.190 331.060 1137.510 331.120 ;
        RECT 1136.270 330.920 1137.510 331.060 ;
        RECT 1136.270 330.860 1136.590 330.920 ;
        RECT 1137.190 330.860 1137.510 330.920 ;
        RECT 1136.270 207.100 1136.590 207.360 ;
        RECT 1136.360 206.620 1136.500 207.100 ;
        RECT 1136.730 206.620 1137.050 206.680 ;
        RECT 1136.360 206.480 1137.050 206.620 ;
        RECT 1136.730 206.420 1137.050 206.480 ;
        RECT 1136.730 186.220 1137.050 186.280 ;
        RECT 1136.535 186.080 1137.050 186.220 ;
        RECT 1136.730 186.020 1137.050 186.080 ;
        RECT 1136.745 138.280 1137.035 138.325 ;
        RECT 1137.190 138.280 1137.510 138.340 ;
        RECT 1136.745 138.140 1137.510 138.280 ;
        RECT 1136.745 138.095 1137.035 138.140 ;
        RECT 1137.190 138.080 1137.510 138.140 ;
        RECT 1137.190 127.740 1137.510 127.800 ;
        RECT 1662.970 127.740 1663.290 127.800 ;
        RECT 1137.190 127.600 1663.290 127.740 ;
        RECT 1137.190 127.540 1137.510 127.600 ;
        RECT 1662.970 127.540 1663.290 127.600 ;
      LAYER via ;
        RECT 1137.220 448.500 1137.480 448.760 ;
        RECT 1137.220 434.900 1137.480 435.160 ;
        RECT 1135.380 410.080 1135.640 410.340 ;
        RECT 1137.220 410.080 1137.480 410.340 ;
        RECT 1136.760 352.280 1137.020 352.540 ;
        RECT 1136.300 351.600 1136.560 351.860 ;
        RECT 1136.300 330.860 1136.560 331.120 ;
        RECT 1137.220 330.860 1137.480 331.120 ;
        RECT 1136.300 207.100 1136.560 207.360 ;
        RECT 1136.760 206.420 1137.020 206.680 ;
        RECT 1136.760 186.020 1137.020 186.280 ;
        RECT 1137.220 138.080 1137.480 138.340 ;
        RECT 1137.220 127.540 1137.480 127.800 ;
        RECT 1663.000 127.540 1663.260 127.800 ;
      LAYER met2 ;
        RECT 1137.350 510.340 1137.630 514.000 ;
        RECT 1137.280 510.000 1137.630 510.340 ;
        RECT 1137.280 448.790 1137.420 510.000 ;
        RECT 1137.220 448.470 1137.480 448.790 ;
        RECT 1137.220 434.870 1137.480 435.190 ;
        RECT 1137.280 410.370 1137.420 434.870 ;
        RECT 1135.380 410.050 1135.640 410.370 ;
        RECT 1137.220 410.050 1137.480 410.370 ;
        RECT 1135.440 386.765 1135.580 410.050 ;
        RECT 1135.370 386.395 1135.650 386.765 ;
        RECT 1136.290 386.650 1136.570 386.765 ;
        RECT 1136.290 386.510 1136.960 386.650 ;
        RECT 1136.290 386.395 1136.570 386.510 ;
        RECT 1136.820 352.570 1136.960 386.510 ;
        RECT 1136.760 352.250 1137.020 352.570 ;
        RECT 1136.300 351.570 1136.560 351.890 ;
        RECT 1136.360 339.165 1136.500 351.570 ;
        RECT 1136.290 338.795 1136.570 339.165 ;
        RECT 1136.290 338.115 1136.570 338.485 ;
        RECT 1136.360 331.150 1136.500 338.115 ;
        RECT 1136.300 330.830 1136.560 331.150 ;
        RECT 1137.220 330.830 1137.480 331.150 ;
        RECT 1137.280 307.205 1137.420 330.830 ;
        RECT 1137.210 306.835 1137.490 307.205 ;
        RECT 1136.750 241.810 1137.030 241.925 ;
        RECT 1136.360 241.670 1137.030 241.810 ;
        RECT 1136.360 207.390 1136.500 241.670 ;
        RECT 1136.750 241.555 1137.030 241.670 ;
        RECT 1136.300 207.070 1136.560 207.390 ;
        RECT 1136.760 206.390 1137.020 206.710 ;
        RECT 1136.820 186.310 1136.960 206.390 ;
        RECT 1136.760 185.990 1137.020 186.310 ;
        RECT 1137.220 138.050 1137.480 138.370 ;
        RECT 1137.280 127.830 1137.420 138.050 ;
        RECT 1137.220 127.510 1137.480 127.830 ;
        RECT 1663.000 127.510 1663.260 127.830 ;
        RECT 1663.060 17.410 1663.200 127.510 ;
        RECT 1663.060 17.270 1668.260 17.410 ;
        RECT 1668.120 2.400 1668.260 17.270 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
      LAYER via2 ;
        RECT 1135.370 386.440 1135.650 386.720 ;
        RECT 1136.290 386.440 1136.570 386.720 ;
        RECT 1136.290 338.840 1136.570 339.120 ;
        RECT 1136.290 338.160 1136.570 338.440 ;
        RECT 1137.210 306.880 1137.490 307.160 ;
        RECT 1136.750 241.600 1137.030 241.880 ;
      LAYER met3 ;
        RECT 1135.345 386.730 1135.675 386.745 ;
        RECT 1136.265 386.730 1136.595 386.745 ;
        RECT 1135.345 386.430 1136.595 386.730 ;
        RECT 1135.345 386.415 1135.675 386.430 ;
        RECT 1136.265 386.415 1136.595 386.430 ;
        RECT 1136.265 338.815 1136.595 339.145 ;
        RECT 1136.280 338.465 1136.580 338.815 ;
        RECT 1136.265 338.135 1136.595 338.465 ;
        RECT 1137.185 307.180 1137.515 307.185 ;
        RECT 1137.185 307.170 1137.770 307.180 ;
        RECT 1136.960 306.870 1137.770 307.170 ;
        RECT 1137.185 306.860 1137.770 306.870 ;
        RECT 1137.185 306.855 1137.515 306.860 ;
        RECT 1136.725 241.890 1137.055 241.905 ;
        RECT 1137.390 241.890 1137.770 241.900 ;
        RECT 1136.725 241.590 1137.770 241.890 ;
        RECT 1136.725 241.575 1137.055 241.590 ;
        RECT 1137.390 241.580 1137.770 241.590 ;
      LAYER via3 ;
        RECT 1137.420 306.860 1137.740 307.180 ;
        RECT 1137.420 241.580 1137.740 241.900 ;
      LAYER met4 ;
        RECT 1137.415 306.855 1137.745 307.185 ;
        RECT 1137.430 241.905 1137.730 306.855 ;
        RECT 1137.415 241.575 1137.745 241.905 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 134.540 1152.230 134.600 ;
        RECT 1683.670 134.540 1683.990 134.600 ;
        RECT 1151.910 134.400 1683.990 134.540 ;
        RECT 1151.910 134.340 1152.230 134.400 ;
        RECT 1683.670 134.340 1683.990 134.400 ;
      LAYER via ;
        RECT 1151.940 134.340 1152.200 134.600 ;
        RECT 1683.700 134.340 1683.960 134.600 ;
      LAYER met2 ;
        RECT 1149.770 510.410 1150.050 514.000 ;
        RECT 1149.770 510.270 1152.140 510.410 ;
        RECT 1149.770 510.000 1150.050 510.270 ;
        RECT 1152.000 134.630 1152.140 510.270 ;
        RECT 1151.940 134.310 1152.200 134.630 ;
        RECT 1683.700 134.310 1683.960 134.630 ;
        RECT 1683.760 17.410 1683.900 134.310 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 481.305 282.965 481.475 331.075 ;
        RECT 481.305 234.685 481.475 282.455 ;
      LAYER mcon ;
        RECT 481.305 330.905 481.475 331.075 ;
        RECT 481.305 282.285 481.475 282.455 ;
      LAYER met1 ;
        RECT 481.690 427.960 482.010 428.020 ;
        RECT 482.150 427.960 482.470 428.020 ;
        RECT 481.690 427.820 482.470 427.960 ;
        RECT 481.690 427.760 482.010 427.820 ;
        RECT 482.150 427.760 482.470 427.820 ;
        RECT 481.245 331.060 481.535 331.105 ;
        RECT 481.690 331.060 482.010 331.120 ;
        RECT 481.245 330.920 482.010 331.060 ;
        RECT 481.245 330.875 481.535 330.920 ;
        RECT 481.690 330.860 482.010 330.920 ;
        RECT 481.230 283.120 481.550 283.180 ;
        RECT 481.035 282.980 481.550 283.120 ;
        RECT 481.230 282.920 481.550 282.980 ;
        RECT 481.230 282.440 481.550 282.500 ;
        RECT 481.035 282.300 481.550 282.440 ;
        RECT 481.230 282.240 481.550 282.300 ;
        RECT 481.245 234.840 481.535 234.885 ;
        RECT 481.690 234.840 482.010 234.900 ;
        RECT 481.245 234.700 482.010 234.840 ;
        RECT 481.245 234.655 481.535 234.700 ;
        RECT 481.690 234.640 482.010 234.700 ;
        RECT 481.690 207.300 482.010 207.360 ;
        RECT 481.320 207.160 482.010 207.300 ;
        RECT 481.320 207.020 481.460 207.160 ;
        RECT 481.690 207.100 482.010 207.160 ;
        RECT 481.230 206.760 481.550 207.020 ;
        RECT 481.230 159.020 481.550 159.080 ;
        RECT 480.860 158.880 481.550 159.020 ;
        RECT 480.860 158.740 481.000 158.880 ;
        RECT 481.230 158.820 481.550 158.880 ;
        RECT 480.770 158.480 481.090 158.740 ;
        RECT 480.770 113.800 481.090 113.860 ;
        RECT 717.670 113.800 717.990 113.860 ;
        RECT 480.770 113.660 717.990 113.800 ;
        RECT 480.770 113.600 481.090 113.660 ;
        RECT 717.670 113.600 717.990 113.660 ;
        RECT 717.670 62.120 717.990 62.180 ;
        RECT 722.270 62.120 722.590 62.180 ;
        RECT 717.670 61.980 722.590 62.120 ;
        RECT 717.670 61.920 717.990 61.980 ;
        RECT 722.270 61.920 722.590 61.980 ;
      LAYER via ;
        RECT 481.720 427.760 481.980 428.020 ;
        RECT 482.180 427.760 482.440 428.020 ;
        RECT 481.720 330.860 481.980 331.120 ;
        RECT 481.260 282.920 481.520 283.180 ;
        RECT 481.260 282.240 481.520 282.500 ;
        RECT 481.720 234.640 481.980 234.900 ;
        RECT 481.720 207.100 481.980 207.360 ;
        RECT 481.260 206.760 481.520 207.020 ;
        RECT 481.260 158.820 481.520 159.080 ;
        RECT 480.800 158.480 481.060 158.740 ;
        RECT 480.800 113.600 481.060 113.860 ;
        RECT 717.700 113.600 717.960 113.860 ;
        RECT 717.700 61.920 717.960 62.180 ;
        RECT 722.300 61.920 722.560 62.180 ;
      LAYER met2 ;
        RECT 481.850 510.410 482.130 514.000 ;
        RECT 481.320 510.270 482.130 510.410 ;
        RECT 481.320 483.325 481.460 510.270 ;
        RECT 481.850 510.000 482.130 510.270 ;
        RECT 481.250 482.955 481.530 483.325 ;
        RECT 482.170 482.955 482.450 483.325 ;
        RECT 482.240 428.050 482.380 482.955 ;
        RECT 481.720 427.730 481.980 428.050 ;
        RECT 482.180 427.730 482.440 428.050 ;
        RECT 481.780 403.765 481.920 427.730 ;
        RECT 481.710 403.395 481.990 403.765 ;
        RECT 481.710 338.115 481.990 338.485 ;
        RECT 481.780 331.150 481.920 338.115 ;
        RECT 481.720 330.830 481.980 331.150 ;
        RECT 481.260 282.890 481.520 283.210 ;
        RECT 481.320 282.530 481.460 282.890 ;
        RECT 481.260 282.210 481.520 282.530 ;
        RECT 481.720 234.610 481.980 234.930 ;
        RECT 481.780 207.390 481.920 234.610 ;
        RECT 481.720 207.070 481.980 207.390 ;
        RECT 481.260 206.730 481.520 207.050 ;
        RECT 481.320 159.110 481.460 206.730 ;
        RECT 481.260 158.790 481.520 159.110 ;
        RECT 480.800 158.450 481.060 158.770 ;
        RECT 480.860 113.890 481.000 158.450 ;
        RECT 480.800 113.570 481.060 113.890 ;
        RECT 717.700 113.570 717.960 113.890 ;
        RECT 717.760 62.210 717.900 113.570 ;
        RECT 717.700 61.890 717.960 62.210 ;
        RECT 722.300 61.890 722.560 62.210 ;
        RECT 722.360 2.400 722.500 61.890 ;
        RECT 722.150 -4.800 722.710 2.400 ;
      LAYER via2 ;
        RECT 481.250 483.000 481.530 483.280 ;
        RECT 482.170 483.000 482.450 483.280 ;
        RECT 481.710 403.440 481.990 403.720 ;
        RECT 481.710 338.160 481.990 338.440 ;
      LAYER met3 ;
        RECT 481.225 483.290 481.555 483.305 ;
        RECT 482.145 483.290 482.475 483.305 ;
        RECT 481.225 482.990 482.475 483.290 ;
        RECT 481.225 482.975 481.555 482.990 ;
        RECT 482.145 482.975 482.475 482.990 ;
        RECT 481.685 403.740 482.015 403.745 ;
        RECT 481.430 403.730 482.015 403.740 ;
        RECT 481.230 403.430 482.015 403.730 ;
        RECT 481.430 403.420 482.015 403.430 ;
        RECT 481.685 403.415 482.015 403.420 ;
        RECT 481.430 339.130 481.810 339.140 ;
        RECT 481.430 338.830 482.690 339.130 ;
        RECT 481.430 338.820 481.810 338.830 ;
        RECT 481.685 338.450 482.015 338.465 ;
        RECT 482.390 338.450 482.690 338.830 ;
        RECT 481.685 338.150 482.690 338.450 ;
        RECT 481.685 338.135 482.015 338.150 ;
      LAYER via3 ;
        RECT 481.460 403.420 481.780 403.740 ;
        RECT 481.460 338.820 481.780 339.140 ;
      LAYER met4 ;
        RECT 481.455 403.415 481.785 403.745 ;
        RECT 481.470 339.145 481.770 403.415 ;
        RECT 481.455 338.815 481.785 339.145 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.030 496.980 1162.350 497.040 ;
        RECT 1165.710 496.980 1166.030 497.040 ;
        RECT 1162.030 496.840 1166.030 496.980 ;
        RECT 1162.030 496.780 1162.350 496.840 ;
        RECT 1165.710 496.780 1166.030 496.840 ;
        RECT 1165.710 30.840 1166.030 30.900 ;
        RECT 1703.450 30.840 1703.770 30.900 ;
        RECT 1165.710 30.700 1703.770 30.840 ;
        RECT 1165.710 30.640 1166.030 30.700 ;
        RECT 1703.450 30.640 1703.770 30.700 ;
      LAYER via ;
        RECT 1162.060 496.780 1162.320 497.040 ;
        RECT 1165.740 496.780 1166.000 497.040 ;
        RECT 1165.740 30.640 1166.000 30.900 ;
        RECT 1703.480 30.640 1703.740 30.900 ;
      LAYER met2 ;
        RECT 1162.190 510.340 1162.470 514.000 ;
        RECT 1162.120 510.000 1162.470 510.340 ;
        RECT 1162.120 497.070 1162.260 510.000 ;
        RECT 1162.060 496.750 1162.320 497.070 ;
        RECT 1165.740 496.750 1166.000 497.070 ;
        RECT 1165.800 30.930 1165.940 496.750 ;
        RECT 1165.740 30.610 1166.000 30.930 ;
        RECT 1703.480 30.610 1703.740 30.930 ;
        RECT 1703.540 2.400 1703.680 30.610 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1174.450 503.440 1174.770 503.500 ;
        RECT 1183.190 503.440 1183.510 503.500 ;
        RECT 1174.450 503.300 1183.510 503.440 ;
        RECT 1174.450 503.240 1174.770 503.300 ;
        RECT 1183.190 503.240 1183.510 503.300 ;
        RECT 1183.190 141.340 1183.510 141.400 ;
        RECT 1718.170 141.340 1718.490 141.400 ;
        RECT 1183.190 141.200 1718.490 141.340 ;
        RECT 1183.190 141.140 1183.510 141.200 ;
        RECT 1718.170 141.140 1718.490 141.200 ;
      LAYER via ;
        RECT 1174.480 503.240 1174.740 503.500 ;
        RECT 1183.220 503.240 1183.480 503.500 ;
        RECT 1183.220 141.140 1183.480 141.400 ;
        RECT 1718.200 141.140 1718.460 141.400 ;
      LAYER met2 ;
        RECT 1174.610 510.340 1174.890 514.000 ;
        RECT 1174.540 510.000 1174.890 510.340 ;
        RECT 1174.540 503.530 1174.680 510.000 ;
        RECT 1174.480 503.210 1174.740 503.530 ;
        RECT 1183.220 503.210 1183.480 503.530 ;
        RECT 1183.280 141.430 1183.420 503.210 ;
        RECT 1183.220 141.110 1183.480 141.430 ;
        RECT 1718.200 141.110 1718.460 141.430 ;
        RECT 1718.260 17.410 1718.400 141.110 ;
        RECT 1718.260 17.270 1721.620 17.410 ;
        RECT 1721.480 2.400 1721.620 17.270 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.870 503.440 1187.190 503.500 ;
        RECT 1193.310 503.440 1193.630 503.500 ;
        RECT 1186.870 503.300 1193.630 503.440 ;
        RECT 1186.870 503.240 1187.190 503.300 ;
        RECT 1193.310 503.240 1193.630 503.300 ;
        RECT 1193.310 210.360 1193.630 210.420 ;
        RECT 1738.870 210.360 1739.190 210.420 ;
        RECT 1193.310 210.220 1739.190 210.360 ;
        RECT 1193.310 210.160 1193.630 210.220 ;
        RECT 1738.870 210.160 1739.190 210.220 ;
      LAYER via ;
        RECT 1186.900 503.240 1187.160 503.500 ;
        RECT 1193.340 503.240 1193.600 503.500 ;
        RECT 1193.340 210.160 1193.600 210.420 ;
        RECT 1738.900 210.160 1739.160 210.420 ;
      LAYER met2 ;
        RECT 1187.030 510.340 1187.310 514.000 ;
        RECT 1186.960 510.000 1187.310 510.340 ;
        RECT 1186.960 503.530 1187.100 510.000 ;
        RECT 1186.900 503.210 1187.160 503.530 ;
        RECT 1193.340 503.210 1193.600 503.530 ;
        RECT 1193.400 210.450 1193.540 503.210 ;
        RECT 1193.340 210.130 1193.600 210.450 ;
        RECT 1738.900 210.130 1739.160 210.450 ;
        RECT 1738.960 17.410 1739.100 210.130 ;
        RECT 1738.960 17.270 1739.560 17.410 ;
        RECT 1739.420 2.400 1739.560 17.270 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1199.365 386.665 1199.535 409.275 ;
        RECT 1198.905 338.045 1199.075 386.155 ;
        RECT 1199.365 289.765 1199.535 314.755 ;
        RECT 1198.445 241.485 1198.615 255.595 ;
      LAYER mcon ;
        RECT 1199.365 409.105 1199.535 409.275 ;
        RECT 1198.905 385.985 1199.075 386.155 ;
        RECT 1199.365 314.585 1199.535 314.755 ;
        RECT 1198.445 255.425 1198.615 255.595 ;
      LAYER met1 ;
        RECT 1199.290 435.100 1199.610 435.160 ;
        RECT 1199.750 435.100 1200.070 435.160 ;
        RECT 1199.290 434.960 1200.070 435.100 ;
        RECT 1199.290 434.900 1199.610 434.960 ;
        RECT 1199.750 434.900 1200.070 434.960 ;
        RECT 1199.290 409.260 1199.610 409.320 ;
        RECT 1199.095 409.120 1199.610 409.260 ;
        RECT 1199.290 409.060 1199.610 409.120 ;
        RECT 1199.290 386.820 1199.610 386.880 ;
        RECT 1199.095 386.680 1199.610 386.820 ;
        RECT 1199.290 386.620 1199.610 386.680 ;
        RECT 1198.830 386.140 1199.150 386.200 ;
        RECT 1198.635 386.000 1199.150 386.140 ;
        RECT 1198.830 385.940 1199.150 386.000 ;
        RECT 1198.845 338.200 1199.135 338.245 ;
        RECT 1199.290 338.200 1199.610 338.260 ;
        RECT 1198.845 338.060 1199.610 338.200 ;
        RECT 1198.845 338.015 1199.135 338.060 ;
        RECT 1199.290 338.000 1199.610 338.060 ;
        RECT 1199.290 314.740 1199.610 314.800 ;
        RECT 1199.095 314.600 1199.610 314.740 ;
        RECT 1199.290 314.540 1199.610 314.600 ;
        RECT 1198.370 289.920 1198.690 289.980 ;
        RECT 1199.305 289.920 1199.595 289.965 ;
        RECT 1198.370 289.780 1199.595 289.920 ;
        RECT 1198.370 289.720 1198.690 289.780 ;
        RECT 1199.305 289.735 1199.595 289.780 ;
        RECT 1198.370 255.580 1198.690 255.640 ;
        RECT 1198.175 255.440 1198.690 255.580 ;
        RECT 1198.370 255.380 1198.690 255.440 ;
        RECT 1198.370 241.640 1198.690 241.700 ;
        RECT 1198.175 241.500 1198.690 241.640 ;
        RECT 1198.370 241.440 1198.690 241.500 ;
        RECT 1198.370 217.160 1198.690 217.220 ;
        RECT 1752.670 217.160 1752.990 217.220 ;
        RECT 1198.370 217.020 1752.990 217.160 ;
        RECT 1198.370 216.960 1198.690 217.020 ;
        RECT 1752.670 216.960 1752.990 217.020 ;
      LAYER via ;
        RECT 1199.320 434.900 1199.580 435.160 ;
        RECT 1199.780 434.900 1200.040 435.160 ;
        RECT 1199.320 409.060 1199.580 409.320 ;
        RECT 1199.320 386.620 1199.580 386.880 ;
        RECT 1198.860 385.940 1199.120 386.200 ;
        RECT 1199.320 338.000 1199.580 338.260 ;
        RECT 1199.320 314.540 1199.580 314.800 ;
        RECT 1198.400 289.720 1198.660 289.980 ;
        RECT 1198.400 255.380 1198.660 255.640 ;
        RECT 1198.400 241.440 1198.660 241.700 ;
        RECT 1198.400 216.960 1198.660 217.220 ;
        RECT 1752.700 216.960 1752.960 217.220 ;
      LAYER met2 ;
        RECT 1199.450 510.410 1199.730 514.000 ;
        RECT 1198.920 510.270 1199.730 510.410 ;
        RECT 1198.920 483.325 1199.060 510.270 ;
        RECT 1199.450 510.000 1199.730 510.270 ;
        RECT 1198.850 482.955 1199.130 483.325 ;
        RECT 1199.770 482.955 1200.050 483.325 ;
        RECT 1199.840 435.190 1199.980 482.955 ;
        RECT 1199.320 434.870 1199.580 435.190 ;
        RECT 1199.780 434.870 1200.040 435.190 ;
        RECT 1199.380 409.350 1199.520 434.870 ;
        RECT 1199.320 409.030 1199.580 409.350 ;
        RECT 1199.320 386.650 1199.580 386.910 ;
        RECT 1198.920 386.590 1199.580 386.650 ;
        RECT 1198.920 386.510 1199.520 386.590 ;
        RECT 1198.920 386.230 1199.060 386.510 ;
        RECT 1198.860 385.910 1199.120 386.230 ;
        RECT 1199.320 337.970 1199.580 338.290 ;
        RECT 1199.380 314.830 1199.520 337.970 ;
        RECT 1199.320 314.510 1199.580 314.830 ;
        RECT 1198.400 289.690 1198.660 290.010 ;
        RECT 1198.460 255.670 1198.600 289.690 ;
        RECT 1198.400 255.350 1198.660 255.670 ;
        RECT 1198.400 241.410 1198.660 241.730 ;
        RECT 1198.460 217.250 1198.600 241.410 ;
        RECT 1198.400 216.930 1198.660 217.250 ;
        RECT 1752.700 216.930 1752.960 217.250 ;
        RECT 1752.760 17.410 1752.900 216.930 ;
        RECT 1752.760 17.270 1757.040 17.410 ;
        RECT 1756.900 2.400 1757.040 17.270 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
      LAYER via2 ;
        RECT 1198.850 483.000 1199.130 483.280 ;
        RECT 1199.770 483.000 1200.050 483.280 ;
      LAYER met3 ;
        RECT 1198.825 483.290 1199.155 483.305 ;
        RECT 1199.745 483.290 1200.075 483.305 ;
        RECT 1198.825 482.990 1200.075 483.290 ;
        RECT 1198.825 482.975 1199.155 482.990 ;
        RECT 1199.745 482.975 1200.075 482.990 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.010 224.300 1214.330 224.360 ;
        RECT 1773.370 224.300 1773.690 224.360 ;
        RECT 1214.010 224.160 1773.690 224.300 ;
        RECT 1214.010 224.100 1214.330 224.160 ;
        RECT 1773.370 224.100 1773.690 224.160 ;
      LAYER via ;
        RECT 1214.040 224.100 1214.300 224.360 ;
        RECT 1773.400 224.100 1773.660 224.360 ;
      LAYER met2 ;
        RECT 1211.410 510.410 1211.690 514.000 ;
        RECT 1211.410 510.270 1214.240 510.410 ;
        RECT 1211.410 510.000 1211.690 510.270 ;
        RECT 1214.100 224.390 1214.240 510.270 ;
        RECT 1214.040 224.070 1214.300 224.390 ;
        RECT 1773.400 224.070 1773.660 224.390 ;
        RECT 1773.460 17.410 1773.600 224.070 ;
        RECT 1773.460 17.270 1774.980 17.410 ;
        RECT 1774.840 2.400 1774.980 17.270 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1223.670 496.980 1223.990 497.040 ;
        RECT 1227.810 496.980 1228.130 497.040 ;
        RECT 1223.670 496.840 1228.130 496.980 ;
        RECT 1223.670 496.780 1223.990 496.840 ;
        RECT 1227.810 496.780 1228.130 496.840 ;
        RECT 1227.810 231.100 1228.130 231.160 ;
        RECT 1787.170 231.100 1787.490 231.160 ;
        RECT 1227.810 230.960 1787.490 231.100 ;
        RECT 1227.810 230.900 1228.130 230.960 ;
        RECT 1787.170 230.900 1787.490 230.960 ;
      LAYER via ;
        RECT 1223.700 496.780 1223.960 497.040 ;
        RECT 1227.840 496.780 1228.100 497.040 ;
        RECT 1227.840 230.900 1228.100 231.160 ;
        RECT 1787.200 230.900 1787.460 231.160 ;
      LAYER met2 ;
        RECT 1223.830 510.340 1224.110 514.000 ;
        RECT 1223.760 510.000 1224.110 510.340 ;
        RECT 1223.760 497.070 1223.900 510.000 ;
        RECT 1223.700 496.750 1223.960 497.070 ;
        RECT 1227.840 496.750 1228.100 497.070 ;
        RECT 1227.900 231.190 1228.040 496.750 ;
        RECT 1227.840 230.870 1228.100 231.190 ;
        RECT 1787.200 230.870 1787.460 231.190 ;
        RECT 1787.260 17.410 1787.400 230.870 ;
        RECT 1787.260 17.270 1792.920 17.410 ;
        RECT 1792.780 2.400 1792.920 17.270 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.090 496.980 1236.410 497.040 ;
        RECT 1241.150 496.980 1241.470 497.040 ;
        RECT 1236.090 496.840 1241.470 496.980 ;
        RECT 1236.090 496.780 1236.410 496.840 ;
        RECT 1241.150 496.780 1241.470 496.840 ;
        RECT 1241.150 148.480 1241.470 148.540 ;
        RECT 1807.870 148.480 1808.190 148.540 ;
        RECT 1241.150 148.340 1808.190 148.480 ;
        RECT 1241.150 148.280 1241.470 148.340 ;
        RECT 1807.870 148.280 1808.190 148.340 ;
      LAYER via ;
        RECT 1236.120 496.780 1236.380 497.040 ;
        RECT 1241.180 496.780 1241.440 497.040 ;
        RECT 1241.180 148.280 1241.440 148.540 ;
        RECT 1807.900 148.280 1808.160 148.540 ;
      LAYER met2 ;
        RECT 1236.250 510.340 1236.530 514.000 ;
        RECT 1236.180 510.000 1236.530 510.340 ;
        RECT 1236.180 497.070 1236.320 510.000 ;
        RECT 1236.120 496.750 1236.380 497.070 ;
        RECT 1241.180 496.750 1241.440 497.070 ;
        RECT 1241.240 148.570 1241.380 496.750 ;
        RECT 1241.180 148.250 1241.440 148.570 ;
        RECT 1807.900 148.250 1808.160 148.570 ;
        RECT 1807.960 17.410 1808.100 148.250 ;
        RECT 1807.960 17.270 1810.860 17.410 ;
        RECT 1810.720 2.400 1810.860 17.270 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.510 237.900 1248.830 237.960 ;
        RECT 1828.570 237.900 1828.890 237.960 ;
        RECT 1248.510 237.760 1828.890 237.900 ;
        RECT 1248.510 237.700 1248.830 237.760 ;
        RECT 1828.570 237.700 1828.890 237.760 ;
      LAYER via ;
        RECT 1248.540 237.700 1248.800 237.960 ;
        RECT 1828.600 237.700 1828.860 237.960 ;
      LAYER met2 ;
        RECT 1248.670 510.340 1248.950 514.000 ;
        RECT 1248.600 510.000 1248.950 510.340 ;
        RECT 1248.600 237.990 1248.740 510.000 ;
        RECT 1248.540 237.670 1248.800 237.990 ;
        RECT 1828.600 237.670 1828.860 237.990 ;
        RECT 1828.660 2.400 1828.800 237.670 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1261.850 245.040 1262.170 245.100 ;
        RECT 1842.370 245.040 1842.690 245.100 ;
        RECT 1261.850 244.900 1842.690 245.040 ;
        RECT 1261.850 244.840 1262.170 244.900 ;
        RECT 1842.370 244.840 1842.690 244.900 ;
      LAYER via ;
        RECT 1261.880 244.840 1262.140 245.100 ;
        RECT 1842.400 244.840 1842.660 245.100 ;
      LAYER met2 ;
        RECT 1261.090 510.410 1261.370 514.000 ;
        RECT 1261.090 510.270 1262.080 510.410 ;
        RECT 1261.090 510.000 1261.370 510.270 ;
        RECT 1261.940 245.130 1262.080 510.270 ;
        RECT 1261.880 244.810 1262.140 245.130 ;
        RECT 1842.400 244.810 1842.660 245.130 ;
        RECT 1842.460 17.410 1842.600 244.810 ;
        RECT 1842.460 17.270 1846.280 17.410 ;
        RECT 1846.140 2.400 1846.280 17.270 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 155.280 1276.430 155.340 ;
        RECT 1863.070 155.280 1863.390 155.340 ;
        RECT 1276.110 155.140 1863.390 155.280 ;
        RECT 1276.110 155.080 1276.430 155.140 ;
        RECT 1863.070 155.080 1863.390 155.140 ;
      LAYER via ;
        RECT 1276.140 155.080 1276.400 155.340 ;
        RECT 1863.100 155.080 1863.360 155.340 ;
      LAYER met2 ;
        RECT 1273.510 510.410 1273.790 514.000 ;
        RECT 1273.510 510.270 1276.340 510.410 ;
        RECT 1273.510 510.000 1273.790 510.270 ;
        RECT 1276.200 155.370 1276.340 510.270 ;
        RECT 1276.140 155.050 1276.400 155.370 ;
        RECT 1863.100 155.050 1863.360 155.370 ;
        RECT 1863.160 17.410 1863.300 155.050 ;
        RECT 1863.160 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 120.600 496.270 120.660 ;
        RECT 738.370 120.600 738.690 120.660 ;
        RECT 495.950 120.460 738.690 120.600 ;
        RECT 495.950 120.400 496.270 120.460 ;
        RECT 738.370 120.400 738.690 120.460 ;
      LAYER via ;
        RECT 495.980 120.400 496.240 120.660 ;
        RECT 738.400 120.400 738.660 120.660 ;
      LAYER met2 ;
        RECT 494.270 510.410 494.550 514.000 ;
        RECT 494.270 510.270 496.180 510.410 ;
        RECT 494.270 510.000 494.550 510.270 ;
        RECT 496.040 120.690 496.180 510.270 ;
        RECT 495.980 120.370 496.240 120.690 ;
        RECT 738.400 120.370 738.660 120.690 ;
        RECT 738.460 16.900 738.600 120.370 ;
        RECT 738.460 16.760 740.440 16.900 ;
        RECT 740.300 2.400 740.440 16.760 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.450 410.620 1289.770 410.680 ;
        RECT 1876.870 410.620 1877.190 410.680 ;
        RECT 1289.450 410.480 1877.190 410.620 ;
        RECT 1289.450 410.420 1289.770 410.480 ;
        RECT 1876.870 410.420 1877.190 410.480 ;
      LAYER via ;
        RECT 1289.480 410.420 1289.740 410.680 ;
        RECT 1876.900 410.420 1877.160 410.680 ;
      LAYER met2 ;
        RECT 1285.930 510.410 1286.210 514.000 ;
        RECT 1285.930 510.270 1289.680 510.410 ;
        RECT 1285.930 510.000 1286.210 510.270 ;
        RECT 1289.540 410.710 1289.680 510.270 ;
        RECT 1289.480 410.390 1289.740 410.710 ;
        RECT 1876.900 410.390 1877.160 410.710 ;
        RECT 1876.960 17.410 1877.100 410.390 ;
        RECT 1876.960 17.270 1882.160 17.410 ;
        RECT 1882.020 2.400 1882.160 17.270 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1298.190 496.980 1298.510 497.040 ;
        RECT 1303.710 496.980 1304.030 497.040 ;
        RECT 1298.190 496.840 1304.030 496.980 ;
        RECT 1298.190 496.780 1298.510 496.840 ;
        RECT 1303.710 496.780 1304.030 496.840 ;
        RECT 1303.710 162.080 1304.030 162.140 ;
        RECT 1897.570 162.080 1897.890 162.140 ;
        RECT 1303.710 161.940 1897.890 162.080 ;
        RECT 1303.710 161.880 1304.030 161.940 ;
        RECT 1897.570 161.880 1897.890 161.940 ;
      LAYER via ;
        RECT 1298.220 496.780 1298.480 497.040 ;
        RECT 1303.740 496.780 1304.000 497.040 ;
        RECT 1303.740 161.880 1304.000 162.140 ;
        RECT 1897.600 161.880 1897.860 162.140 ;
      LAYER met2 ;
        RECT 1298.350 510.340 1298.630 514.000 ;
        RECT 1298.280 510.000 1298.630 510.340 ;
        RECT 1298.280 497.070 1298.420 510.000 ;
        RECT 1298.220 496.750 1298.480 497.070 ;
        RECT 1303.740 496.750 1304.000 497.070 ;
        RECT 1303.800 162.170 1303.940 496.750 ;
        RECT 1303.740 161.850 1304.000 162.170 ;
        RECT 1897.600 161.850 1897.860 162.170 ;
        RECT 1897.660 17.410 1897.800 161.850 ;
        RECT 1897.660 17.270 1900.100 17.410 ;
        RECT 1899.960 2.400 1900.100 17.270 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 501.060 1310.930 501.120 ;
        RECT 1459.190 501.060 1459.510 501.120 ;
        RECT 1310.610 500.920 1459.510 501.060 ;
        RECT 1310.610 500.860 1310.930 500.920 ;
        RECT 1459.190 500.860 1459.510 500.920 ;
        RECT 1459.190 24.380 1459.510 24.440 ;
        RECT 1917.810 24.380 1918.130 24.440 ;
        RECT 1459.190 24.240 1918.130 24.380 ;
        RECT 1459.190 24.180 1459.510 24.240 ;
        RECT 1917.810 24.180 1918.130 24.240 ;
      LAYER via ;
        RECT 1310.640 500.860 1310.900 501.120 ;
        RECT 1459.220 500.860 1459.480 501.120 ;
        RECT 1459.220 24.180 1459.480 24.440 ;
        RECT 1917.840 24.180 1918.100 24.440 ;
      LAYER met2 ;
        RECT 1310.770 510.340 1311.050 514.000 ;
        RECT 1310.700 510.000 1311.050 510.340 ;
        RECT 1310.700 501.150 1310.840 510.000 ;
        RECT 1310.640 500.830 1310.900 501.150 ;
        RECT 1459.220 500.830 1459.480 501.150 ;
        RECT 1459.280 24.470 1459.420 500.830 ;
        RECT 1459.220 24.150 1459.480 24.470 ;
        RECT 1917.840 24.150 1918.100 24.470 ;
        RECT 1917.900 2.400 1918.040 24.150 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 168.880 1324.730 168.940 ;
        RECT 1932.070 168.880 1932.390 168.940 ;
        RECT 1324.410 168.740 1932.390 168.880 ;
        RECT 1324.410 168.680 1324.730 168.740 ;
        RECT 1932.070 168.680 1932.390 168.740 ;
      LAYER via ;
        RECT 1324.440 168.680 1324.700 168.940 ;
        RECT 1932.100 168.680 1932.360 168.940 ;
      LAYER met2 ;
        RECT 1322.730 510.410 1323.010 514.000 ;
        RECT 1322.730 510.270 1324.640 510.410 ;
        RECT 1322.730 510.000 1323.010 510.270 ;
        RECT 1324.500 168.970 1324.640 510.270 ;
        RECT 1324.440 168.650 1324.700 168.970 ;
        RECT 1932.100 168.650 1932.360 168.970 ;
        RECT 1932.160 17.410 1932.300 168.650 ;
        RECT 1932.160 17.270 1935.520 17.410 ;
        RECT 1935.380 2.400 1935.520 17.270 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 251.840 1338.530 251.900 ;
        RECT 1952.770 251.840 1953.090 251.900 ;
        RECT 1338.210 251.700 1953.090 251.840 ;
        RECT 1338.210 251.640 1338.530 251.700 ;
        RECT 1952.770 251.640 1953.090 251.700 ;
      LAYER via ;
        RECT 1338.240 251.640 1338.500 251.900 ;
        RECT 1952.800 251.640 1953.060 251.900 ;
      LAYER met2 ;
        RECT 1335.150 510.410 1335.430 514.000 ;
        RECT 1335.150 510.270 1338.440 510.410 ;
        RECT 1335.150 510.000 1335.430 510.270 ;
        RECT 1338.300 251.930 1338.440 510.270 ;
        RECT 1338.240 251.610 1338.500 251.930 ;
        RECT 1952.800 251.610 1953.060 251.930 ;
        RECT 1952.860 7.890 1953.000 251.610 ;
        RECT 1952.860 7.750 1953.460 7.890 ;
        RECT 1953.320 2.400 1953.460 7.750 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.410 499.700 1347.730 499.760 ;
        RECT 1351.550 499.700 1351.870 499.760 ;
        RECT 1347.410 499.560 1351.870 499.700 ;
        RECT 1347.410 499.500 1347.730 499.560 ;
        RECT 1351.550 499.500 1351.870 499.560 ;
        RECT 1351.550 258.980 1351.870 259.040 ;
        RECT 1966.570 258.980 1966.890 259.040 ;
        RECT 1351.550 258.840 1966.890 258.980 ;
        RECT 1351.550 258.780 1351.870 258.840 ;
        RECT 1966.570 258.780 1966.890 258.840 ;
      LAYER via ;
        RECT 1347.440 499.500 1347.700 499.760 ;
        RECT 1351.580 499.500 1351.840 499.760 ;
        RECT 1351.580 258.780 1351.840 259.040 ;
        RECT 1966.600 258.780 1966.860 259.040 ;
      LAYER met2 ;
        RECT 1347.570 510.340 1347.850 514.000 ;
        RECT 1347.500 510.000 1347.850 510.340 ;
        RECT 1347.500 499.790 1347.640 510.000 ;
        RECT 1347.440 499.470 1347.700 499.790 ;
        RECT 1351.580 499.470 1351.840 499.790 ;
        RECT 1351.640 259.070 1351.780 499.470 ;
        RECT 1351.580 258.750 1351.840 259.070 ;
        RECT 1966.600 258.750 1966.860 259.070 ;
        RECT 1966.660 17.410 1966.800 258.750 ;
        RECT 1966.660 17.270 1971.400 17.410 ;
        RECT 1971.260 2.400 1971.400 17.270 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.830 503.440 1360.150 503.500 ;
        RECT 1365.810 503.440 1366.130 503.500 ;
        RECT 1359.830 503.300 1366.130 503.440 ;
        RECT 1359.830 503.240 1360.150 503.300 ;
        RECT 1365.810 503.240 1366.130 503.300 ;
        RECT 1365.810 265.780 1366.130 265.840 ;
        RECT 1987.270 265.780 1987.590 265.840 ;
        RECT 1365.810 265.640 1987.590 265.780 ;
        RECT 1365.810 265.580 1366.130 265.640 ;
        RECT 1987.270 265.580 1987.590 265.640 ;
      LAYER via ;
        RECT 1359.860 503.240 1360.120 503.500 ;
        RECT 1365.840 503.240 1366.100 503.500 ;
        RECT 1365.840 265.580 1366.100 265.840 ;
        RECT 1987.300 265.580 1987.560 265.840 ;
      LAYER met2 ;
        RECT 1359.990 510.340 1360.270 514.000 ;
        RECT 1359.920 510.000 1360.270 510.340 ;
        RECT 1359.920 503.530 1360.060 510.000 ;
        RECT 1359.860 503.210 1360.120 503.530 ;
        RECT 1365.840 503.210 1366.100 503.530 ;
        RECT 1365.900 265.870 1366.040 503.210 ;
        RECT 1365.840 265.550 1366.100 265.870 ;
        RECT 1987.300 265.550 1987.560 265.870 ;
        RECT 1987.360 17.410 1987.500 265.550 ;
        RECT 1987.360 17.270 1989.340 17.410 ;
        RECT 1989.200 2.400 1989.340 17.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1372.785 338.045 1372.955 355.895 ;
      LAYER mcon ;
        RECT 1372.785 355.725 1372.955 355.895 ;
      LAYER met1 ;
        RECT 1371.790 448.700 1372.110 448.760 ;
        RECT 1372.710 448.700 1373.030 448.760 ;
        RECT 1371.790 448.560 1373.030 448.700 ;
        RECT 1371.790 448.500 1372.110 448.560 ;
        RECT 1372.710 448.500 1373.030 448.560 ;
        RECT 1372.710 355.880 1373.030 355.940 ;
        RECT 1372.515 355.740 1373.030 355.880 ;
        RECT 1372.710 355.680 1373.030 355.740 ;
        RECT 1372.710 338.200 1373.030 338.260 ;
        RECT 1372.515 338.060 1373.030 338.200 ;
        RECT 1372.710 338.000 1373.030 338.060 ;
        RECT 1371.790 337.520 1372.110 337.580 ;
        RECT 1372.710 337.520 1373.030 337.580 ;
        RECT 1371.790 337.380 1373.030 337.520 ;
        RECT 1371.790 337.320 1372.110 337.380 ;
        RECT 1372.710 337.320 1373.030 337.380 ;
        RECT 1371.790 273.260 1372.110 273.320 ;
        RECT 2001.070 273.260 2001.390 273.320 ;
        RECT 1371.790 273.120 2001.390 273.260 ;
        RECT 1371.790 273.060 1372.110 273.120 ;
        RECT 2001.070 273.060 2001.390 273.120 ;
        RECT 2001.070 20.980 2001.390 21.040 ;
        RECT 2006.590 20.980 2006.910 21.040 ;
        RECT 2001.070 20.840 2006.910 20.980 ;
        RECT 2001.070 20.780 2001.390 20.840 ;
        RECT 2006.590 20.780 2006.910 20.840 ;
      LAYER via ;
        RECT 1371.820 448.500 1372.080 448.760 ;
        RECT 1372.740 448.500 1373.000 448.760 ;
        RECT 1372.740 355.680 1373.000 355.940 ;
        RECT 1372.740 338.000 1373.000 338.260 ;
        RECT 1371.820 337.320 1372.080 337.580 ;
        RECT 1372.740 337.320 1373.000 337.580 ;
        RECT 1371.820 273.060 1372.080 273.320 ;
        RECT 2001.100 273.060 2001.360 273.320 ;
        RECT 2001.100 20.780 2001.360 21.040 ;
        RECT 2006.620 20.780 2006.880 21.040 ;
      LAYER met2 ;
        RECT 1372.410 510.410 1372.690 514.000 ;
        RECT 1371.880 510.270 1372.690 510.410 ;
        RECT 1371.880 483.325 1372.020 510.270 ;
        RECT 1372.410 510.000 1372.690 510.270 ;
        RECT 1371.810 482.955 1372.090 483.325 ;
        RECT 1372.730 482.955 1373.010 483.325 ;
        RECT 1372.800 448.790 1372.940 482.955 ;
        RECT 1371.820 448.530 1372.080 448.790 ;
        RECT 1371.820 448.470 1372.480 448.530 ;
        RECT 1372.740 448.470 1373.000 448.790 ;
        RECT 1371.880 448.390 1372.480 448.470 ;
        RECT 1372.340 447.850 1372.480 448.390 ;
        RECT 1372.340 447.710 1372.940 447.850 ;
        RECT 1372.800 355.970 1372.940 447.710 ;
        RECT 1372.740 355.650 1373.000 355.970 ;
        RECT 1372.740 337.970 1373.000 338.290 ;
        RECT 1372.800 337.610 1372.940 337.970 ;
        RECT 1371.820 337.290 1372.080 337.610 ;
        RECT 1372.740 337.290 1373.000 337.610 ;
        RECT 1371.880 273.350 1372.020 337.290 ;
        RECT 1371.820 273.030 1372.080 273.350 ;
        RECT 2001.100 273.030 2001.360 273.350 ;
        RECT 2001.160 21.070 2001.300 273.030 ;
        RECT 2001.100 20.750 2001.360 21.070 ;
        RECT 2006.620 20.750 2006.880 21.070 ;
        RECT 2006.680 2.400 2006.820 20.750 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 1371.810 483.000 1372.090 483.280 ;
        RECT 1372.730 483.000 1373.010 483.280 ;
      LAYER met3 ;
        RECT 1371.785 483.290 1372.115 483.305 ;
        RECT 1372.705 483.290 1373.035 483.305 ;
        RECT 1371.785 482.990 1373.035 483.290 ;
        RECT 1371.785 482.975 1372.115 482.990 ;
        RECT 1372.705 482.975 1373.035 482.990 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.050 438.160 1386.370 438.220 ;
        RECT 2021.770 438.160 2022.090 438.220 ;
        RECT 1386.050 438.020 2022.090 438.160 ;
        RECT 1386.050 437.960 1386.370 438.020 ;
        RECT 2021.770 437.960 2022.090 438.020 ;
      LAYER via ;
        RECT 1386.080 437.960 1386.340 438.220 ;
        RECT 2021.800 437.960 2022.060 438.220 ;
      LAYER met2 ;
        RECT 1384.830 510.410 1385.110 514.000 ;
        RECT 1384.830 510.270 1386.280 510.410 ;
        RECT 1384.830 510.000 1385.110 510.270 ;
        RECT 1386.140 438.250 1386.280 510.270 ;
        RECT 1386.080 437.930 1386.340 438.250 ;
        RECT 2021.800 437.930 2022.060 438.250 ;
        RECT 2021.860 17.410 2022.000 437.930 ;
        RECT 2021.860 17.270 2024.760 17.410 ;
        RECT 2024.620 2.400 2024.760 17.270 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 176.360 1400.630 176.420 ;
        RECT 2042.930 176.360 2043.250 176.420 ;
        RECT 1400.310 176.220 2043.250 176.360 ;
        RECT 1400.310 176.160 1400.630 176.220 ;
        RECT 2042.930 176.160 2043.250 176.220 ;
      LAYER via ;
        RECT 1400.340 176.160 1400.600 176.420 ;
        RECT 2042.960 176.160 2043.220 176.420 ;
      LAYER met2 ;
        RECT 1397.250 510.410 1397.530 514.000 ;
        RECT 1397.250 510.270 1400.540 510.410 ;
        RECT 1397.250 510.000 1397.530 510.270 ;
        RECT 1400.400 176.450 1400.540 510.270 ;
        RECT 1400.340 176.130 1400.600 176.450 ;
        RECT 2042.960 176.130 2043.220 176.450 ;
        RECT 2043.020 17.410 2043.160 176.130 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 127.740 510.530 127.800 ;
        RECT 752.630 127.740 752.950 127.800 ;
        RECT 510.210 127.600 752.950 127.740 ;
        RECT 510.210 127.540 510.530 127.600 ;
        RECT 752.630 127.540 752.950 127.600 ;
      LAYER via ;
        RECT 510.240 127.540 510.500 127.800 ;
        RECT 752.660 127.540 752.920 127.800 ;
      LAYER met2 ;
        RECT 506.690 510.410 506.970 514.000 ;
        RECT 506.690 510.270 510.440 510.410 ;
        RECT 506.690 510.000 506.970 510.270 ;
        RECT 510.300 127.830 510.440 510.270 ;
        RECT 510.240 127.510 510.500 127.830 ;
        RECT 752.660 127.510 752.920 127.830 ;
        RECT 752.720 16.900 752.860 127.510 ;
        RECT 752.720 16.760 757.920 16.900 ;
        RECT 757.780 2.400 757.920 16.760 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.510 498.680 1409.830 498.740 ;
        RECT 1414.110 498.680 1414.430 498.740 ;
        RECT 1409.510 498.540 1414.430 498.680 ;
        RECT 1409.510 498.480 1409.830 498.540 ;
        RECT 1414.110 498.480 1414.430 498.540 ;
        RECT 1414.110 362.680 1414.430 362.740 ;
        RECT 2056.270 362.680 2056.590 362.740 ;
        RECT 1414.110 362.540 2056.590 362.680 ;
        RECT 1414.110 362.480 1414.430 362.540 ;
        RECT 2056.270 362.480 2056.590 362.540 ;
      LAYER via ;
        RECT 1409.540 498.480 1409.800 498.740 ;
        RECT 1414.140 498.480 1414.400 498.740 ;
        RECT 1414.140 362.480 1414.400 362.740 ;
        RECT 2056.300 362.480 2056.560 362.740 ;
      LAYER met2 ;
        RECT 1409.670 510.340 1409.950 514.000 ;
        RECT 1409.600 510.000 1409.950 510.340 ;
        RECT 1409.600 498.770 1409.740 510.000 ;
        RECT 1409.540 498.450 1409.800 498.770 ;
        RECT 1414.140 498.450 1414.400 498.770 ;
        RECT 1414.200 362.770 1414.340 498.450 ;
        RECT 1414.140 362.450 1414.400 362.770 ;
        RECT 2056.300 362.450 2056.560 362.770 ;
        RECT 2056.360 17.410 2056.500 362.450 ;
        RECT 2056.360 17.270 2060.640 17.410 ;
        RECT 2060.500 2.400 2060.640 17.270 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.930 496.980 1422.250 497.040 ;
        RECT 1427.910 496.980 1428.230 497.040 ;
        RECT 1421.930 496.840 1428.230 496.980 ;
        RECT 1421.930 496.780 1422.250 496.840 ;
        RECT 1427.910 496.780 1428.230 496.840 ;
        RECT 1427.910 355.880 1428.230 355.940 ;
        RECT 2076.970 355.880 2077.290 355.940 ;
        RECT 1427.910 355.740 2077.290 355.880 ;
        RECT 1427.910 355.680 1428.230 355.740 ;
        RECT 2076.970 355.680 2077.290 355.740 ;
      LAYER via ;
        RECT 1421.960 496.780 1422.220 497.040 ;
        RECT 1427.940 496.780 1428.200 497.040 ;
        RECT 1427.940 355.680 1428.200 355.940 ;
        RECT 2077.000 355.680 2077.260 355.940 ;
      LAYER met2 ;
        RECT 1422.090 510.340 1422.370 514.000 ;
        RECT 1422.020 510.000 1422.370 510.340 ;
        RECT 1422.020 497.070 1422.160 510.000 ;
        RECT 1421.960 496.750 1422.220 497.070 ;
        RECT 1427.940 496.750 1428.200 497.070 ;
        RECT 1428.000 355.970 1428.140 496.750 ;
        RECT 1427.940 355.650 1428.200 355.970 ;
        RECT 2077.000 355.650 2077.260 355.970 ;
        RECT 2077.060 17.410 2077.200 355.650 ;
        RECT 2077.060 17.270 2078.580 17.410 ;
        RECT 2078.440 2.400 2078.580 17.270 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 280.060 1435.130 280.120 ;
        RECT 2090.770 280.060 2091.090 280.120 ;
        RECT 1434.810 279.920 2091.090 280.060 ;
        RECT 1434.810 279.860 1435.130 279.920 ;
        RECT 2090.770 279.860 2091.090 279.920 ;
      LAYER via ;
        RECT 1434.840 279.860 1435.100 280.120 ;
        RECT 2090.800 279.860 2091.060 280.120 ;
      LAYER met2 ;
        RECT 1434.510 510.340 1434.790 514.000 ;
        RECT 1434.440 510.000 1434.790 510.340 ;
        RECT 1434.440 497.490 1434.580 510.000 ;
        RECT 1434.440 497.350 1435.040 497.490 ;
        RECT 1434.900 280.150 1435.040 497.350 ;
        RECT 1434.840 279.830 1435.100 280.150 ;
        RECT 2090.800 279.830 2091.060 280.150 ;
        RECT 2090.860 17.410 2091.000 279.830 ;
        RECT 2090.860 17.270 2096.060 17.410 ;
        RECT 2095.920 2.400 2096.060 17.270 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1446.310 500.720 1446.630 500.780 ;
        RECT 1610.990 500.720 1611.310 500.780 ;
        RECT 1446.310 500.580 1611.310 500.720 ;
        RECT 1446.310 500.520 1446.630 500.580 ;
        RECT 1610.990 500.520 1611.310 500.580 ;
        RECT 1610.990 348.740 1611.310 348.800 ;
        RECT 2111.470 348.740 2111.790 348.800 ;
        RECT 1610.990 348.600 2111.790 348.740 ;
        RECT 1610.990 348.540 1611.310 348.600 ;
        RECT 2111.470 348.540 2111.790 348.600 ;
      LAYER via ;
        RECT 1446.340 500.520 1446.600 500.780 ;
        RECT 1611.020 500.520 1611.280 500.780 ;
        RECT 1611.020 348.540 1611.280 348.800 ;
        RECT 2111.500 348.540 2111.760 348.800 ;
      LAYER met2 ;
        RECT 1446.470 510.340 1446.750 514.000 ;
        RECT 1446.400 510.000 1446.750 510.340 ;
        RECT 1446.400 500.810 1446.540 510.000 ;
        RECT 1446.340 500.490 1446.600 500.810 ;
        RECT 1611.020 500.490 1611.280 500.810 ;
        RECT 1611.080 348.830 1611.220 500.490 ;
        RECT 1611.020 348.510 1611.280 348.830 ;
        RECT 2111.500 348.510 2111.760 348.830 ;
        RECT 2111.560 17.410 2111.700 348.510 ;
        RECT 2111.560 17.270 2114.000 17.410 ;
        RECT 2113.860 2.400 2114.000 17.270 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 342.280 1462.730 342.340 ;
        RECT 2125.270 342.280 2125.590 342.340 ;
        RECT 1462.410 342.140 2125.590 342.280 ;
        RECT 1462.410 342.080 1462.730 342.140 ;
        RECT 2125.270 342.080 2125.590 342.140 ;
        RECT 2125.270 16.900 2125.590 16.960 ;
        RECT 2131.710 16.900 2132.030 16.960 ;
        RECT 2125.270 16.760 2132.030 16.900 ;
        RECT 2125.270 16.700 2125.590 16.760 ;
        RECT 2131.710 16.700 2132.030 16.760 ;
      LAYER via ;
        RECT 1462.440 342.080 1462.700 342.340 ;
        RECT 2125.300 342.080 2125.560 342.340 ;
        RECT 2125.300 16.700 2125.560 16.960 ;
        RECT 2131.740 16.700 2132.000 16.960 ;
      LAYER met2 ;
        RECT 1458.890 510.410 1459.170 514.000 ;
        RECT 1458.890 510.270 1462.640 510.410 ;
        RECT 1458.890 510.000 1459.170 510.270 ;
        RECT 1462.500 342.370 1462.640 510.270 ;
        RECT 1462.440 342.050 1462.700 342.370 ;
        RECT 2125.300 342.050 2125.560 342.370 ;
        RECT 2125.360 16.990 2125.500 342.050 ;
        RECT 2125.300 16.670 2125.560 16.990 ;
        RECT 2131.740 16.670 2132.000 16.990 ;
        RECT 2131.800 2.400 2131.940 16.670 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.150 496.980 1471.470 497.040 ;
        RECT 1476.210 496.980 1476.530 497.040 ;
        RECT 1471.150 496.840 1476.530 496.980 ;
        RECT 1471.150 496.780 1471.470 496.840 ;
        RECT 1476.210 496.780 1476.530 496.840 ;
        RECT 1476.210 334.800 1476.530 334.860 ;
        RECT 2145.970 334.800 2146.290 334.860 ;
        RECT 1476.210 334.660 2146.290 334.800 ;
        RECT 1476.210 334.600 1476.530 334.660 ;
        RECT 2145.970 334.600 2146.290 334.660 ;
      LAYER via ;
        RECT 1471.180 496.780 1471.440 497.040 ;
        RECT 1476.240 496.780 1476.500 497.040 ;
        RECT 1476.240 334.600 1476.500 334.860 ;
        RECT 2146.000 334.600 2146.260 334.860 ;
      LAYER met2 ;
        RECT 1471.310 510.340 1471.590 514.000 ;
        RECT 1471.240 510.000 1471.590 510.340 ;
        RECT 1471.240 497.070 1471.380 510.000 ;
        RECT 1471.180 496.750 1471.440 497.070 ;
        RECT 1476.240 496.750 1476.500 497.070 ;
        RECT 1476.300 334.890 1476.440 496.750 ;
        RECT 1476.240 334.570 1476.500 334.890 ;
        RECT 2146.000 334.570 2146.260 334.890 ;
        RECT 2146.060 17.410 2146.200 334.570 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.570 496.980 1483.890 497.040 ;
        RECT 1489.550 496.980 1489.870 497.040 ;
        RECT 1483.570 496.840 1489.870 496.980 ;
        RECT 1483.570 496.780 1483.890 496.840 ;
        RECT 1489.550 496.780 1489.870 496.840 ;
        RECT 1489.550 328.000 1489.870 328.060 ;
        RECT 2166.670 328.000 2166.990 328.060 ;
        RECT 1489.550 327.860 2166.990 328.000 ;
        RECT 1489.550 327.800 1489.870 327.860 ;
        RECT 2166.670 327.800 2166.990 327.860 ;
      LAYER via ;
        RECT 1483.600 496.780 1483.860 497.040 ;
        RECT 1489.580 496.780 1489.840 497.040 ;
        RECT 1489.580 327.800 1489.840 328.060 ;
        RECT 2166.700 327.800 2166.960 328.060 ;
      LAYER met2 ;
        RECT 1483.730 510.340 1484.010 514.000 ;
        RECT 1483.660 510.000 1484.010 510.340 ;
        RECT 1483.660 497.070 1483.800 510.000 ;
        RECT 1483.600 496.750 1483.860 497.070 ;
        RECT 1489.580 496.750 1489.840 497.070 ;
        RECT 1489.640 328.090 1489.780 496.750 ;
        RECT 1489.580 327.770 1489.840 328.090 ;
        RECT 2166.700 327.770 2166.960 328.090 ;
        RECT 2166.760 17.410 2166.900 327.770 ;
        RECT 2166.760 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 286.520 1497.230 286.580 ;
        RECT 2180.470 286.520 2180.790 286.580 ;
        RECT 1496.910 286.380 2180.790 286.520 ;
        RECT 1496.910 286.320 1497.230 286.380 ;
        RECT 2180.470 286.320 2180.790 286.380 ;
      LAYER via ;
        RECT 1496.940 286.320 1497.200 286.580 ;
        RECT 2180.500 286.320 2180.760 286.580 ;
      LAYER met2 ;
        RECT 1496.150 510.410 1496.430 514.000 ;
        RECT 1496.150 510.270 1497.140 510.410 ;
        RECT 1496.150 510.000 1496.430 510.270 ;
        RECT 1497.000 286.610 1497.140 510.270 ;
        RECT 1496.940 286.290 1497.200 286.610 ;
        RECT 2180.500 286.290 2180.760 286.610 ;
        RECT 2180.560 17.410 2180.700 286.290 ;
        RECT 2180.560 17.270 2185.300 17.410 ;
        RECT 2185.160 2.400 2185.300 17.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.710 321.200 1511.030 321.260 ;
        RECT 2201.170 321.200 2201.490 321.260 ;
        RECT 1510.710 321.060 2201.490 321.200 ;
        RECT 1510.710 321.000 1511.030 321.060 ;
        RECT 2201.170 321.000 2201.490 321.060 ;
      LAYER via ;
        RECT 1510.740 321.000 1511.000 321.260 ;
        RECT 2201.200 321.000 2201.460 321.260 ;
      LAYER met2 ;
        RECT 1508.570 510.410 1508.850 514.000 ;
        RECT 1508.570 510.270 1510.940 510.410 ;
        RECT 1508.570 510.000 1508.850 510.270 ;
        RECT 1510.800 321.290 1510.940 510.270 ;
        RECT 1510.740 320.970 1511.000 321.290 ;
        RECT 2201.200 320.970 2201.460 321.290 ;
        RECT 2201.260 17.410 2201.400 320.970 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1520.830 496.980 1521.150 497.040 ;
        RECT 1524.510 496.980 1524.830 497.040 ;
        RECT 1520.830 496.840 1524.830 496.980 ;
        RECT 1520.830 496.780 1521.150 496.840 ;
        RECT 1524.510 496.780 1524.830 496.840 ;
        RECT 1524.510 100.200 1524.830 100.260 ;
        RECT 2215.430 100.200 2215.750 100.260 ;
        RECT 1524.510 100.060 2215.750 100.200 ;
        RECT 1524.510 100.000 1524.830 100.060 ;
        RECT 2215.430 100.000 2215.750 100.060 ;
      LAYER via ;
        RECT 1520.860 496.780 1521.120 497.040 ;
        RECT 1524.540 496.780 1524.800 497.040 ;
        RECT 1524.540 100.000 1524.800 100.260 ;
        RECT 2215.460 100.000 2215.720 100.260 ;
      LAYER met2 ;
        RECT 1520.990 510.340 1521.270 514.000 ;
        RECT 1520.920 510.000 1521.270 510.340 ;
        RECT 1520.920 497.070 1521.060 510.000 ;
        RECT 1520.860 496.750 1521.120 497.070 ;
        RECT 1524.540 496.750 1524.800 497.070 ;
        RECT 1524.600 100.290 1524.740 496.750 ;
        RECT 1524.540 99.970 1524.800 100.290 ;
        RECT 2215.460 99.970 2215.720 100.290 ;
        RECT 2215.520 17.410 2215.660 99.970 ;
        RECT 2215.520 17.270 2221.180 17.410 ;
        RECT 2221.040 2.400 2221.180 17.270 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 518.950 498.000 519.270 498.060 ;
        RECT 524.010 498.000 524.330 498.060 ;
        RECT 518.950 497.860 524.330 498.000 ;
        RECT 518.950 497.800 519.270 497.860 ;
        RECT 524.010 497.800 524.330 497.860 ;
        RECT 524.010 134.540 524.330 134.600 ;
        RECT 772.870 134.540 773.190 134.600 ;
        RECT 524.010 134.400 773.190 134.540 ;
        RECT 524.010 134.340 524.330 134.400 ;
        RECT 772.870 134.340 773.190 134.400 ;
      LAYER via ;
        RECT 518.980 497.800 519.240 498.060 ;
        RECT 524.040 497.800 524.300 498.060 ;
        RECT 524.040 134.340 524.300 134.600 ;
        RECT 772.900 134.340 773.160 134.600 ;
      LAYER met2 ;
        RECT 519.110 510.340 519.390 514.000 ;
        RECT 519.040 510.000 519.390 510.340 ;
        RECT 519.040 498.090 519.180 510.000 ;
        RECT 518.980 497.770 519.240 498.090 ;
        RECT 524.040 497.770 524.300 498.090 ;
        RECT 524.100 134.630 524.240 497.770 ;
        RECT 524.040 134.310 524.300 134.630 ;
        RECT 772.900 134.310 773.160 134.630 ;
        RECT 772.960 17.410 773.100 134.310 ;
        RECT 772.960 17.270 775.860 17.410 ;
        RECT 775.720 2.400 775.860 17.270 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1533.250 497.660 1533.570 497.720 ;
        RECT 1569.590 497.660 1569.910 497.720 ;
        RECT 1533.250 497.520 1569.910 497.660 ;
        RECT 1533.250 497.460 1533.570 497.520 ;
        RECT 1569.590 497.460 1569.910 497.520 ;
        RECT 1569.590 314.400 1569.910 314.460 ;
        RECT 2235.670 314.400 2235.990 314.460 ;
        RECT 1569.590 314.260 2235.990 314.400 ;
        RECT 1569.590 314.200 1569.910 314.260 ;
        RECT 2235.670 314.200 2235.990 314.260 ;
      LAYER via ;
        RECT 1533.280 497.460 1533.540 497.720 ;
        RECT 1569.620 497.460 1569.880 497.720 ;
        RECT 1569.620 314.200 1569.880 314.460 ;
        RECT 2235.700 314.200 2235.960 314.460 ;
      LAYER met2 ;
        RECT 1533.410 510.340 1533.690 514.000 ;
        RECT 1533.340 510.000 1533.690 510.340 ;
        RECT 1533.340 497.750 1533.480 510.000 ;
        RECT 1533.280 497.430 1533.540 497.750 ;
        RECT 1569.620 497.430 1569.880 497.750 ;
        RECT 1569.680 314.490 1569.820 497.430 ;
        RECT 1569.620 314.170 1569.880 314.490 ;
        RECT 2235.700 314.170 2235.960 314.490 ;
        RECT 2235.760 17.410 2235.900 314.170 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.670 496.980 1545.990 497.040 ;
        RECT 1552.110 496.980 1552.430 497.040 ;
        RECT 1545.670 496.840 1552.430 496.980 ;
        RECT 1545.670 496.780 1545.990 496.840 ;
        RECT 1552.110 496.780 1552.430 496.840 ;
        RECT 1552.110 307.260 1552.430 307.320 ;
        RECT 2256.370 307.260 2256.690 307.320 ;
        RECT 1552.110 307.120 2256.690 307.260 ;
        RECT 1552.110 307.060 1552.430 307.120 ;
        RECT 2256.370 307.060 2256.690 307.120 ;
      LAYER via ;
        RECT 1545.700 496.780 1545.960 497.040 ;
        RECT 1552.140 496.780 1552.400 497.040 ;
        RECT 1552.140 307.060 1552.400 307.320 ;
        RECT 2256.400 307.060 2256.660 307.320 ;
      LAYER met2 ;
        RECT 1545.830 510.340 1546.110 514.000 ;
        RECT 1545.760 510.000 1546.110 510.340 ;
        RECT 1545.760 497.070 1545.900 510.000 ;
        RECT 1545.700 496.750 1545.960 497.070 ;
        RECT 1552.140 496.750 1552.400 497.070 ;
        RECT 1552.200 307.350 1552.340 496.750 ;
        RECT 1552.140 307.030 1552.400 307.350 ;
        RECT 2256.400 307.030 2256.660 307.350 ;
        RECT 2256.460 2.400 2256.600 307.030 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1557.630 497.320 1557.950 497.380 ;
        RECT 1590.290 497.320 1590.610 497.380 ;
        RECT 1557.630 497.180 1590.610 497.320 ;
        RECT 1557.630 497.120 1557.950 497.180 ;
        RECT 1590.290 497.120 1590.610 497.180 ;
        RECT 1590.290 107.340 1590.610 107.400 ;
        RECT 2270.170 107.340 2270.490 107.400 ;
        RECT 1590.290 107.200 2270.490 107.340 ;
        RECT 1590.290 107.140 1590.610 107.200 ;
        RECT 2270.170 107.140 2270.490 107.200 ;
      LAYER via ;
        RECT 1557.660 497.120 1557.920 497.380 ;
        RECT 1590.320 497.120 1590.580 497.380 ;
        RECT 1590.320 107.140 1590.580 107.400 ;
        RECT 2270.200 107.140 2270.460 107.400 ;
      LAYER met2 ;
        RECT 1557.790 510.340 1558.070 514.000 ;
        RECT 1557.720 510.000 1558.070 510.340 ;
        RECT 1557.720 497.410 1557.860 510.000 ;
        RECT 1557.660 497.090 1557.920 497.410 ;
        RECT 1590.320 497.090 1590.580 497.410 ;
        RECT 1590.380 107.430 1590.520 497.090 ;
        RECT 1590.320 107.110 1590.580 107.430 ;
        RECT 2270.200 107.110 2270.460 107.430 ;
        RECT 2270.260 17.410 2270.400 107.110 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 183.160 1573.130 183.220 ;
        RECT 2290.870 183.160 2291.190 183.220 ;
        RECT 1572.810 183.020 2291.190 183.160 ;
        RECT 1572.810 182.960 1573.130 183.020 ;
        RECT 2290.870 182.960 2291.190 183.020 ;
      LAYER via ;
        RECT 1572.840 182.960 1573.100 183.220 ;
        RECT 2290.900 182.960 2291.160 183.220 ;
      LAYER met2 ;
        RECT 1570.210 510.410 1570.490 514.000 ;
        RECT 1570.210 510.270 1573.040 510.410 ;
        RECT 1570.210 510.000 1570.490 510.270 ;
        RECT 1572.900 183.250 1573.040 510.270 ;
        RECT 1572.840 182.930 1573.100 183.250 ;
        RECT 2290.900 182.930 2291.160 183.250 ;
        RECT 2290.960 17.410 2291.100 182.930 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.470 496.980 1582.790 497.040 ;
        RECT 1586.150 496.980 1586.470 497.040 ;
        RECT 1582.470 496.840 1586.470 496.980 ;
        RECT 1582.470 496.780 1582.790 496.840 ;
        RECT 1586.150 496.780 1586.470 496.840 ;
        RECT 1586.150 300.120 1586.470 300.180 ;
        RECT 2304.670 300.120 2304.990 300.180 ;
        RECT 1586.150 299.980 2304.990 300.120 ;
        RECT 1586.150 299.920 1586.470 299.980 ;
        RECT 2304.670 299.920 2304.990 299.980 ;
      LAYER via ;
        RECT 1582.500 496.780 1582.760 497.040 ;
        RECT 1586.180 496.780 1586.440 497.040 ;
        RECT 1586.180 299.920 1586.440 300.180 ;
        RECT 2304.700 299.920 2304.960 300.180 ;
      LAYER met2 ;
        RECT 1582.630 510.340 1582.910 514.000 ;
        RECT 1582.560 510.000 1582.910 510.340 ;
        RECT 1582.560 497.070 1582.700 510.000 ;
        RECT 1582.500 496.750 1582.760 497.070 ;
        RECT 1586.180 496.750 1586.440 497.070 ;
        RECT 1586.240 300.210 1586.380 496.750 ;
        RECT 1586.180 299.890 1586.440 300.210 ;
        RECT 2304.700 299.890 2304.960 300.210 ;
        RECT 2304.760 17.410 2304.900 299.890 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1594.890 496.980 1595.210 497.040 ;
        RECT 1599.950 496.980 1600.270 497.040 ;
        RECT 1594.890 496.840 1600.270 496.980 ;
        RECT 1594.890 496.780 1595.210 496.840 ;
        RECT 1599.950 496.780 1600.270 496.840 ;
        RECT 1599.950 293.660 1600.270 293.720 ;
        RECT 2325.370 293.660 2325.690 293.720 ;
        RECT 1599.950 293.520 2325.690 293.660 ;
        RECT 1599.950 293.460 1600.270 293.520 ;
        RECT 2325.370 293.460 2325.690 293.520 ;
      LAYER via ;
        RECT 1594.920 496.780 1595.180 497.040 ;
        RECT 1599.980 496.780 1600.240 497.040 ;
        RECT 1599.980 293.460 1600.240 293.720 ;
        RECT 2325.400 293.460 2325.660 293.720 ;
      LAYER met2 ;
        RECT 1595.050 510.340 1595.330 514.000 ;
        RECT 1594.980 510.000 1595.330 510.340 ;
        RECT 1594.980 497.070 1595.120 510.000 ;
        RECT 1594.920 496.750 1595.180 497.070 ;
        RECT 1599.980 496.750 1600.240 497.070 ;
        RECT 1600.040 293.750 1600.180 496.750 ;
        RECT 1599.980 293.430 1600.240 293.750 ;
        RECT 2325.400 293.430 2325.660 293.750 ;
        RECT 2325.460 17.410 2325.600 293.430 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1606.850 114.140 1607.170 114.200 ;
        RECT 2339.630 114.140 2339.950 114.200 ;
        RECT 1606.850 114.000 2339.950 114.140 ;
        RECT 1606.850 113.940 1607.170 114.000 ;
        RECT 2339.630 113.940 2339.950 114.000 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.610 16.900 2345.930 16.960 ;
        RECT 2339.630 16.760 2345.930 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.610 16.700 2345.930 16.760 ;
      LAYER via ;
        RECT 1606.880 113.940 1607.140 114.200 ;
        RECT 2339.660 113.940 2339.920 114.200 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.640 16.700 2345.900 16.960 ;
      LAYER met2 ;
        RECT 1607.470 510.410 1607.750 514.000 ;
        RECT 1606.940 510.270 1607.750 510.410 ;
        RECT 1606.940 114.230 1607.080 510.270 ;
        RECT 1607.470 510.000 1607.750 510.270 ;
        RECT 1606.880 113.910 1607.140 114.230 ;
        RECT 2339.660 113.910 2339.920 114.230 ;
        RECT 2339.720 16.990 2339.860 113.910 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.640 16.670 2345.900 16.990 ;
        RECT 2345.700 2.400 2345.840 16.670 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1620.650 120.940 1620.970 121.000 ;
        RECT 2359.870 120.940 2360.190 121.000 ;
        RECT 1620.650 120.800 2360.190 120.940 ;
        RECT 1620.650 120.740 1620.970 120.800 ;
        RECT 2359.870 120.740 2360.190 120.800 ;
      LAYER via ;
        RECT 1620.680 120.740 1620.940 121.000 ;
        RECT 2359.900 120.740 2360.160 121.000 ;
      LAYER met2 ;
        RECT 1619.890 510.410 1620.170 514.000 ;
        RECT 1619.890 510.270 1620.880 510.410 ;
        RECT 1619.890 510.000 1620.170 510.270 ;
        RECT 1620.740 121.030 1620.880 510.270 ;
        RECT 1620.680 120.710 1620.940 121.030 ;
        RECT 2359.900 120.710 2360.160 121.030 ;
        RECT 2359.960 17.410 2360.100 120.710 ;
        RECT 2359.960 17.270 2363.780 17.410 ;
        RECT 2363.640 2.400 2363.780 17.270 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.910 197.100 1635.230 197.160 ;
        RECT 2380.570 197.100 2380.890 197.160 ;
        RECT 1634.910 196.960 2380.890 197.100 ;
        RECT 1634.910 196.900 1635.230 196.960 ;
        RECT 2380.570 196.900 2380.890 196.960 ;
      LAYER via ;
        RECT 1634.940 196.900 1635.200 197.160 ;
        RECT 2380.600 196.900 2380.860 197.160 ;
      LAYER met2 ;
        RECT 1632.310 510.410 1632.590 514.000 ;
        RECT 1632.310 510.270 1635.140 510.410 ;
        RECT 1632.310 510.000 1632.590 510.270 ;
        RECT 1635.000 197.190 1635.140 510.270 ;
        RECT 1634.940 196.870 1635.200 197.190 ;
        RECT 2380.600 196.870 2380.860 197.190 ;
        RECT 2380.660 17.410 2380.800 196.870 ;
        RECT 2380.660 17.270 2381.720 17.410 ;
        RECT 2381.580 2.400 2381.720 17.270 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1644.570 496.980 1644.890 497.040 ;
        RECT 1659.290 496.980 1659.610 497.040 ;
        RECT 1644.570 496.840 1659.610 496.980 ;
        RECT 1644.570 496.780 1644.890 496.840 ;
        RECT 1659.290 496.780 1659.610 496.840 ;
        RECT 1659.290 189.960 1659.610 190.020 ;
        RECT 2394.370 189.960 2394.690 190.020 ;
        RECT 1659.290 189.820 2394.690 189.960 ;
        RECT 1659.290 189.760 1659.610 189.820 ;
        RECT 2394.370 189.760 2394.690 189.820 ;
      LAYER via ;
        RECT 1644.600 496.780 1644.860 497.040 ;
        RECT 1659.320 496.780 1659.580 497.040 ;
        RECT 1659.320 189.760 1659.580 190.020 ;
        RECT 2394.400 189.760 2394.660 190.020 ;
      LAYER met2 ;
        RECT 1644.730 510.340 1645.010 514.000 ;
        RECT 1644.660 510.000 1645.010 510.340 ;
        RECT 1644.660 497.070 1644.800 510.000 ;
        RECT 1644.600 496.750 1644.860 497.070 ;
        RECT 1659.320 496.750 1659.580 497.070 ;
        RECT 1659.380 190.050 1659.520 496.750 ;
        RECT 1659.320 189.730 1659.580 190.050 ;
        RECT 2394.400 189.730 2394.660 190.050 ;
        RECT 2394.460 17.410 2394.600 189.730 ;
        RECT 2394.460 17.270 2399.660 17.410 ;
        RECT 2399.520 2.400 2399.660 17.270 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.450 148.140 530.770 148.200 ;
        RECT 794.030 148.140 794.350 148.200 ;
        RECT 530.450 148.000 794.350 148.140 ;
        RECT 530.450 147.940 530.770 148.000 ;
        RECT 794.030 147.940 794.350 148.000 ;
      LAYER via ;
        RECT 530.480 147.940 530.740 148.200 ;
        RECT 794.060 147.940 794.320 148.200 ;
      LAYER met2 ;
        RECT 531.070 510.410 531.350 514.000 ;
        RECT 530.540 510.270 531.350 510.410 ;
        RECT 530.540 148.230 530.680 510.270 ;
        RECT 531.070 510.000 531.350 510.270 ;
        RECT 530.480 147.910 530.740 148.230 ;
        RECT 794.060 147.910 794.320 148.230 ;
        RECT 794.120 7.210 794.260 147.910 ;
        RECT 793.660 7.070 794.260 7.210 ;
        RECT 793.660 2.400 793.800 7.070 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 427.410 72.320 427.730 72.380 ;
        RECT 634.870 72.320 635.190 72.380 ;
        RECT 427.410 72.180 635.190 72.320 ;
        RECT 427.410 72.120 427.730 72.180 ;
        RECT 634.870 72.120 635.190 72.180 ;
        RECT 634.870 2.960 635.190 3.020 ;
        RECT 639.010 2.960 639.330 3.020 ;
        RECT 634.870 2.820 639.330 2.960 ;
        RECT 634.870 2.760 635.190 2.820 ;
        RECT 639.010 2.760 639.330 2.820 ;
      LAYER via ;
        RECT 427.440 72.120 427.700 72.380 ;
        RECT 634.900 72.120 635.160 72.380 ;
        RECT 634.900 2.760 635.160 3.020 ;
        RECT 639.040 2.760 639.300 3.020 ;
      LAYER met2 ;
        RECT 423.890 510.410 424.170 514.000 ;
        RECT 423.890 510.270 427.640 510.410 ;
        RECT 423.890 510.000 424.170 510.270 ;
        RECT 427.500 72.410 427.640 510.270 ;
        RECT 427.440 72.090 427.700 72.410 ;
        RECT 634.900 72.090 635.160 72.410 ;
        RECT 634.960 3.050 635.100 72.090 ;
        RECT 634.900 2.730 635.160 3.050 ;
        RECT 639.040 2.730 639.300 3.050 ;
        RECT 639.100 2.400 639.240 2.730 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 128.080 1662.830 128.140 ;
        RECT 2421.970 128.080 2422.290 128.140 ;
        RECT 1662.510 127.940 2422.290 128.080 ;
        RECT 1662.510 127.880 1662.830 127.940 ;
        RECT 2421.970 127.880 2422.290 127.940 ;
      LAYER via ;
        RECT 1662.540 127.880 1662.800 128.140 ;
        RECT 2422.000 127.880 2422.260 128.140 ;
      LAYER met2 ;
        RECT 1661.290 510.410 1661.570 514.000 ;
        RECT 1661.290 510.270 1662.740 510.410 ;
        RECT 1661.290 510.000 1661.570 510.270 ;
        RECT 1662.600 128.170 1662.740 510.270 ;
        RECT 1662.540 127.850 1662.800 128.170 ;
        RECT 2422.000 127.850 2422.260 128.170 ;
        RECT 2422.060 17.410 2422.200 127.850 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 134.880 1676.630 134.940 ;
        RECT 2435.770 134.880 2436.090 134.940 ;
        RECT 1676.310 134.740 2436.090 134.880 ;
        RECT 1676.310 134.680 1676.630 134.740 ;
        RECT 2435.770 134.680 2436.090 134.740 ;
        RECT 2435.770 62.120 2436.090 62.180 ;
        RECT 2440.830 62.120 2441.150 62.180 ;
        RECT 2435.770 61.980 2441.150 62.120 ;
        RECT 2435.770 61.920 2436.090 61.980 ;
        RECT 2440.830 61.920 2441.150 61.980 ;
      LAYER via ;
        RECT 1676.340 134.680 1676.600 134.940 ;
        RECT 2435.800 134.680 2436.060 134.940 ;
        RECT 2435.800 61.920 2436.060 62.180 ;
        RECT 2440.860 61.920 2441.120 62.180 ;
      LAYER met2 ;
        RECT 1673.250 510.410 1673.530 514.000 ;
        RECT 1673.250 510.270 1676.540 510.410 ;
        RECT 1673.250 510.000 1673.530 510.270 ;
        RECT 1676.400 134.970 1676.540 510.270 ;
        RECT 1676.340 134.650 1676.600 134.970 ;
        RECT 2435.800 134.650 2436.060 134.970 ;
        RECT 2435.860 62.210 2436.000 134.650 ;
        RECT 2435.800 61.890 2436.060 62.210 ;
        RECT 2440.860 61.890 2441.120 62.210 ;
        RECT 2440.920 2.400 2441.060 61.890 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2456.545 48.365 2456.715 96.475 ;
      LAYER mcon ;
        RECT 2456.545 96.305 2456.715 96.475 ;
      LAYER met1 ;
        RECT 1685.510 496.980 1685.830 497.040 ;
        RECT 1689.650 496.980 1689.970 497.040 ;
        RECT 1685.510 496.840 1689.970 496.980 ;
        RECT 1685.510 496.780 1685.830 496.840 ;
        RECT 1689.650 496.780 1689.970 496.840 ;
        RECT 1689.650 141.680 1689.970 141.740 ;
        RECT 2456.470 141.680 2456.790 141.740 ;
        RECT 1689.650 141.540 2456.790 141.680 ;
        RECT 1689.650 141.480 1689.970 141.540 ;
        RECT 2456.470 141.480 2456.790 141.540 ;
        RECT 2456.470 96.460 2456.790 96.520 ;
        RECT 2456.275 96.320 2456.790 96.460 ;
        RECT 2456.470 96.260 2456.790 96.320 ;
        RECT 2456.485 48.520 2456.775 48.565 ;
        RECT 2458.770 48.520 2459.090 48.580 ;
        RECT 2456.485 48.380 2459.090 48.520 ;
        RECT 2456.485 48.335 2456.775 48.380 ;
        RECT 2458.770 48.320 2459.090 48.380 ;
      LAYER via ;
        RECT 1685.540 496.780 1685.800 497.040 ;
        RECT 1689.680 496.780 1689.940 497.040 ;
        RECT 1689.680 141.480 1689.940 141.740 ;
        RECT 2456.500 141.480 2456.760 141.740 ;
        RECT 2456.500 96.260 2456.760 96.520 ;
        RECT 2458.800 48.320 2459.060 48.580 ;
      LAYER met2 ;
        RECT 1685.670 510.340 1685.950 514.000 ;
        RECT 1685.600 510.000 1685.950 510.340 ;
        RECT 1685.600 497.070 1685.740 510.000 ;
        RECT 1685.540 496.750 1685.800 497.070 ;
        RECT 1689.680 496.750 1689.940 497.070 ;
        RECT 1689.740 141.770 1689.880 496.750 ;
        RECT 1689.680 141.450 1689.940 141.770 ;
        RECT 2456.500 141.450 2456.760 141.770 ;
        RECT 2456.560 96.550 2456.700 141.450 ;
        RECT 2456.500 96.230 2456.760 96.550 ;
        RECT 2458.800 48.290 2459.060 48.610 ;
        RECT 2458.860 2.400 2459.000 48.290 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1697.930 496.980 1698.250 497.040 ;
        RECT 1703.910 496.980 1704.230 497.040 ;
        RECT 1697.930 496.840 1704.230 496.980 ;
        RECT 1697.930 496.780 1698.250 496.840 ;
        RECT 1703.910 496.780 1704.230 496.840 ;
        RECT 1703.910 210.700 1704.230 210.760 ;
        RECT 2470.270 210.700 2470.590 210.760 ;
        RECT 1703.910 210.560 2470.590 210.700 ;
        RECT 1703.910 210.500 1704.230 210.560 ;
        RECT 2470.270 210.500 2470.590 210.560 ;
        RECT 2470.270 38.320 2470.590 38.380 ;
        RECT 2476.710 38.320 2477.030 38.380 ;
        RECT 2470.270 38.180 2477.030 38.320 ;
        RECT 2470.270 38.120 2470.590 38.180 ;
        RECT 2476.710 38.120 2477.030 38.180 ;
      LAYER via ;
        RECT 1697.960 496.780 1698.220 497.040 ;
        RECT 1703.940 496.780 1704.200 497.040 ;
        RECT 1703.940 210.500 1704.200 210.760 ;
        RECT 2470.300 210.500 2470.560 210.760 ;
        RECT 2470.300 38.120 2470.560 38.380 ;
        RECT 2476.740 38.120 2477.000 38.380 ;
      LAYER met2 ;
        RECT 1698.090 510.340 1698.370 514.000 ;
        RECT 1698.020 510.000 1698.370 510.340 ;
        RECT 1698.020 497.070 1698.160 510.000 ;
        RECT 1697.960 496.750 1698.220 497.070 ;
        RECT 1703.940 496.750 1704.200 497.070 ;
        RECT 1704.000 210.790 1704.140 496.750 ;
        RECT 1703.940 210.470 1704.200 210.790 ;
        RECT 2470.300 210.470 2470.560 210.790 ;
        RECT 2470.360 38.410 2470.500 210.470 ;
        RECT 2470.300 38.090 2470.560 38.410 ;
        RECT 2476.740 38.090 2477.000 38.410 ;
        RECT 2476.800 2.400 2476.940 38.090 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1710.425 434.945 1710.595 492.915 ;
        RECT 1709.505 282.965 1709.675 331.075 ;
      LAYER mcon ;
        RECT 1710.425 492.745 1710.595 492.915 ;
        RECT 1709.505 330.905 1709.675 331.075 ;
      LAYER met1 ;
        RECT 1710.350 492.900 1710.670 492.960 ;
        RECT 1710.155 492.760 1710.670 492.900 ;
        RECT 1710.350 492.700 1710.670 492.760 ;
        RECT 1710.350 435.100 1710.670 435.160 ;
        RECT 1710.155 434.960 1710.670 435.100 ;
        RECT 1710.350 434.900 1710.670 434.960 ;
        RECT 1708.510 410.280 1708.830 410.340 ;
        RECT 1710.350 410.280 1710.670 410.340 ;
        RECT 1708.510 410.140 1710.670 410.280 ;
        RECT 1708.510 410.080 1708.830 410.140 ;
        RECT 1710.350 410.080 1710.670 410.140 ;
        RECT 1709.890 352.480 1710.210 352.540 ;
        RECT 1709.520 352.340 1710.210 352.480 ;
        RECT 1709.520 351.860 1709.660 352.340 ;
        RECT 1709.890 352.280 1710.210 352.340 ;
        RECT 1709.430 351.600 1709.750 351.860 ;
        RECT 1709.430 331.060 1709.750 331.120 ;
        RECT 1709.235 330.920 1709.750 331.060 ;
        RECT 1709.430 330.860 1709.750 330.920 ;
        RECT 1709.445 283.120 1709.735 283.165 ;
        RECT 1710.350 283.120 1710.670 283.180 ;
        RECT 1709.445 282.980 1710.670 283.120 ;
        RECT 1709.445 282.935 1709.735 282.980 ;
        RECT 1710.350 282.920 1710.670 282.980 ;
        RECT 1710.350 255.380 1710.670 255.640 ;
        RECT 1710.440 254.960 1710.580 255.380 ;
        RECT 1710.350 254.700 1710.670 254.960 ;
        RECT 1710.350 217.500 1710.670 217.560 ;
        RECT 2490.970 217.500 2491.290 217.560 ;
        RECT 1710.350 217.360 2491.290 217.500 ;
        RECT 1710.350 217.300 1710.670 217.360 ;
        RECT 2490.970 217.300 2491.290 217.360 ;
      LAYER via ;
        RECT 1710.380 492.700 1710.640 492.960 ;
        RECT 1710.380 434.900 1710.640 435.160 ;
        RECT 1708.540 410.080 1708.800 410.340 ;
        RECT 1710.380 410.080 1710.640 410.340 ;
        RECT 1709.920 352.280 1710.180 352.540 ;
        RECT 1709.460 351.600 1709.720 351.860 ;
        RECT 1709.460 330.860 1709.720 331.120 ;
        RECT 1710.380 282.920 1710.640 283.180 ;
        RECT 1710.380 255.380 1710.640 255.640 ;
        RECT 1710.380 254.700 1710.640 254.960 ;
        RECT 1710.380 217.300 1710.640 217.560 ;
        RECT 2491.000 217.300 2491.260 217.560 ;
      LAYER met2 ;
        RECT 1710.510 510.340 1710.790 514.000 ;
        RECT 1710.440 510.000 1710.790 510.340 ;
        RECT 1710.440 492.990 1710.580 510.000 ;
        RECT 1710.380 492.670 1710.640 492.990 ;
        RECT 1710.380 434.870 1710.640 435.190 ;
        RECT 1710.440 410.370 1710.580 434.870 ;
        RECT 1708.540 410.050 1708.800 410.370 ;
        RECT 1710.380 410.050 1710.640 410.370 ;
        RECT 1708.600 386.765 1708.740 410.050 ;
        RECT 1708.530 386.395 1708.810 386.765 ;
        RECT 1709.450 386.650 1709.730 386.765 ;
        RECT 1709.450 386.510 1710.120 386.650 ;
        RECT 1709.450 386.395 1709.730 386.510 ;
        RECT 1709.980 352.570 1710.120 386.510 ;
        RECT 1709.920 352.250 1710.180 352.570 ;
        RECT 1709.460 351.570 1709.720 351.890 ;
        RECT 1709.520 339.165 1709.660 351.570 ;
        RECT 1709.450 338.795 1709.730 339.165 ;
        RECT 1709.450 338.115 1709.730 338.485 ;
        RECT 1709.520 331.150 1709.660 338.115 ;
        RECT 1709.460 330.830 1709.720 331.150 ;
        RECT 1710.380 282.890 1710.640 283.210 ;
        RECT 1710.440 255.670 1710.580 282.890 ;
        RECT 1710.380 255.350 1710.640 255.670 ;
        RECT 1710.380 254.670 1710.640 254.990 ;
        RECT 1710.440 217.590 1710.580 254.670 ;
        RECT 1710.380 217.270 1710.640 217.590 ;
        RECT 2491.000 217.270 2491.260 217.590 ;
        RECT 2491.060 17.410 2491.200 217.270 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 1708.530 386.440 1708.810 386.720 ;
        RECT 1709.450 386.440 1709.730 386.720 ;
        RECT 1709.450 338.840 1709.730 339.120 ;
        RECT 1709.450 338.160 1709.730 338.440 ;
      LAYER met3 ;
        RECT 1708.505 386.730 1708.835 386.745 ;
        RECT 1709.425 386.730 1709.755 386.745 ;
        RECT 1708.505 386.430 1709.755 386.730 ;
        RECT 1708.505 386.415 1708.835 386.430 ;
        RECT 1709.425 386.415 1709.755 386.430 ;
        RECT 1709.425 338.815 1709.755 339.145 ;
        RECT 1709.440 338.465 1709.740 338.815 ;
        RECT 1709.425 338.135 1709.755 338.465 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.610 224.640 1724.930 224.700 ;
        RECT 2511.670 224.640 2511.990 224.700 ;
        RECT 1724.610 224.500 2511.990 224.640 ;
        RECT 1724.610 224.440 1724.930 224.500 ;
        RECT 2511.670 224.440 2511.990 224.500 ;
      LAYER via ;
        RECT 1724.640 224.440 1724.900 224.700 ;
        RECT 2511.700 224.440 2511.960 224.700 ;
      LAYER met2 ;
        RECT 1722.930 510.410 1723.210 514.000 ;
        RECT 1722.930 510.270 1724.840 510.410 ;
        RECT 1722.930 510.000 1723.210 510.270 ;
        RECT 1724.700 224.730 1724.840 510.270 ;
        RECT 1724.640 224.410 1724.900 224.730 ;
        RECT 2511.700 224.410 2511.960 224.730 ;
        RECT 2511.760 17.410 2511.900 224.410 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.410 231.440 1738.730 231.500 ;
        RECT 2525.470 231.440 2525.790 231.500 ;
        RECT 1738.410 231.300 2525.790 231.440 ;
        RECT 1738.410 231.240 1738.730 231.300 ;
        RECT 2525.470 231.240 2525.790 231.300 ;
        RECT 2525.470 62.120 2525.790 62.180 ;
        RECT 2530.070 62.120 2530.390 62.180 ;
        RECT 2525.470 61.980 2530.390 62.120 ;
        RECT 2525.470 61.920 2525.790 61.980 ;
        RECT 2530.070 61.920 2530.390 61.980 ;
      LAYER via ;
        RECT 1738.440 231.240 1738.700 231.500 ;
        RECT 2525.500 231.240 2525.760 231.500 ;
        RECT 2525.500 61.920 2525.760 62.180 ;
        RECT 2530.100 61.920 2530.360 62.180 ;
      LAYER met2 ;
        RECT 1735.350 510.410 1735.630 514.000 ;
        RECT 1735.350 510.270 1738.640 510.410 ;
        RECT 1735.350 510.000 1735.630 510.270 ;
        RECT 1738.500 231.530 1738.640 510.270 ;
        RECT 1738.440 231.210 1738.700 231.530 ;
        RECT 2525.500 231.210 2525.760 231.530 ;
        RECT 2525.560 62.210 2525.700 231.210 ;
        RECT 2525.500 61.890 2525.760 62.210 ;
        RECT 2530.100 61.890 2530.360 62.210 ;
        RECT 2530.160 2.400 2530.300 61.890 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2546.245 186.405 2546.415 234.515 ;
        RECT 2546.245 48.365 2546.415 137.955 ;
      LAYER mcon ;
        RECT 2546.245 234.345 2546.415 234.515 ;
        RECT 2546.245 137.785 2546.415 137.955 ;
      LAYER met1 ;
        RECT 1747.610 503.440 1747.930 503.500 ;
        RECT 1751.750 503.440 1752.070 503.500 ;
        RECT 1747.610 503.300 1752.070 503.440 ;
        RECT 1747.610 503.240 1747.930 503.300 ;
        RECT 1751.750 503.240 1752.070 503.300 ;
        RECT 1751.750 238.240 1752.070 238.300 ;
        RECT 2546.170 238.240 2546.490 238.300 ;
        RECT 1751.750 238.100 2546.490 238.240 ;
        RECT 1751.750 238.040 1752.070 238.100 ;
        RECT 2546.170 238.040 2546.490 238.100 ;
        RECT 2546.170 234.500 2546.490 234.560 ;
        RECT 2545.975 234.360 2546.490 234.500 ;
        RECT 2546.170 234.300 2546.490 234.360 ;
        RECT 2546.170 186.560 2546.490 186.620 ;
        RECT 2545.975 186.420 2546.490 186.560 ;
        RECT 2546.170 186.360 2546.490 186.420 ;
        RECT 2546.170 137.940 2546.490 138.000 ;
        RECT 2545.975 137.800 2546.490 137.940 ;
        RECT 2546.170 137.740 2546.490 137.800 ;
        RECT 2546.185 48.520 2546.475 48.565 ;
        RECT 2548.010 48.520 2548.330 48.580 ;
        RECT 2546.185 48.380 2548.330 48.520 ;
        RECT 2546.185 48.335 2546.475 48.380 ;
        RECT 2548.010 48.320 2548.330 48.380 ;
      LAYER via ;
        RECT 1747.640 503.240 1747.900 503.500 ;
        RECT 1751.780 503.240 1752.040 503.500 ;
        RECT 1751.780 238.040 1752.040 238.300 ;
        RECT 2546.200 238.040 2546.460 238.300 ;
        RECT 2546.200 234.300 2546.460 234.560 ;
        RECT 2546.200 186.360 2546.460 186.620 ;
        RECT 2546.200 137.740 2546.460 138.000 ;
        RECT 2548.040 48.320 2548.300 48.580 ;
      LAYER met2 ;
        RECT 1747.770 510.340 1748.050 514.000 ;
        RECT 1747.700 510.000 1748.050 510.340 ;
        RECT 1747.700 503.530 1747.840 510.000 ;
        RECT 1747.640 503.210 1747.900 503.530 ;
        RECT 1751.780 503.210 1752.040 503.530 ;
        RECT 1751.840 238.330 1751.980 503.210 ;
        RECT 1751.780 238.010 1752.040 238.330 ;
        RECT 2546.200 238.010 2546.460 238.330 ;
        RECT 2546.260 234.590 2546.400 238.010 ;
        RECT 2546.200 234.270 2546.460 234.590 ;
        RECT 2546.200 186.330 2546.460 186.650 ;
        RECT 2546.260 138.030 2546.400 186.330 ;
        RECT 2546.200 137.710 2546.460 138.030 ;
        RECT 2548.040 48.290 2548.300 48.610 ;
        RECT 2548.100 2.400 2548.240 48.290 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1760.030 496.980 1760.350 497.040 ;
        RECT 1765.550 496.980 1765.870 497.040 ;
        RECT 1760.030 496.840 1765.870 496.980 ;
        RECT 1760.030 496.780 1760.350 496.840 ;
        RECT 1765.550 496.780 1765.870 496.840 ;
        RECT 1765.550 245.380 1765.870 245.440 ;
        RECT 2559.970 245.380 2560.290 245.440 ;
        RECT 1765.550 245.240 2560.290 245.380 ;
        RECT 1765.550 245.180 1765.870 245.240 ;
        RECT 2559.970 245.180 2560.290 245.240 ;
        RECT 2559.970 38.320 2560.290 38.380 ;
        RECT 2565.950 38.320 2566.270 38.380 ;
        RECT 2559.970 38.180 2566.270 38.320 ;
        RECT 2559.970 38.120 2560.290 38.180 ;
        RECT 2565.950 38.120 2566.270 38.180 ;
      LAYER via ;
        RECT 1760.060 496.780 1760.320 497.040 ;
        RECT 1765.580 496.780 1765.840 497.040 ;
        RECT 1765.580 245.180 1765.840 245.440 ;
        RECT 2560.000 245.180 2560.260 245.440 ;
        RECT 2560.000 38.120 2560.260 38.380 ;
        RECT 2565.980 38.120 2566.240 38.380 ;
      LAYER met2 ;
        RECT 1760.190 510.340 1760.470 514.000 ;
        RECT 1760.120 510.000 1760.470 510.340 ;
        RECT 1760.120 497.070 1760.260 510.000 ;
        RECT 1760.060 496.750 1760.320 497.070 ;
        RECT 1765.580 496.750 1765.840 497.070 ;
        RECT 1765.640 245.470 1765.780 496.750 ;
        RECT 1765.580 245.150 1765.840 245.470 ;
        RECT 2560.000 245.150 2560.260 245.470 ;
        RECT 2560.060 38.410 2560.200 245.150 ;
        RECT 2560.000 38.090 2560.260 38.410 ;
        RECT 2565.980 38.090 2566.240 38.410 ;
        RECT 2566.040 2.400 2566.180 38.090 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2580.745 48.365 2580.915 96.475 ;
      LAYER mcon ;
        RECT 2580.745 96.305 2580.915 96.475 ;
      LAYER met1 ;
        RECT 1772.910 155.620 1773.230 155.680 ;
        RECT 2580.670 155.620 2580.990 155.680 ;
        RECT 1772.910 155.480 2580.990 155.620 ;
        RECT 1772.910 155.420 1773.230 155.480 ;
        RECT 2580.670 155.420 2580.990 155.480 ;
        RECT 2580.670 96.460 2580.990 96.520 ;
        RECT 2580.475 96.320 2580.990 96.460 ;
        RECT 2580.670 96.260 2580.990 96.320 ;
        RECT 2580.685 48.520 2580.975 48.565 ;
        RECT 2583.890 48.520 2584.210 48.580 ;
        RECT 2580.685 48.380 2584.210 48.520 ;
        RECT 2580.685 48.335 2580.975 48.380 ;
        RECT 2583.890 48.320 2584.210 48.380 ;
      LAYER via ;
        RECT 1772.940 155.420 1773.200 155.680 ;
        RECT 2580.700 155.420 2580.960 155.680 ;
        RECT 2580.700 96.260 2580.960 96.520 ;
        RECT 2583.920 48.320 2584.180 48.580 ;
      LAYER met2 ;
        RECT 1772.610 510.340 1772.890 514.000 ;
        RECT 1772.540 510.000 1772.890 510.340 ;
        RECT 1772.540 497.490 1772.680 510.000 ;
        RECT 1772.540 497.350 1773.140 497.490 ;
        RECT 1773.000 155.710 1773.140 497.350 ;
        RECT 1772.940 155.390 1773.200 155.710 ;
        RECT 2580.700 155.390 2580.960 155.710 ;
        RECT 2580.760 96.550 2580.900 155.390 ;
        RECT 2580.700 96.230 2580.960 96.550 ;
        RECT 2583.920 48.290 2584.180 48.610 ;
        RECT 2583.980 2.400 2584.120 48.290 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 547.470 496.980 547.790 497.040 ;
        RECT 555.290 496.980 555.610 497.040 ;
        RECT 547.470 496.840 555.610 496.980 ;
        RECT 547.470 496.780 547.790 496.840 ;
        RECT 555.290 496.780 555.610 496.840 ;
        RECT 555.290 155.280 555.610 155.340 ;
        RECT 814.270 155.280 814.590 155.340 ;
        RECT 555.290 155.140 814.590 155.280 ;
        RECT 555.290 155.080 555.610 155.140 ;
        RECT 814.270 155.080 814.590 155.140 ;
      LAYER via ;
        RECT 547.500 496.780 547.760 497.040 ;
        RECT 555.320 496.780 555.580 497.040 ;
        RECT 555.320 155.080 555.580 155.340 ;
        RECT 814.300 155.080 814.560 155.340 ;
      LAYER met2 ;
        RECT 547.630 510.340 547.910 514.000 ;
        RECT 547.560 510.000 547.910 510.340 ;
        RECT 547.560 497.070 547.700 510.000 ;
        RECT 547.500 496.750 547.760 497.070 ;
        RECT 555.320 496.750 555.580 497.070 ;
        RECT 555.380 155.370 555.520 496.750 ;
        RECT 555.320 155.050 555.580 155.370 ;
        RECT 814.300 155.050 814.560 155.370 ;
        RECT 814.360 17.410 814.500 155.050 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.710 162.420 1787.030 162.480 ;
        RECT 2601.370 162.420 2601.690 162.480 ;
        RECT 1786.710 162.280 2601.690 162.420 ;
        RECT 1786.710 162.220 1787.030 162.280 ;
        RECT 2601.370 162.220 2601.690 162.280 ;
      LAYER via ;
        RECT 1786.740 162.220 1787.000 162.480 ;
        RECT 2601.400 162.220 2601.660 162.480 ;
      LAYER met2 ;
        RECT 1784.570 510.410 1784.850 514.000 ;
        RECT 1784.570 510.270 1786.940 510.410 ;
        RECT 1784.570 510.000 1784.850 510.270 ;
        RECT 1786.800 162.510 1786.940 510.270 ;
        RECT 1786.740 162.190 1787.000 162.510 ;
        RECT 2601.400 162.190 2601.660 162.510 ;
        RECT 2601.460 2.400 2601.600 162.190 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1796.830 496.980 1797.150 497.040 ;
        RECT 1800.510 496.980 1800.830 497.040 ;
        RECT 1796.830 496.840 1800.830 496.980 ;
        RECT 1796.830 496.780 1797.150 496.840 ;
        RECT 1800.510 496.780 1800.830 496.840 ;
        RECT 1800.510 169.220 1800.830 169.280 ;
        RECT 2615.170 169.220 2615.490 169.280 ;
        RECT 1800.510 169.080 2615.490 169.220 ;
        RECT 1800.510 169.020 1800.830 169.080 ;
        RECT 2615.170 169.020 2615.490 169.080 ;
        RECT 2615.170 62.120 2615.490 62.180 ;
        RECT 2619.310 62.120 2619.630 62.180 ;
        RECT 2615.170 61.980 2619.630 62.120 ;
        RECT 2615.170 61.920 2615.490 61.980 ;
        RECT 2619.310 61.920 2619.630 61.980 ;
      LAYER via ;
        RECT 1796.860 496.780 1797.120 497.040 ;
        RECT 1800.540 496.780 1800.800 497.040 ;
        RECT 1800.540 169.020 1800.800 169.280 ;
        RECT 2615.200 169.020 2615.460 169.280 ;
        RECT 2615.200 61.920 2615.460 62.180 ;
        RECT 2619.340 61.920 2619.600 62.180 ;
      LAYER met2 ;
        RECT 1796.990 510.340 1797.270 514.000 ;
        RECT 1796.920 510.000 1797.270 510.340 ;
        RECT 1796.920 497.070 1797.060 510.000 ;
        RECT 1796.860 496.750 1797.120 497.070 ;
        RECT 1800.540 496.750 1800.800 497.070 ;
        RECT 1800.600 169.310 1800.740 496.750 ;
        RECT 1800.540 168.990 1800.800 169.310 ;
        RECT 2615.200 168.990 2615.460 169.310 ;
        RECT 2615.260 62.210 2615.400 168.990 ;
        RECT 2615.200 61.890 2615.460 62.210 ;
        RECT 2619.340 61.890 2619.600 62.210 ;
        RECT 2619.400 2.400 2619.540 61.890 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2635.945 186.405 2636.115 234.515 ;
        RECT 2635.945 89.845 2636.115 137.955 ;
      LAYER mcon ;
        RECT 2635.945 234.345 2636.115 234.515 ;
        RECT 2635.945 137.785 2636.115 137.955 ;
      LAYER met1 ;
        RECT 1809.250 496.980 1809.570 497.040 ;
        RECT 1813.850 496.980 1814.170 497.040 ;
        RECT 1809.250 496.840 1814.170 496.980 ;
        RECT 1809.250 496.780 1809.570 496.840 ;
        RECT 1813.850 496.780 1814.170 496.840 ;
        RECT 1813.850 252.180 1814.170 252.240 ;
        RECT 2635.870 252.180 2636.190 252.240 ;
        RECT 1813.850 252.040 2636.190 252.180 ;
        RECT 1813.850 251.980 1814.170 252.040 ;
        RECT 2635.870 251.980 2636.190 252.040 ;
        RECT 2635.870 234.500 2636.190 234.560 ;
        RECT 2635.675 234.360 2636.190 234.500 ;
        RECT 2635.870 234.300 2636.190 234.360 ;
        RECT 2635.870 186.560 2636.190 186.620 ;
        RECT 2635.675 186.420 2636.190 186.560 ;
        RECT 2635.870 186.360 2636.190 186.420 ;
        RECT 2635.870 137.940 2636.190 138.000 ;
        RECT 2635.675 137.800 2636.190 137.940 ;
        RECT 2635.870 137.740 2636.190 137.800 ;
        RECT 2635.870 90.000 2636.190 90.060 ;
        RECT 2635.675 89.860 2636.190 90.000 ;
        RECT 2635.870 89.800 2636.190 89.860 ;
        RECT 2635.870 74.360 2636.190 74.420 ;
        RECT 2636.790 74.360 2637.110 74.420 ;
        RECT 2635.870 74.220 2637.110 74.360 ;
        RECT 2635.870 74.160 2636.190 74.220 ;
        RECT 2636.790 74.160 2637.110 74.220 ;
        RECT 2637.250 47.980 2637.570 48.240 ;
        RECT 2637.340 47.560 2637.480 47.980 ;
        RECT 2637.250 47.300 2637.570 47.560 ;
      LAYER via ;
        RECT 1809.280 496.780 1809.540 497.040 ;
        RECT 1813.880 496.780 1814.140 497.040 ;
        RECT 1813.880 251.980 1814.140 252.240 ;
        RECT 2635.900 251.980 2636.160 252.240 ;
        RECT 2635.900 234.300 2636.160 234.560 ;
        RECT 2635.900 186.360 2636.160 186.620 ;
        RECT 2635.900 137.740 2636.160 138.000 ;
        RECT 2635.900 89.800 2636.160 90.060 ;
        RECT 2635.900 74.160 2636.160 74.420 ;
        RECT 2636.820 74.160 2637.080 74.420 ;
        RECT 2637.280 47.980 2637.540 48.240 ;
        RECT 2637.280 47.300 2637.540 47.560 ;
      LAYER met2 ;
        RECT 1809.410 510.340 1809.690 514.000 ;
        RECT 1809.340 510.000 1809.690 510.340 ;
        RECT 1809.340 497.070 1809.480 510.000 ;
        RECT 1809.280 496.750 1809.540 497.070 ;
        RECT 1813.880 496.750 1814.140 497.070 ;
        RECT 1813.940 252.270 1814.080 496.750 ;
        RECT 1813.880 251.950 1814.140 252.270 ;
        RECT 2635.900 251.950 2636.160 252.270 ;
        RECT 2635.960 234.590 2636.100 251.950 ;
        RECT 2635.900 234.270 2636.160 234.590 ;
        RECT 2635.900 186.330 2636.160 186.650 ;
        RECT 2635.960 138.030 2636.100 186.330 ;
        RECT 2635.900 137.710 2636.160 138.030 ;
        RECT 2635.900 89.770 2636.160 90.090 ;
        RECT 2635.960 74.450 2636.100 89.770 ;
        RECT 2635.900 74.130 2636.160 74.450 ;
        RECT 2636.820 74.130 2637.080 74.450 ;
        RECT 2636.880 61.610 2637.020 74.130 ;
        RECT 2636.880 61.470 2637.480 61.610 ;
        RECT 2637.340 48.270 2637.480 61.470 ;
        RECT 2637.280 47.950 2637.540 48.270 ;
        RECT 2637.280 47.270 2637.540 47.590 ;
        RECT 2637.340 2.400 2637.480 47.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1821.670 497.320 1821.990 497.380 ;
        RECT 1838.690 497.320 1839.010 497.380 ;
        RECT 1821.670 497.180 1839.010 497.320 ;
        RECT 1821.670 497.120 1821.990 497.180 ;
        RECT 1838.690 497.120 1839.010 497.180 ;
        RECT 1838.690 258.640 1839.010 258.700 ;
        RECT 2649.670 258.640 2649.990 258.700 ;
        RECT 1838.690 258.500 2649.990 258.640 ;
        RECT 1838.690 258.440 1839.010 258.500 ;
        RECT 2649.670 258.440 2649.990 258.500 ;
        RECT 2649.670 62.120 2649.990 62.180 ;
        RECT 2655.190 62.120 2655.510 62.180 ;
        RECT 2649.670 61.980 2655.510 62.120 ;
        RECT 2649.670 61.920 2649.990 61.980 ;
        RECT 2655.190 61.920 2655.510 61.980 ;
      LAYER via ;
        RECT 1821.700 497.120 1821.960 497.380 ;
        RECT 1838.720 497.120 1838.980 497.380 ;
        RECT 1838.720 258.440 1838.980 258.700 ;
        RECT 2649.700 258.440 2649.960 258.700 ;
        RECT 2649.700 61.920 2649.960 62.180 ;
        RECT 2655.220 61.920 2655.480 62.180 ;
      LAYER met2 ;
        RECT 1821.830 510.340 1822.110 514.000 ;
        RECT 1821.760 510.000 1822.110 510.340 ;
        RECT 1821.760 497.410 1821.900 510.000 ;
        RECT 1821.700 497.090 1821.960 497.410 ;
        RECT 1838.720 497.090 1838.980 497.410 ;
        RECT 1838.780 258.730 1838.920 497.090 ;
        RECT 1838.720 258.410 1838.980 258.730 ;
        RECT 2649.700 258.410 2649.960 258.730 ;
        RECT 2649.760 62.210 2649.900 258.410 ;
        RECT 2649.700 61.890 2649.960 62.210 ;
        RECT 2655.220 61.890 2655.480 62.210 ;
        RECT 2655.280 2.400 2655.420 61.890 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 265.440 1835.330 265.500 ;
        RECT 2670.370 265.440 2670.690 265.500 ;
        RECT 1835.010 265.300 2670.690 265.440 ;
        RECT 1835.010 265.240 1835.330 265.300 ;
        RECT 2670.370 265.240 2670.690 265.300 ;
      LAYER via ;
        RECT 1835.040 265.240 1835.300 265.500 ;
        RECT 2670.400 265.240 2670.660 265.500 ;
      LAYER met2 ;
        RECT 1834.250 510.410 1834.530 514.000 ;
        RECT 1834.250 510.270 1835.240 510.410 ;
        RECT 1834.250 510.000 1834.530 510.270 ;
        RECT 1835.100 265.530 1835.240 510.270 ;
        RECT 1835.040 265.210 1835.300 265.530 ;
        RECT 2670.400 265.210 2670.660 265.530 ;
        RECT 2670.460 17.410 2670.600 265.210 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.810 272.580 1849.130 272.640 ;
        RECT 2684.630 272.580 2684.950 272.640 ;
        RECT 1848.810 272.440 2684.950 272.580 ;
        RECT 1848.810 272.380 1849.130 272.440 ;
        RECT 2684.630 272.380 2684.950 272.440 ;
        RECT 2684.630 17.920 2684.950 17.980 ;
        RECT 2690.610 17.920 2690.930 17.980 ;
        RECT 2684.630 17.780 2690.930 17.920 ;
        RECT 2684.630 17.720 2684.950 17.780 ;
        RECT 2690.610 17.720 2690.930 17.780 ;
      LAYER via ;
        RECT 1848.840 272.380 1849.100 272.640 ;
        RECT 2684.660 272.380 2684.920 272.640 ;
        RECT 2684.660 17.720 2684.920 17.980 ;
        RECT 2690.640 17.720 2690.900 17.980 ;
      LAYER met2 ;
        RECT 1846.670 510.410 1846.950 514.000 ;
        RECT 1846.670 510.270 1849.040 510.410 ;
        RECT 1846.670 510.000 1846.950 510.270 ;
        RECT 1848.900 272.670 1849.040 510.270 ;
        RECT 1848.840 272.350 1849.100 272.670 ;
        RECT 2684.660 272.350 2684.920 272.670 ;
        RECT 2684.720 18.010 2684.860 272.350 ;
        RECT 2684.660 17.690 2684.920 18.010 ;
        RECT 2690.640 17.690 2690.900 18.010 ;
        RECT 2690.700 2.400 2690.840 17.690 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1862.610 176.020 1862.930 176.080 ;
        RECT 2704.870 176.020 2705.190 176.080 ;
        RECT 1862.610 175.880 2705.190 176.020 ;
        RECT 1862.610 175.820 1862.930 175.880 ;
        RECT 2704.870 175.820 2705.190 175.880 ;
      LAYER via ;
        RECT 1862.640 175.820 1862.900 176.080 ;
        RECT 2704.900 175.820 2705.160 176.080 ;
      LAYER met2 ;
        RECT 1859.090 510.410 1859.370 514.000 ;
        RECT 1859.090 510.270 1862.840 510.410 ;
        RECT 1859.090 510.000 1859.370 510.270 ;
        RECT 1862.700 176.110 1862.840 510.270 ;
        RECT 1862.640 175.790 1862.900 176.110 ;
        RECT 2704.900 175.790 2705.160 176.110 ;
        RECT 2704.960 16.730 2705.100 175.790 ;
        RECT 2704.960 16.590 2708.780 16.730 ;
        RECT 2708.640 2.400 2708.780 16.590 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2726.565 2.805 2726.735 48.195 ;
      LAYER mcon ;
        RECT 2726.565 48.025 2726.735 48.195 ;
      LAYER met1 ;
        RECT 1871.350 503.440 1871.670 503.500 ;
        RECT 1875.950 503.440 1876.270 503.500 ;
        RECT 1871.350 503.300 1876.270 503.440 ;
        RECT 1871.350 503.240 1871.670 503.300 ;
        RECT 1875.950 503.240 1876.270 503.300 ;
        RECT 1875.950 362.340 1876.270 362.400 ;
        RECT 2725.570 362.340 2725.890 362.400 ;
        RECT 1875.950 362.200 2725.890 362.340 ;
        RECT 1875.950 362.140 1876.270 362.200 ;
        RECT 2725.570 362.140 2725.890 362.200 ;
        RECT 2725.570 62.260 2725.890 62.520 ;
        RECT 2725.660 61.780 2725.800 62.260 ;
        RECT 2726.490 61.780 2726.810 61.840 ;
        RECT 2725.660 61.640 2726.810 61.780 ;
        RECT 2726.490 61.580 2726.810 61.640 ;
        RECT 2726.490 48.180 2726.810 48.240 ;
        RECT 2726.295 48.040 2726.810 48.180 ;
        RECT 2726.490 47.980 2726.810 48.040 ;
        RECT 2726.490 2.960 2726.810 3.020 ;
        RECT 2726.295 2.820 2726.810 2.960 ;
        RECT 2726.490 2.760 2726.810 2.820 ;
      LAYER via ;
        RECT 1871.380 503.240 1871.640 503.500 ;
        RECT 1875.980 503.240 1876.240 503.500 ;
        RECT 1875.980 362.140 1876.240 362.400 ;
        RECT 2725.600 362.140 2725.860 362.400 ;
        RECT 2725.600 62.260 2725.860 62.520 ;
        RECT 2726.520 61.580 2726.780 61.840 ;
        RECT 2726.520 47.980 2726.780 48.240 ;
        RECT 2726.520 2.760 2726.780 3.020 ;
      LAYER met2 ;
        RECT 1871.510 510.340 1871.790 514.000 ;
        RECT 1871.440 510.000 1871.790 510.340 ;
        RECT 1871.440 503.530 1871.580 510.000 ;
        RECT 1871.380 503.210 1871.640 503.530 ;
        RECT 1875.980 503.210 1876.240 503.530 ;
        RECT 1876.040 362.430 1876.180 503.210 ;
        RECT 1875.980 362.110 1876.240 362.430 ;
        RECT 2725.600 362.110 2725.860 362.430 ;
        RECT 2725.660 62.550 2725.800 362.110 ;
        RECT 2725.600 62.230 2725.860 62.550 ;
        RECT 2726.520 61.550 2726.780 61.870 ;
        RECT 2726.580 48.270 2726.720 61.550 ;
        RECT 2726.520 47.950 2726.780 48.270 ;
        RECT 2726.520 2.730 2726.780 3.050 ;
        RECT 2726.580 2.400 2726.720 2.730 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2744.505 2.805 2744.675 48.195 ;
      LAYER mcon ;
        RECT 2744.505 48.025 2744.675 48.195 ;
      LAYER met1 ;
        RECT 1883.770 499.360 1884.090 499.420 ;
        RECT 1889.750 499.360 1890.070 499.420 ;
        RECT 1883.770 499.220 1890.070 499.360 ;
        RECT 1883.770 499.160 1884.090 499.220 ;
        RECT 1889.750 499.160 1890.070 499.220 ;
        RECT 1889.750 355.200 1890.070 355.260 ;
        RECT 2739.370 355.200 2739.690 355.260 ;
        RECT 1889.750 355.060 2739.690 355.200 ;
        RECT 1889.750 355.000 1890.070 355.060 ;
        RECT 2739.370 355.000 2739.690 355.060 ;
        RECT 2739.370 96.460 2739.690 96.520 ;
        RECT 2744.430 96.460 2744.750 96.520 ;
        RECT 2739.370 96.320 2744.750 96.460 ;
        RECT 2739.370 96.260 2739.690 96.320 ;
        RECT 2744.430 96.260 2744.750 96.320 ;
        RECT 2744.430 48.180 2744.750 48.240 ;
        RECT 2744.235 48.040 2744.750 48.180 ;
        RECT 2744.430 47.980 2744.750 48.040 ;
        RECT 2744.430 2.960 2744.750 3.020 ;
        RECT 2744.235 2.820 2744.750 2.960 ;
        RECT 2744.430 2.760 2744.750 2.820 ;
      LAYER via ;
        RECT 1883.800 499.160 1884.060 499.420 ;
        RECT 1889.780 499.160 1890.040 499.420 ;
        RECT 1889.780 355.000 1890.040 355.260 ;
        RECT 2739.400 355.000 2739.660 355.260 ;
        RECT 2739.400 96.260 2739.660 96.520 ;
        RECT 2744.460 96.260 2744.720 96.520 ;
        RECT 2744.460 47.980 2744.720 48.240 ;
        RECT 2744.460 2.760 2744.720 3.020 ;
      LAYER met2 ;
        RECT 1883.930 510.340 1884.210 514.000 ;
        RECT 1883.860 510.000 1884.210 510.340 ;
        RECT 1883.860 499.450 1884.000 510.000 ;
        RECT 1883.800 499.130 1884.060 499.450 ;
        RECT 1889.780 499.130 1890.040 499.450 ;
        RECT 1889.840 355.290 1889.980 499.130 ;
        RECT 1889.780 354.970 1890.040 355.290 ;
        RECT 2739.400 354.970 2739.660 355.290 ;
        RECT 2739.460 96.550 2739.600 354.970 ;
        RECT 2739.400 96.230 2739.660 96.550 ;
        RECT 2744.460 96.230 2744.720 96.550 ;
        RECT 2744.520 48.270 2744.660 96.230 ;
        RECT 2744.460 47.950 2744.720 48.270 ;
        RECT 2744.460 2.730 2744.720 3.050 ;
        RECT 2744.520 2.400 2744.660 2.730 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1895.730 501.060 1896.050 501.120 ;
        RECT 2018.090 501.060 2018.410 501.120 ;
        RECT 1895.730 500.920 2018.410 501.060 ;
        RECT 1895.730 500.860 1896.050 500.920 ;
        RECT 2018.090 500.860 2018.410 500.920 ;
        RECT 2018.090 279.380 2018.410 279.440 ;
        RECT 2760.070 279.380 2760.390 279.440 ;
        RECT 2018.090 279.240 2760.390 279.380 ;
        RECT 2018.090 279.180 2018.410 279.240 ;
        RECT 2760.070 279.180 2760.390 279.240 ;
        RECT 2760.530 61.780 2760.850 61.840 ;
        RECT 2761.910 61.780 2762.230 61.840 ;
        RECT 2760.530 61.640 2762.230 61.780 ;
        RECT 2760.530 61.580 2760.850 61.640 ;
        RECT 2761.910 61.580 2762.230 61.640 ;
      LAYER via ;
        RECT 1895.760 500.860 1896.020 501.120 ;
        RECT 2018.120 500.860 2018.380 501.120 ;
        RECT 2018.120 279.180 2018.380 279.440 ;
        RECT 2760.100 279.180 2760.360 279.440 ;
        RECT 2760.560 61.580 2760.820 61.840 ;
        RECT 2761.940 61.580 2762.200 61.840 ;
      LAYER met2 ;
        RECT 1895.890 510.340 1896.170 514.000 ;
        RECT 1895.820 510.000 1896.170 510.340 ;
        RECT 1895.820 501.150 1895.960 510.000 ;
        RECT 1895.760 500.830 1896.020 501.150 ;
        RECT 2018.120 500.830 2018.380 501.150 ;
        RECT 2018.180 279.470 2018.320 500.830 ;
        RECT 2018.120 279.150 2018.380 279.470 ;
        RECT 2760.100 279.150 2760.360 279.470 ;
        RECT 2760.160 72.490 2760.300 279.150 ;
        RECT 2760.160 72.350 2760.760 72.490 ;
        RECT 2760.620 61.870 2760.760 72.350 ;
        RECT 2760.560 61.550 2760.820 61.870 ;
        RECT 2761.940 61.550 2762.200 61.870 ;
        RECT 2762.000 2.400 2762.140 61.550 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 559.890 496.980 560.210 497.040 ;
        RECT 575.990 496.980 576.310 497.040 ;
        RECT 559.890 496.840 576.310 496.980 ;
        RECT 559.890 496.780 560.210 496.840 ;
        RECT 575.990 496.780 576.310 496.840 ;
        RECT 575.990 162.080 576.310 162.140 ;
        RECT 835.430 162.080 835.750 162.140 ;
        RECT 575.990 161.940 835.750 162.080 ;
        RECT 575.990 161.880 576.310 161.940 ;
        RECT 835.430 161.880 835.750 161.940 ;
      LAYER via ;
        RECT 559.920 496.780 560.180 497.040 ;
        RECT 576.020 496.780 576.280 497.040 ;
        RECT 576.020 161.880 576.280 162.140 ;
        RECT 835.460 161.880 835.720 162.140 ;
      LAYER met2 ;
        RECT 560.050 510.340 560.330 514.000 ;
        RECT 559.980 510.000 560.330 510.340 ;
        RECT 559.980 497.070 560.120 510.000 ;
        RECT 559.920 496.750 560.180 497.070 ;
        RECT 576.020 496.750 576.280 497.070 ;
        RECT 576.080 162.170 576.220 496.750 ;
        RECT 576.020 161.850 576.280 162.170 ;
        RECT 835.460 161.850 835.720 162.170 ;
        RECT 835.520 2.400 835.660 161.850 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.910 348.400 1911.230 348.460 ;
        RECT 2773.870 348.400 2774.190 348.460 ;
        RECT 1910.910 348.260 2774.190 348.400 ;
        RECT 1910.910 348.200 1911.230 348.260 ;
        RECT 2773.870 348.200 2774.190 348.260 ;
        RECT 2773.870 37.980 2774.190 38.040 ;
        RECT 2779.850 37.980 2780.170 38.040 ;
        RECT 2773.870 37.840 2780.170 37.980 ;
        RECT 2773.870 37.780 2774.190 37.840 ;
        RECT 2779.850 37.780 2780.170 37.840 ;
      LAYER via ;
        RECT 1910.940 348.200 1911.200 348.460 ;
        RECT 2773.900 348.200 2774.160 348.460 ;
        RECT 2773.900 37.780 2774.160 38.040 ;
        RECT 2779.880 37.780 2780.140 38.040 ;
      LAYER met2 ;
        RECT 1908.310 510.410 1908.590 514.000 ;
        RECT 1908.310 510.270 1911.140 510.410 ;
        RECT 1908.310 510.000 1908.590 510.270 ;
        RECT 1911.000 348.490 1911.140 510.270 ;
        RECT 1910.940 348.170 1911.200 348.490 ;
        RECT 2773.900 348.170 2774.160 348.490 ;
        RECT 2773.960 38.070 2774.100 348.170 ;
        RECT 2773.900 37.750 2774.160 38.070 ;
        RECT 2779.880 37.750 2780.140 38.070 ;
        RECT 2779.940 2.400 2780.080 37.750 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1920.570 500.040 1920.890 500.100 ;
        RECT 2466.590 500.040 2466.910 500.100 ;
        RECT 1920.570 499.900 2466.910 500.040 ;
        RECT 1920.570 499.840 1920.890 499.900 ;
        RECT 2466.590 499.840 2466.910 499.900 ;
        RECT 2466.590 24.040 2466.910 24.100 ;
        RECT 2797.790 24.040 2798.110 24.100 ;
        RECT 2466.590 23.900 2798.110 24.040 ;
        RECT 2466.590 23.840 2466.910 23.900 ;
        RECT 2797.790 23.840 2798.110 23.900 ;
      LAYER via ;
        RECT 1920.600 499.840 1920.860 500.100 ;
        RECT 2466.620 499.840 2466.880 500.100 ;
        RECT 2466.620 23.840 2466.880 24.100 ;
        RECT 2797.820 23.840 2798.080 24.100 ;
      LAYER met2 ;
        RECT 1920.730 510.340 1921.010 514.000 ;
        RECT 1920.660 510.000 1921.010 510.340 ;
        RECT 1920.660 500.130 1920.800 510.000 ;
        RECT 1920.600 499.810 1920.860 500.130 ;
        RECT 2466.620 499.810 2466.880 500.130 ;
        RECT 2466.680 24.130 2466.820 499.810 ;
        RECT 2466.620 23.810 2466.880 24.130 ;
        RECT 2797.820 23.810 2798.080 24.130 ;
        RECT 2797.880 2.400 2798.020 23.810 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1932.990 496.980 1933.310 497.040 ;
        RECT 1938.050 496.980 1938.370 497.040 ;
        RECT 1932.990 496.840 1938.370 496.980 ;
        RECT 1932.990 496.780 1933.310 496.840 ;
        RECT 1938.050 496.780 1938.370 496.840 ;
        RECT 1938.050 341.600 1938.370 341.660 ;
        RECT 2815.270 341.600 2815.590 341.660 ;
        RECT 1938.050 341.460 2815.590 341.600 ;
        RECT 1938.050 341.400 1938.370 341.460 ;
        RECT 2815.270 341.400 2815.590 341.460 ;
      LAYER via ;
        RECT 1933.020 496.780 1933.280 497.040 ;
        RECT 1938.080 496.780 1938.340 497.040 ;
        RECT 1938.080 341.400 1938.340 341.660 ;
        RECT 2815.300 341.400 2815.560 341.660 ;
      LAYER met2 ;
        RECT 1933.150 510.340 1933.430 514.000 ;
        RECT 1933.080 510.000 1933.430 510.340 ;
        RECT 1933.080 497.070 1933.220 510.000 ;
        RECT 1933.020 496.750 1933.280 497.070 ;
        RECT 1938.080 496.750 1938.340 497.070 ;
        RECT 1938.140 341.690 1938.280 496.750 ;
        RECT 1938.080 341.370 1938.340 341.690 ;
        RECT 2815.300 341.370 2815.560 341.690 ;
        RECT 2815.360 37.130 2815.500 341.370 ;
        RECT 2815.360 36.990 2815.960 37.130 ;
        RECT 2815.820 2.400 2815.960 36.990 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1945.410 334.460 1945.730 334.520 ;
        RECT 2829.070 334.460 2829.390 334.520 ;
        RECT 1945.410 334.320 2829.390 334.460 ;
        RECT 1945.410 334.260 1945.730 334.320 ;
        RECT 2829.070 334.260 2829.390 334.320 ;
        RECT 2829.070 62.120 2829.390 62.180 ;
        RECT 2833.670 62.120 2833.990 62.180 ;
        RECT 2829.070 61.980 2833.990 62.120 ;
        RECT 2829.070 61.920 2829.390 61.980 ;
        RECT 2833.670 61.920 2833.990 61.980 ;
      LAYER via ;
        RECT 1945.440 334.260 1945.700 334.520 ;
        RECT 2829.100 334.260 2829.360 334.520 ;
        RECT 2829.100 61.920 2829.360 62.180 ;
        RECT 2833.700 61.920 2833.960 62.180 ;
      LAYER met2 ;
        RECT 1945.570 510.340 1945.850 514.000 ;
        RECT 1945.500 510.000 1945.850 510.340 ;
        RECT 1945.500 334.550 1945.640 510.000 ;
        RECT 1945.440 334.230 1945.700 334.550 ;
        RECT 2829.100 334.230 2829.360 334.550 ;
        RECT 2829.160 62.210 2829.300 334.230 ;
        RECT 2829.100 61.890 2829.360 62.210 ;
        RECT 2833.700 61.890 2833.960 62.210 ;
        RECT 2833.760 2.400 2833.900 61.890 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2849.845 282.965 2850.015 327.675 ;
        RECT 2849.845 186.405 2850.015 234.515 ;
        RECT 2849.845 48.365 2850.015 137.955 ;
      LAYER mcon ;
        RECT 2849.845 327.505 2850.015 327.675 ;
        RECT 2849.845 234.345 2850.015 234.515 ;
        RECT 2849.845 137.785 2850.015 137.955 ;
      LAYER met1 ;
        RECT 1959.210 327.660 1959.530 327.720 ;
        RECT 2849.785 327.660 2850.075 327.705 ;
        RECT 1959.210 327.520 2850.075 327.660 ;
        RECT 1959.210 327.460 1959.530 327.520 ;
        RECT 2849.785 327.475 2850.075 327.520 ;
        RECT 2849.770 283.120 2850.090 283.180 ;
        RECT 2849.575 282.980 2850.090 283.120 ;
        RECT 2849.770 282.920 2850.090 282.980 ;
        RECT 2849.770 234.500 2850.090 234.560 ;
        RECT 2849.575 234.360 2850.090 234.500 ;
        RECT 2849.770 234.300 2850.090 234.360 ;
        RECT 2849.770 186.560 2850.090 186.620 ;
        RECT 2849.575 186.420 2850.090 186.560 ;
        RECT 2849.770 186.360 2850.090 186.420 ;
        RECT 2849.770 137.940 2850.090 138.000 ;
        RECT 2849.575 137.800 2850.090 137.940 ;
        RECT 2849.770 137.740 2850.090 137.800 ;
        RECT 2849.785 48.520 2850.075 48.565 ;
        RECT 2851.150 48.520 2851.470 48.580 ;
        RECT 2849.785 48.380 2851.470 48.520 ;
        RECT 2849.785 48.335 2850.075 48.380 ;
        RECT 2851.150 48.320 2851.470 48.380 ;
      LAYER via ;
        RECT 1959.240 327.460 1959.500 327.720 ;
        RECT 2849.800 282.920 2850.060 283.180 ;
        RECT 2849.800 234.300 2850.060 234.560 ;
        RECT 2849.800 186.360 2850.060 186.620 ;
        RECT 2849.800 137.740 2850.060 138.000 ;
        RECT 2851.180 48.320 2851.440 48.580 ;
      LAYER met2 ;
        RECT 1957.990 510.410 1958.270 514.000 ;
        RECT 1957.990 510.270 1959.440 510.410 ;
        RECT 1957.990 510.000 1958.270 510.270 ;
        RECT 1959.300 327.750 1959.440 510.270 ;
        RECT 1959.240 327.430 1959.500 327.750 ;
        RECT 2849.800 282.890 2850.060 283.210 ;
        RECT 2849.860 234.590 2850.000 282.890 ;
        RECT 2849.800 234.270 2850.060 234.590 ;
        RECT 2849.800 186.330 2850.060 186.650 ;
        RECT 2849.860 138.030 2850.000 186.330 ;
        RECT 2849.800 137.710 2850.060 138.030 ;
        RECT 2851.180 48.290 2851.440 48.610 ;
        RECT 2851.240 2.400 2851.380 48.290 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 286.180 1973.330 286.240 ;
        RECT 2863.570 286.180 2863.890 286.240 ;
        RECT 1973.010 286.040 2863.890 286.180 ;
        RECT 1973.010 285.980 1973.330 286.040 ;
        RECT 2863.570 285.980 2863.890 286.040 ;
      LAYER via ;
        RECT 1973.040 285.980 1973.300 286.240 ;
        RECT 2863.600 285.980 2863.860 286.240 ;
      LAYER met2 ;
        RECT 1970.410 510.410 1970.690 514.000 ;
        RECT 1970.410 510.270 1973.240 510.410 ;
        RECT 1970.410 510.000 1970.690 510.270 ;
        RECT 1973.100 286.270 1973.240 510.270 ;
        RECT 1973.040 285.950 1973.300 286.270 ;
        RECT 2863.600 285.950 2863.860 286.270 ;
        RECT 2863.660 18.090 2863.800 285.950 ;
        RECT 2863.660 17.950 2869.320 18.090 ;
        RECT 2869.180 2.400 2869.320 17.950 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1982.670 496.980 1982.990 497.040 ;
        RECT 1990.490 496.980 1990.810 497.040 ;
        RECT 1982.670 496.840 1990.810 496.980 ;
        RECT 1982.670 496.780 1982.990 496.840 ;
        RECT 1990.490 496.780 1990.810 496.840 ;
        RECT 1990.490 320.860 1990.810 320.920 ;
        RECT 2884.270 320.860 2884.590 320.920 ;
        RECT 1990.490 320.720 2884.590 320.860 ;
        RECT 1990.490 320.660 1990.810 320.720 ;
        RECT 2884.270 320.660 2884.590 320.720 ;
        RECT 2884.270 2.960 2884.590 3.020 ;
        RECT 2887.030 2.960 2887.350 3.020 ;
        RECT 2884.270 2.820 2887.350 2.960 ;
        RECT 2884.270 2.760 2884.590 2.820 ;
        RECT 2887.030 2.760 2887.350 2.820 ;
      LAYER via ;
        RECT 1982.700 496.780 1982.960 497.040 ;
        RECT 1990.520 496.780 1990.780 497.040 ;
        RECT 1990.520 320.660 1990.780 320.920 ;
        RECT 2884.300 320.660 2884.560 320.920 ;
        RECT 2884.300 2.760 2884.560 3.020 ;
        RECT 2887.060 2.760 2887.320 3.020 ;
      LAYER met2 ;
        RECT 1982.830 510.340 1983.110 514.000 ;
        RECT 1982.760 510.000 1983.110 510.340 ;
        RECT 1982.760 497.070 1982.900 510.000 ;
        RECT 1982.700 496.750 1982.960 497.070 ;
        RECT 1990.520 496.750 1990.780 497.070 ;
        RECT 1990.580 320.950 1990.720 496.750 ;
        RECT 1990.520 320.630 1990.780 320.950 ;
        RECT 2884.300 320.630 2884.560 320.950 ;
        RECT 2884.360 3.050 2884.500 320.630 ;
        RECT 2884.300 2.730 2884.560 3.050 ;
        RECT 2887.060 2.730 2887.320 3.050 ;
        RECT 2887.120 2.400 2887.260 2.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 496.980 1995.410 497.040 ;
        RECT 2000.610 496.980 2000.930 497.040 ;
        RECT 1995.090 496.840 2000.930 496.980 ;
        RECT 1995.090 496.780 1995.410 496.840 ;
        RECT 2000.610 496.780 2000.930 496.840 ;
        RECT 2000.610 314.060 2000.930 314.120 ;
        RECT 2894.390 314.060 2894.710 314.120 ;
        RECT 2000.610 313.920 2894.710 314.060 ;
        RECT 2000.610 313.860 2000.930 313.920 ;
        RECT 2894.390 313.860 2894.710 313.920 ;
        RECT 2894.390 15.880 2894.710 15.940 ;
        RECT 2904.970 15.880 2905.290 15.940 ;
        RECT 2894.390 15.740 2905.290 15.880 ;
        RECT 2894.390 15.680 2894.710 15.740 ;
        RECT 2904.970 15.680 2905.290 15.740 ;
      LAYER via ;
        RECT 1995.120 496.780 1995.380 497.040 ;
        RECT 2000.640 496.780 2000.900 497.040 ;
        RECT 2000.640 313.860 2000.900 314.120 ;
        RECT 2894.420 313.860 2894.680 314.120 ;
        RECT 2894.420 15.680 2894.680 15.940 ;
        RECT 2905.000 15.680 2905.260 15.940 ;
      LAYER met2 ;
        RECT 1995.250 510.340 1995.530 514.000 ;
        RECT 1995.180 510.000 1995.530 510.340 ;
        RECT 1995.180 497.070 1995.320 510.000 ;
        RECT 1995.120 496.750 1995.380 497.070 ;
        RECT 2000.640 496.750 2000.900 497.070 ;
        RECT 2000.700 314.150 2000.840 496.750 ;
        RECT 2000.640 313.830 2000.900 314.150 ;
        RECT 2894.420 313.830 2894.680 314.150 ;
        RECT 2894.480 15.970 2894.620 313.830 ;
        RECT 2894.420 15.650 2894.680 15.970 ;
        RECT 2905.000 15.650 2905.260 15.970 ;
        RECT 2905.060 2.400 2905.200 15.650 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 572.310 168.880 572.630 168.940 ;
        RECT 848.770 168.880 849.090 168.940 ;
        RECT 572.310 168.740 849.090 168.880 ;
        RECT 572.310 168.680 572.630 168.740 ;
        RECT 848.770 168.680 849.090 168.740 ;
      LAYER via ;
        RECT 572.340 168.680 572.600 168.940 ;
        RECT 848.800 168.680 849.060 168.940 ;
      LAYER met2 ;
        RECT 572.470 510.340 572.750 514.000 ;
        RECT 572.400 510.000 572.750 510.340 ;
        RECT 572.400 168.970 572.540 510.000 ;
        RECT 572.340 168.650 572.600 168.970 ;
        RECT 848.800 168.650 849.060 168.970 ;
        RECT 848.860 17.410 849.000 168.650 ;
        RECT 848.860 17.270 853.140 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 585.650 176.020 585.970 176.080 ;
        RECT 869.470 176.020 869.790 176.080 ;
        RECT 585.650 175.880 869.790 176.020 ;
        RECT 585.650 175.820 585.970 175.880 ;
        RECT 869.470 175.820 869.790 175.880 ;
      LAYER via ;
        RECT 585.680 175.820 585.940 176.080 ;
        RECT 869.500 175.820 869.760 176.080 ;
      LAYER met2 ;
        RECT 584.890 510.410 585.170 514.000 ;
        RECT 584.890 510.270 585.880 510.410 ;
        RECT 584.890 510.000 585.170 510.270 ;
        RECT 585.740 176.110 585.880 510.270 ;
        RECT 585.680 175.790 585.940 176.110 ;
        RECT 869.500 175.790 869.760 176.110 ;
        RECT 869.560 17.410 869.700 175.790 ;
        RECT 869.560 17.270 871.080 17.410 ;
        RECT 870.940 2.400 871.080 17.270 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 599.910 182.820 600.230 182.880 ;
        RECT 883.270 182.820 883.590 182.880 ;
        RECT 599.910 182.680 883.590 182.820 ;
        RECT 599.910 182.620 600.230 182.680 ;
        RECT 883.270 182.620 883.590 182.680 ;
      LAYER via ;
        RECT 599.940 182.620 600.200 182.880 ;
        RECT 883.300 182.620 883.560 182.880 ;
      LAYER met2 ;
        RECT 597.310 510.410 597.590 514.000 ;
        RECT 597.310 510.270 600.140 510.410 ;
        RECT 597.310 510.000 597.590 510.270 ;
        RECT 600.000 182.910 600.140 510.270 ;
        RECT 599.940 182.590 600.200 182.910 ;
        RECT 883.300 182.590 883.560 182.910 ;
        RECT 883.360 17.410 883.500 182.590 ;
        RECT 883.360 17.270 889.020 17.410 ;
        RECT 888.880 2.400 889.020 17.270 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.570 496.980 609.890 497.040 ;
        RECT 613.710 496.980 614.030 497.040 ;
        RECT 609.570 496.840 614.030 496.980 ;
        RECT 609.570 496.780 609.890 496.840 ;
        RECT 613.710 496.780 614.030 496.840 ;
        RECT 613.710 189.620 614.030 189.680 ;
        RECT 903.970 189.620 904.290 189.680 ;
        RECT 613.710 189.480 904.290 189.620 ;
        RECT 613.710 189.420 614.030 189.480 ;
        RECT 903.970 189.420 904.290 189.480 ;
      LAYER via ;
        RECT 609.600 496.780 609.860 497.040 ;
        RECT 613.740 496.780 614.000 497.040 ;
        RECT 613.740 189.420 614.000 189.680 ;
        RECT 904.000 189.420 904.260 189.680 ;
      LAYER met2 ;
        RECT 609.730 510.340 610.010 514.000 ;
        RECT 609.660 510.000 610.010 510.340 ;
        RECT 609.660 497.070 609.800 510.000 ;
        RECT 609.600 496.750 609.860 497.070 ;
        RECT 613.740 496.750 614.000 497.070 ;
        RECT 613.800 189.710 613.940 496.750 ;
        RECT 613.740 189.390 614.000 189.710 ;
        RECT 904.000 189.390 904.260 189.710 ;
        RECT 904.060 17.410 904.200 189.390 ;
        RECT 904.060 17.270 906.960 17.410 ;
        RECT 906.820 2.400 906.960 17.270 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 621.990 496.980 622.310 497.040 ;
        RECT 627.510 496.980 627.830 497.040 ;
        RECT 621.990 496.840 627.830 496.980 ;
        RECT 621.990 496.780 622.310 496.840 ;
        RECT 627.510 496.780 627.830 496.840 ;
        RECT 627.510 24.040 627.830 24.100 ;
        RECT 724.570 24.040 724.890 24.100 ;
        RECT 627.510 23.900 724.890 24.040 ;
        RECT 627.510 23.840 627.830 23.900 ;
        RECT 724.570 23.840 724.890 23.900 ;
        RECT 725.030 24.040 725.350 24.100 ;
        RECT 924.210 24.040 924.530 24.100 ;
        RECT 725.030 23.900 924.530 24.040 ;
        RECT 725.030 23.840 725.350 23.900 ;
        RECT 924.210 23.840 924.530 23.900 ;
      LAYER via ;
        RECT 622.020 496.780 622.280 497.040 ;
        RECT 627.540 496.780 627.800 497.040 ;
        RECT 627.540 23.840 627.800 24.100 ;
        RECT 724.600 23.840 724.860 24.100 ;
        RECT 725.060 23.840 725.320 24.100 ;
        RECT 924.240 23.840 924.500 24.100 ;
      LAYER met2 ;
        RECT 622.150 510.340 622.430 514.000 ;
        RECT 622.080 510.000 622.430 510.340 ;
        RECT 622.080 497.070 622.220 510.000 ;
        RECT 622.020 496.750 622.280 497.070 ;
        RECT 627.540 496.750 627.800 497.070 ;
        RECT 627.600 24.130 627.740 496.750 ;
        RECT 627.540 23.810 627.800 24.130 ;
        RECT 724.600 23.810 724.860 24.130 ;
        RECT 725.060 23.810 725.320 24.130 ;
        RECT 924.240 23.810 924.500 24.130 ;
        RECT 724.660 23.530 724.800 23.810 ;
        RECT 725.120 23.530 725.260 23.810 ;
        RECT 724.660 23.390 725.260 23.530 ;
        RECT 924.300 2.400 924.440 23.810 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 633.950 196.760 634.270 196.820 ;
        RECT 938.470 196.760 938.790 196.820 ;
        RECT 633.950 196.620 938.790 196.760 ;
        RECT 633.950 196.560 634.270 196.620 ;
        RECT 938.470 196.560 938.790 196.620 ;
      LAYER via ;
        RECT 633.980 196.560 634.240 196.820 ;
        RECT 938.500 196.560 938.760 196.820 ;
      LAYER met2 ;
        RECT 634.570 510.410 634.850 514.000 ;
        RECT 634.040 510.270 634.850 510.410 ;
        RECT 634.040 196.850 634.180 510.270 ;
        RECT 634.570 510.000 634.850 510.270 ;
        RECT 633.980 196.530 634.240 196.850 ;
        RECT 938.500 196.530 938.760 196.850 ;
        RECT 938.560 17.410 938.700 196.530 ;
        RECT 938.560 17.270 942.380 17.410 ;
        RECT 942.240 2.400 942.380 17.270 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 647.750 203.560 648.070 203.620 ;
        RECT 959.170 203.560 959.490 203.620 ;
        RECT 647.750 203.420 959.490 203.560 ;
        RECT 647.750 203.360 648.070 203.420 ;
        RECT 959.170 203.360 959.490 203.420 ;
      LAYER via ;
        RECT 647.780 203.360 648.040 203.620 ;
        RECT 959.200 203.360 959.460 203.620 ;
      LAYER met2 ;
        RECT 646.530 510.410 646.810 514.000 ;
        RECT 646.530 510.270 647.980 510.410 ;
        RECT 646.530 510.000 646.810 510.270 ;
        RECT 647.840 203.650 647.980 510.270 ;
        RECT 647.780 203.330 648.040 203.650 ;
        RECT 959.200 203.330 959.460 203.650 ;
        RECT 959.260 17.410 959.400 203.330 ;
        RECT 959.260 17.270 960.320 17.410 ;
        RECT 960.180 2.400 960.320 17.270 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 210.700 662.330 210.760 ;
        RECT 972.970 210.700 973.290 210.760 ;
        RECT 662.010 210.560 973.290 210.700 ;
        RECT 662.010 210.500 662.330 210.560 ;
        RECT 972.970 210.500 973.290 210.560 ;
      LAYER via ;
        RECT 662.040 210.500 662.300 210.760 ;
        RECT 973.000 210.500 973.260 210.760 ;
      LAYER met2 ;
        RECT 658.950 510.410 659.230 514.000 ;
        RECT 658.950 510.270 662.240 510.410 ;
        RECT 658.950 510.000 659.230 510.270 ;
        RECT 662.100 210.790 662.240 510.270 ;
        RECT 662.040 210.470 662.300 210.790 ;
        RECT 973.000 210.470 973.260 210.790 ;
        RECT 973.060 17.410 973.200 210.470 ;
        RECT 973.060 17.270 978.260 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 436.150 497.320 436.470 497.380 ;
        RECT 444.890 497.320 445.210 497.380 ;
        RECT 436.150 497.180 445.210 497.320 ;
        RECT 436.150 497.120 436.470 497.180 ;
        RECT 444.890 497.120 445.210 497.180 ;
        RECT 444.890 107.000 445.210 107.060 ;
        RECT 655.570 107.000 655.890 107.060 ;
        RECT 444.890 106.860 655.890 107.000 ;
        RECT 444.890 106.800 445.210 106.860 ;
        RECT 655.570 106.800 655.890 106.860 ;
        RECT 655.570 2.960 655.890 3.020 ;
        RECT 656.950 2.960 657.270 3.020 ;
        RECT 655.570 2.820 657.270 2.960 ;
        RECT 655.570 2.760 655.890 2.820 ;
        RECT 656.950 2.760 657.270 2.820 ;
      LAYER via ;
        RECT 436.180 497.120 436.440 497.380 ;
        RECT 444.920 497.120 445.180 497.380 ;
        RECT 444.920 106.800 445.180 107.060 ;
        RECT 655.600 106.800 655.860 107.060 ;
        RECT 655.600 2.760 655.860 3.020 ;
        RECT 656.980 2.760 657.240 3.020 ;
      LAYER met2 ;
        RECT 436.310 510.340 436.590 514.000 ;
        RECT 436.240 510.000 436.590 510.340 ;
        RECT 436.240 497.410 436.380 510.000 ;
        RECT 436.180 497.090 436.440 497.410 ;
        RECT 444.920 497.090 445.180 497.410 ;
        RECT 444.980 107.090 445.120 497.090 ;
        RECT 444.920 106.770 445.180 107.090 ;
        RECT 655.600 106.770 655.860 107.090 ;
        RECT 655.660 3.050 655.800 106.770 ;
        RECT 655.600 2.730 655.860 3.050 ;
        RECT 656.980 2.730 657.240 3.050 ;
        RECT 657.040 2.400 657.180 2.730 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 993.745 48.365 993.915 137.275 ;
      LAYER mcon ;
        RECT 993.745 137.105 993.915 137.275 ;
      LAYER met1 ;
        RECT 671.210 496.980 671.530 497.040 ;
        RECT 675.810 496.980 676.130 497.040 ;
        RECT 671.210 496.840 676.130 496.980 ;
        RECT 671.210 496.780 671.530 496.840 ;
        RECT 675.810 496.780 676.130 496.840 ;
        RECT 675.810 217.160 676.130 217.220 ;
        RECT 993.670 217.160 993.990 217.220 ;
        RECT 675.810 217.020 993.990 217.160 ;
        RECT 675.810 216.960 676.130 217.020 ;
        RECT 993.670 216.960 993.990 217.020 ;
        RECT 992.750 193.020 993.070 193.080 ;
        RECT 993.670 193.020 993.990 193.080 ;
        RECT 992.750 192.880 993.990 193.020 ;
        RECT 992.750 192.820 993.070 192.880 ;
        RECT 993.670 192.820 993.990 192.880 ;
        RECT 993.670 137.740 993.990 138.000 ;
        RECT 993.760 137.305 993.900 137.740 ;
        RECT 993.685 137.075 993.975 137.305 ;
        RECT 993.685 48.520 993.975 48.565 ;
        RECT 995.970 48.520 996.290 48.580 ;
        RECT 993.685 48.380 996.290 48.520 ;
        RECT 993.685 48.335 993.975 48.380 ;
        RECT 995.970 48.320 996.290 48.380 ;
      LAYER via ;
        RECT 671.240 496.780 671.500 497.040 ;
        RECT 675.840 496.780 676.100 497.040 ;
        RECT 675.840 216.960 676.100 217.220 ;
        RECT 993.700 216.960 993.960 217.220 ;
        RECT 992.780 192.820 993.040 193.080 ;
        RECT 993.700 192.820 993.960 193.080 ;
        RECT 993.700 137.740 993.960 138.000 ;
        RECT 996.000 48.320 996.260 48.580 ;
      LAYER met2 ;
        RECT 671.370 510.340 671.650 514.000 ;
        RECT 671.300 510.000 671.650 510.340 ;
        RECT 671.300 497.070 671.440 510.000 ;
        RECT 671.240 496.750 671.500 497.070 ;
        RECT 675.840 496.750 676.100 497.070 ;
        RECT 675.900 217.250 676.040 496.750 ;
        RECT 675.840 216.930 676.100 217.250 ;
        RECT 993.700 216.930 993.960 217.250 ;
        RECT 993.760 193.110 993.900 216.930 ;
        RECT 992.780 192.790 993.040 193.110 ;
        RECT 993.700 192.790 993.960 193.110 ;
        RECT 992.840 145.365 992.980 192.790 ;
        RECT 992.770 144.995 993.050 145.365 ;
        RECT 993.690 144.995 993.970 145.365 ;
        RECT 993.760 138.030 993.900 144.995 ;
        RECT 993.700 137.710 993.960 138.030 ;
        RECT 996.000 48.290 996.260 48.610 ;
        RECT 996.060 2.400 996.200 48.290 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 992.770 145.040 993.050 145.320 ;
        RECT 993.690 145.040 993.970 145.320 ;
      LAYER met3 ;
        RECT 992.745 145.330 993.075 145.345 ;
        RECT 993.665 145.330 993.995 145.345 ;
        RECT 992.745 145.030 993.995 145.330 ;
        RECT 992.745 145.015 993.075 145.030 ;
        RECT 993.665 145.015 993.995 145.030 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 683.630 496.980 683.950 497.040 ;
        RECT 689.610 496.980 689.930 497.040 ;
        RECT 683.630 496.840 689.930 496.980 ;
        RECT 683.630 496.780 683.950 496.840 ;
        RECT 689.610 496.780 689.930 496.840 ;
        RECT 689.610 231.440 689.930 231.500 ;
        RECT 1007.470 231.440 1007.790 231.500 ;
        RECT 689.610 231.300 1007.790 231.440 ;
        RECT 689.610 231.240 689.930 231.300 ;
        RECT 1007.470 231.240 1007.790 231.300 ;
        RECT 1007.470 37.980 1007.790 38.040 ;
        RECT 1013.450 37.980 1013.770 38.040 ;
        RECT 1007.470 37.840 1013.770 37.980 ;
        RECT 1007.470 37.780 1007.790 37.840 ;
        RECT 1013.450 37.780 1013.770 37.840 ;
      LAYER via ;
        RECT 683.660 496.780 683.920 497.040 ;
        RECT 689.640 496.780 689.900 497.040 ;
        RECT 689.640 231.240 689.900 231.500 ;
        RECT 1007.500 231.240 1007.760 231.500 ;
        RECT 1007.500 37.780 1007.760 38.040 ;
        RECT 1013.480 37.780 1013.740 38.040 ;
      LAYER met2 ;
        RECT 683.790 510.340 684.070 514.000 ;
        RECT 683.720 510.000 684.070 510.340 ;
        RECT 683.720 497.070 683.860 510.000 ;
        RECT 683.660 496.750 683.920 497.070 ;
        RECT 689.640 496.750 689.900 497.070 ;
        RECT 689.700 231.530 689.840 496.750 ;
        RECT 689.640 231.210 689.900 231.530 ;
        RECT 1007.500 231.210 1007.760 231.530 ;
        RECT 1007.560 38.070 1007.700 231.210 ;
        RECT 1007.500 37.750 1007.760 38.070 ;
        RECT 1013.480 37.750 1013.740 38.070 ;
        RECT 1013.540 2.400 1013.680 37.750 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.050 237.900 696.370 237.960 ;
        RECT 1028.170 237.900 1028.490 237.960 ;
        RECT 696.050 237.760 1028.490 237.900 ;
        RECT 696.050 237.700 696.370 237.760 ;
        RECT 1028.170 237.700 1028.490 237.760 ;
      LAYER via ;
        RECT 696.080 237.700 696.340 237.960 ;
        RECT 1028.200 237.700 1028.460 237.960 ;
      LAYER met2 ;
        RECT 696.210 510.340 696.490 514.000 ;
        RECT 696.140 510.000 696.490 510.340 ;
        RECT 696.140 237.990 696.280 510.000 ;
        RECT 696.080 237.670 696.340 237.990 ;
        RECT 1028.200 237.670 1028.460 237.990 ;
        RECT 1028.260 16.730 1028.400 237.670 ;
        RECT 1028.260 16.590 1031.620 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 245.040 710.170 245.100 ;
        RECT 1049.330 245.040 1049.650 245.100 ;
        RECT 709.850 244.900 1049.650 245.040 ;
        RECT 709.850 244.840 710.170 244.900 ;
        RECT 1049.330 244.840 1049.650 244.900 ;
      LAYER via ;
        RECT 709.880 244.840 710.140 245.100 ;
        RECT 1049.360 244.840 1049.620 245.100 ;
      LAYER met2 ;
        RECT 708.630 510.410 708.910 514.000 ;
        RECT 708.630 510.270 710.080 510.410 ;
        RECT 708.630 510.000 708.910 510.270 ;
        RECT 709.940 245.130 710.080 510.270 ;
        RECT 709.880 244.810 710.140 245.130 ;
        RECT 1049.360 244.810 1049.620 245.130 ;
        RECT 1049.420 2.400 1049.560 244.810 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 724.110 252.180 724.430 252.240 ;
        RECT 1062.670 252.180 1062.990 252.240 ;
        RECT 724.110 252.040 1062.990 252.180 ;
        RECT 724.110 251.980 724.430 252.040 ;
        RECT 1062.670 251.980 1062.990 252.040 ;
      LAYER via ;
        RECT 724.140 251.980 724.400 252.240 ;
        RECT 1062.700 251.980 1062.960 252.240 ;
      LAYER met2 ;
        RECT 721.050 510.410 721.330 514.000 ;
        RECT 721.050 510.270 724.340 510.410 ;
        RECT 721.050 510.000 721.330 510.270 ;
        RECT 724.200 252.270 724.340 510.270 ;
        RECT 724.140 251.950 724.400 252.270 ;
        RECT 1062.700 251.950 1062.960 252.270 ;
        RECT 1062.760 17.410 1062.900 251.950 ;
        RECT 1062.760 17.270 1067.500 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 733.310 496.980 733.630 497.040 ;
        RECT 737.910 496.980 738.230 497.040 ;
        RECT 733.310 496.840 738.230 496.980 ;
        RECT 733.310 496.780 733.630 496.840 ;
        RECT 737.910 496.780 738.230 496.840 ;
        RECT 737.910 258.640 738.230 258.700 ;
        RECT 1083.370 258.640 1083.690 258.700 ;
        RECT 737.910 258.500 1083.690 258.640 ;
        RECT 737.910 258.440 738.230 258.500 ;
        RECT 1083.370 258.440 1083.690 258.500 ;
      LAYER via ;
        RECT 733.340 496.780 733.600 497.040 ;
        RECT 737.940 496.780 738.200 497.040 ;
        RECT 737.940 258.440 738.200 258.700 ;
        RECT 1083.400 258.440 1083.660 258.700 ;
      LAYER met2 ;
        RECT 733.470 510.340 733.750 514.000 ;
        RECT 733.400 510.000 733.750 510.340 ;
        RECT 733.400 497.070 733.540 510.000 ;
        RECT 733.340 496.750 733.600 497.070 ;
        RECT 737.940 496.750 738.200 497.070 ;
        RECT 738.000 258.730 738.140 496.750 ;
        RECT 737.940 258.410 738.200 258.730 ;
        RECT 1083.400 258.410 1083.660 258.730 ;
        RECT 1083.460 17.410 1083.600 258.410 ;
        RECT 1083.460 17.270 1085.440 17.410 ;
        RECT 1085.300 2.400 1085.440 17.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 745.730 498.680 746.050 498.740 ;
        RECT 751.710 498.680 752.030 498.740 ;
        RECT 745.730 498.540 752.030 498.680 ;
        RECT 745.730 498.480 746.050 498.540 ;
        RECT 751.710 498.480 752.030 498.540 ;
        RECT 751.710 265.440 752.030 265.500 ;
        RECT 1097.170 265.440 1097.490 265.500 ;
        RECT 751.710 265.300 1097.490 265.440 ;
        RECT 751.710 265.240 752.030 265.300 ;
        RECT 1097.170 265.240 1097.490 265.300 ;
      LAYER via ;
        RECT 745.760 498.480 746.020 498.740 ;
        RECT 751.740 498.480 752.000 498.740 ;
        RECT 751.740 265.240 752.000 265.500 ;
        RECT 1097.200 265.240 1097.460 265.500 ;
      LAYER met2 ;
        RECT 745.890 510.340 746.170 514.000 ;
        RECT 745.820 510.000 746.170 510.340 ;
        RECT 745.820 498.770 745.960 510.000 ;
        RECT 745.760 498.450 746.020 498.770 ;
        RECT 751.740 498.450 752.000 498.770 ;
        RECT 751.800 265.530 751.940 498.450 ;
        RECT 751.740 265.210 752.000 265.530 ;
        RECT 1097.200 265.210 1097.460 265.530 ;
        RECT 1097.260 17.410 1097.400 265.210 ;
        RECT 1097.260 17.270 1102.920 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 757.765 338.045 757.935 386.155 ;
      LAYER mcon ;
        RECT 757.765 385.985 757.935 386.155 ;
      LAYER met1 ;
        RECT 757.230 448.700 757.550 448.760 ;
        RECT 758.150 448.700 758.470 448.760 ;
        RECT 757.230 448.560 758.470 448.700 ;
        RECT 757.230 448.500 757.550 448.560 ;
        RECT 758.150 448.500 758.470 448.560 ;
        RECT 757.690 386.140 758.010 386.200 ;
        RECT 757.495 386.000 758.010 386.140 ;
        RECT 757.690 385.940 758.010 386.000 ;
        RECT 757.705 338.200 757.995 338.245 ;
        RECT 758.150 338.200 758.470 338.260 ;
        RECT 757.705 338.060 758.470 338.200 ;
        RECT 757.705 338.015 757.995 338.060 ;
        RECT 758.150 338.000 758.470 338.060 ;
        RECT 757.230 337.520 757.550 337.580 ;
        RECT 758.150 337.520 758.470 337.580 ;
        RECT 757.230 337.380 758.470 337.520 ;
        RECT 757.230 337.320 757.550 337.380 ;
        RECT 758.150 337.320 758.470 337.380 ;
        RECT 757.230 272.920 757.550 272.980 ;
        RECT 1117.870 272.920 1118.190 272.980 ;
        RECT 757.230 272.780 1118.190 272.920 ;
        RECT 757.230 272.720 757.550 272.780 ;
        RECT 1117.870 272.720 1118.190 272.780 ;
      LAYER via ;
        RECT 757.260 448.500 757.520 448.760 ;
        RECT 758.180 448.500 758.440 448.760 ;
        RECT 757.720 385.940 757.980 386.200 ;
        RECT 758.180 338.000 758.440 338.260 ;
        RECT 757.260 337.320 757.520 337.580 ;
        RECT 758.180 337.320 758.440 337.580 ;
        RECT 757.260 272.720 757.520 272.980 ;
        RECT 1117.900 272.720 1118.160 272.980 ;
      LAYER met2 ;
        RECT 757.850 510.410 758.130 514.000 ;
        RECT 757.320 510.270 758.130 510.410 ;
        RECT 757.320 483.325 757.460 510.270 ;
        RECT 757.850 510.000 758.130 510.270 ;
        RECT 757.250 482.955 757.530 483.325 ;
        RECT 758.170 482.955 758.450 483.325 ;
        RECT 758.240 448.790 758.380 482.955 ;
        RECT 757.260 448.530 757.520 448.790 ;
        RECT 758.180 448.530 758.440 448.790 ;
        RECT 757.260 448.470 758.440 448.530 ;
        RECT 757.320 448.390 758.380 448.470 ;
        RECT 758.240 401.045 758.380 448.390 ;
        RECT 758.170 400.675 758.450 401.045 ;
        RECT 757.710 386.395 757.990 386.765 ;
        RECT 757.780 386.230 757.920 386.395 ;
        RECT 757.720 385.910 757.980 386.230 ;
        RECT 758.180 337.970 758.440 338.290 ;
        RECT 758.240 337.610 758.380 337.970 ;
        RECT 757.260 337.290 757.520 337.610 ;
        RECT 758.180 337.290 758.440 337.610 ;
        RECT 757.320 273.010 757.460 337.290 ;
        RECT 757.260 272.690 757.520 273.010 ;
        RECT 1117.900 272.690 1118.160 273.010 ;
        RECT 1117.960 17.410 1118.100 272.690 ;
        RECT 1117.960 17.270 1120.860 17.410 ;
        RECT 1120.720 2.400 1120.860 17.270 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 757.250 483.000 757.530 483.280 ;
        RECT 758.170 483.000 758.450 483.280 ;
        RECT 758.170 400.720 758.450 401.000 ;
        RECT 757.710 386.440 757.990 386.720 ;
      LAYER met3 ;
        RECT 757.225 483.290 757.555 483.305 ;
        RECT 758.145 483.290 758.475 483.305 ;
        RECT 757.225 482.990 758.475 483.290 ;
        RECT 757.225 482.975 757.555 482.990 ;
        RECT 758.145 482.975 758.475 482.990 ;
        RECT 757.430 401.010 757.810 401.020 ;
        RECT 758.145 401.010 758.475 401.025 ;
        RECT 757.430 400.710 758.475 401.010 ;
        RECT 757.430 400.700 757.810 400.710 ;
        RECT 758.145 400.695 758.475 400.710 ;
        RECT 757.685 386.740 758.015 386.745 ;
        RECT 757.430 386.730 758.015 386.740 ;
        RECT 757.430 386.430 758.240 386.730 ;
        RECT 757.430 386.420 758.015 386.430 ;
        RECT 757.685 386.415 758.015 386.420 ;
      LAYER via3 ;
        RECT 757.460 400.700 757.780 401.020 ;
        RECT 757.460 386.420 757.780 386.740 ;
      LAYER met4 ;
        RECT 757.455 400.695 757.785 401.025 ;
        RECT 757.470 386.745 757.770 400.695 ;
        RECT 757.455 386.415 757.785 386.745 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 771.950 279.380 772.270 279.440 ;
        RECT 1139.030 279.380 1139.350 279.440 ;
        RECT 771.950 279.240 1139.350 279.380 ;
        RECT 771.950 279.180 772.270 279.240 ;
        RECT 1139.030 279.180 1139.350 279.240 ;
      LAYER via ;
        RECT 771.980 279.180 772.240 279.440 ;
        RECT 1139.060 279.180 1139.320 279.440 ;
      LAYER met2 ;
        RECT 770.270 510.410 770.550 514.000 ;
        RECT 770.270 510.270 772.180 510.410 ;
        RECT 770.270 510.000 770.550 510.270 ;
        RECT 772.040 279.470 772.180 510.270 ;
        RECT 771.980 279.150 772.240 279.470 ;
        RECT 1139.060 279.150 1139.320 279.470 ;
        RECT 1139.120 17.410 1139.260 279.150 ;
        RECT 1138.660 17.270 1139.260 17.410 ;
        RECT 1138.660 2.400 1138.800 17.270 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 286.180 786.530 286.240 ;
        RECT 1152.370 286.180 1152.690 286.240 ;
        RECT 786.210 286.040 1152.690 286.180 ;
        RECT 786.210 285.980 786.530 286.040 ;
        RECT 1152.370 285.980 1152.690 286.040 ;
      LAYER via ;
        RECT 786.240 285.980 786.500 286.240 ;
        RECT 1152.400 285.980 1152.660 286.240 ;
      LAYER met2 ;
        RECT 782.690 510.410 782.970 514.000 ;
        RECT 782.690 510.270 786.440 510.410 ;
        RECT 782.690 510.000 782.970 510.270 ;
        RECT 786.300 286.270 786.440 510.270 ;
        RECT 786.240 285.950 786.500 286.270 ;
        RECT 1152.400 285.950 1152.660 286.270 ;
        RECT 1152.460 17.410 1152.600 285.950 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 503.440 448.890 503.500 ;
        RECT 454.550 503.440 454.870 503.500 ;
        RECT 448.570 503.300 454.870 503.440 ;
        RECT 448.570 503.240 448.890 503.300 ;
        RECT 454.550 503.240 454.870 503.300 ;
        RECT 454.550 141.340 454.870 141.400 ;
        RECT 669.370 141.340 669.690 141.400 ;
        RECT 454.550 141.200 669.690 141.340 ;
        RECT 454.550 141.140 454.870 141.200 ;
        RECT 669.370 141.140 669.690 141.200 ;
        RECT 669.370 62.120 669.690 62.180 ;
        RECT 673.970 62.120 674.290 62.180 ;
        RECT 669.370 61.980 674.290 62.120 ;
        RECT 669.370 61.920 669.690 61.980 ;
        RECT 673.970 61.920 674.290 61.980 ;
      LAYER via ;
        RECT 448.600 503.240 448.860 503.500 ;
        RECT 454.580 503.240 454.840 503.500 ;
        RECT 454.580 141.140 454.840 141.400 ;
        RECT 669.400 141.140 669.660 141.400 ;
        RECT 669.400 61.920 669.660 62.180 ;
        RECT 674.000 61.920 674.260 62.180 ;
      LAYER met2 ;
        RECT 448.730 510.340 449.010 514.000 ;
        RECT 448.660 510.000 449.010 510.340 ;
        RECT 448.660 503.530 448.800 510.000 ;
        RECT 448.600 503.210 448.860 503.530 ;
        RECT 454.580 503.210 454.840 503.530 ;
        RECT 454.640 141.430 454.780 503.210 ;
        RECT 454.580 141.110 454.840 141.430 ;
        RECT 669.400 141.110 669.660 141.430 ;
        RECT 669.460 62.210 669.600 141.110 ;
        RECT 669.400 61.890 669.660 62.210 ;
        RECT 674.000 61.890 674.260 62.210 ;
        RECT 674.060 61.610 674.200 61.890 ;
        RECT 674.060 61.470 674.660 61.610 ;
        RECT 674.520 2.400 674.660 61.470 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 794.950 496.980 795.270 497.040 ;
        RECT 799.550 496.980 799.870 497.040 ;
        RECT 794.950 496.840 799.870 496.980 ;
        RECT 794.950 496.780 795.270 496.840 ;
        RECT 799.550 496.780 799.870 496.840 ;
        RECT 799.550 293.320 799.870 293.380 ;
        RECT 1173.070 293.320 1173.390 293.380 ;
        RECT 799.550 293.180 1173.390 293.320 ;
        RECT 799.550 293.120 799.870 293.180 ;
        RECT 1173.070 293.120 1173.390 293.180 ;
      LAYER via ;
        RECT 794.980 496.780 795.240 497.040 ;
        RECT 799.580 496.780 799.840 497.040 ;
        RECT 799.580 293.120 799.840 293.380 ;
        RECT 1173.100 293.120 1173.360 293.380 ;
      LAYER met2 ;
        RECT 795.110 510.340 795.390 514.000 ;
        RECT 795.040 510.000 795.390 510.340 ;
        RECT 795.040 497.070 795.180 510.000 ;
        RECT 794.980 496.750 795.240 497.070 ;
        RECT 799.580 496.750 799.840 497.070 ;
        RECT 799.640 293.410 799.780 496.750 ;
        RECT 799.580 293.090 799.840 293.410 ;
        RECT 1173.100 293.090 1173.360 293.410 ;
        RECT 1173.160 17.410 1173.300 293.090 ;
        RECT 1173.160 17.270 1174.220 17.410 ;
        RECT 1174.080 2.400 1174.220 17.270 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 807.370 496.980 807.690 497.040 ;
        RECT 813.350 496.980 813.670 497.040 ;
        RECT 807.370 496.840 813.670 496.980 ;
        RECT 807.370 496.780 807.690 496.840 ;
        RECT 813.350 496.780 813.670 496.840 ;
        RECT 813.350 300.120 813.670 300.180 ;
        RECT 1186.870 300.120 1187.190 300.180 ;
        RECT 813.350 299.980 1187.190 300.120 ;
        RECT 813.350 299.920 813.670 299.980 ;
        RECT 1186.870 299.920 1187.190 299.980 ;
      LAYER via ;
        RECT 807.400 496.780 807.660 497.040 ;
        RECT 813.380 496.780 813.640 497.040 ;
        RECT 813.380 299.920 813.640 300.180 ;
        RECT 1186.900 299.920 1187.160 300.180 ;
      LAYER met2 ;
        RECT 807.530 510.340 807.810 514.000 ;
        RECT 807.460 510.000 807.810 510.340 ;
        RECT 807.460 497.070 807.600 510.000 ;
        RECT 807.400 496.750 807.660 497.070 ;
        RECT 813.380 496.750 813.640 497.070 ;
        RECT 813.440 300.210 813.580 496.750 ;
        RECT 813.380 299.890 813.640 300.210 ;
        RECT 1186.900 299.890 1187.160 300.210 ;
        RECT 1186.960 17.410 1187.100 299.890 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 819.790 496.980 820.110 497.040 ;
        RECT 824.390 496.980 824.710 497.040 ;
        RECT 819.790 496.840 824.710 496.980 ;
        RECT 819.790 496.780 820.110 496.840 ;
        RECT 824.390 496.780 824.710 496.840 ;
        RECT 824.390 224.300 824.710 224.360 ;
        RECT 1207.570 224.300 1207.890 224.360 ;
        RECT 824.390 224.160 1207.890 224.300 ;
        RECT 824.390 224.100 824.710 224.160 ;
        RECT 1207.570 224.100 1207.890 224.160 ;
      LAYER via ;
        RECT 819.820 496.780 820.080 497.040 ;
        RECT 824.420 496.780 824.680 497.040 ;
        RECT 824.420 224.100 824.680 224.360 ;
        RECT 1207.600 224.100 1207.860 224.360 ;
      LAYER met2 ;
        RECT 819.950 510.340 820.230 514.000 ;
        RECT 819.880 510.000 820.230 510.340 ;
        RECT 819.880 497.070 820.020 510.000 ;
        RECT 819.820 496.750 820.080 497.070 ;
        RECT 824.420 496.750 824.680 497.070 ;
        RECT 824.480 224.390 824.620 496.750 ;
        RECT 824.420 224.070 824.680 224.390 ;
        RECT 1207.600 224.070 1207.860 224.390 ;
        RECT 1207.660 17.410 1207.800 224.070 ;
        RECT 1207.660 17.270 1210.100 17.410 ;
        RECT 1209.960 2.400 1210.100 17.270 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 834.510 307.260 834.830 307.320 ;
        RECT 1221.370 307.260 1221.690 307.320 ;
        RECT 834.510 307.120 1221.690 307.260 ;
        RECT 834.510 307.060 834.830 307.120 ;
        RECT 1221.370 307.060 1221.690 307.120 ;
        RECT 1221.370 17.580 1221.690 17.640 ;
        RECT 1227.810 17.580 1228.130 17.640 ;
        RECT 1221.370 17.440 1228.130 17.580 ;
        RECT 1221.370 17.380 1221.690 17.440 ;
        RECT 1227.810 17.380 1228.130 17.440 ;
      LAYER via ;
        RECT 834.540 307.060 834.800 307.320 ;
        RECT 1221.400 307.060 1221.660 307.320 ;
        RECT 1221.400 17.380 1221.660 17.640 ;
        RECT 1227.840 17.380 1228.100 17.640 ;
      LAYER met2 ;
        RECT 832.370 510.410 832.650 514.000 ;
        RECT 832.370 510.270 834.740 510.410 ;
        RECT 832.370 510.000 832.650 510.270 ;
        RECT 834.600 307.350 834.740 510.270 ;
        RECT 834.540 307.030 834.800 307.350 ;
        RECT 1221.400 307.030 1221.660 307.350 ;
        RECT 1221.460 17.670 1221.600 307.030 ;
        RECT 1221.400 17.350 1221.660 17.670 ;
        RECT 1227.840 17.350 1228.100 17.670 ;
        RECT 1227.900 2.400 1228.040 17.350 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 844.630 496.980 844.950 497.040 ;
        RECT 848.310 496.980 848.630 497.040 ;
        RECT 844.630 496.840 848.630 496.980 ;
        RECT 844.630 496.780 844.950 496.840 ;
        RECT 848.310 496.780 848.630 496.840 ;
        RECT 848.310 314.060 848.630 314.120 ;
        RECT 1242.070 314.060 1242.390 314.120 ;
        RECT 848.310 313.920 1242.390 314.060 ;
        RECT 848.310 313.860 848.630 313.920 ;
        RECT 1242.070 313.860 1242.390 313.920 ;
      LAYER via ;
        RECT 844.660 496.780 844.920 497.040 ;
        RECT 848.340 496.780 848.600 497.040 ;
        RECT 848.340 313.860 848.600 314.120 ;
        RECT 1242.100 313.860 1242.360 314.120 ;
      LAYER met2 ;
        RECT 844.790 510.340 845.070 514.000 ;
        RECT 844.720 510.000 845.070 510.340 ;
        RECT 844.720 497.070 844.860 510.000 ;
        RECT 844.660 496.750 844.920 497.070 ;
        RECT 848.340 496.750 848.600 497.070 ;
        RECT 848.400 314.150 848.540 496.750 ;
        RECT 848.340 313.830 848.600 314.150 ;
        RECT 1242.100 313.830 1242.360 314.150 ;
        RECT 1242.160 17.410 1242.300 313.830 ;
        RECT 1242.160 17.270 1245.980 17.410 ;
        RECT 1245.840 2.400 1245.980 17.270 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 857.050 496.980 857.370 497.040 ;
        RECT 862.110 496.980 862.430 497.040 ;
        RECT 857.050 496.840 862.430 496.980 ;
        RECT 857.050 496.780 857.370 496.840 ;
        RECT 862.110 496.780 862.430 496.840 ;
        RECT 862.110 320.860 862.430 320.920 ;
        RECT 1262.770 320.860 1263.090 320.920 ;
        RECT 862.110 320.720 1263.090 320.860 ;
        RECT 862.110 320.660 862.430 320.720 ;
        RECT 1262.770 320.660 1263.090 320.720 ;
      LAYER via ;
        RECT 857.080 496.780 857.340 497.040 ;
        RECT 862.140 496.780 862.400 497.040 ;
        RECT 862.140 320.660 862.400 320.920 ;
        RECT 1262.800 320.660 1263.060 320.920 ;
      LAYER met2 ;
        RECT 857.210 510.340 857.490 514.000 ;
        RECT 857.140 510.000 857.490 510.340 ;
        RECT 857.140 497.070 857.280 510.000 ;
        RECT 857.080 496.750 857.340 497.070 ;
        RECT 862.140 496.750 862.400 497.070 ;
        RECT 862.200 320.950 862.340 496.750 ;
        RECT 862.140 320.630 862.400 320.950 ;
        RECT 1262.800 320.630 1263.060 320.950 ;
        RECT 1262.860 17.410 1263.000 320.630 ;
        RECT 1262.860 17.270 1263.460 17.410 ;
        RECT 1263.320 2.400 1263.460 17.270 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 868.550 328.000 868.870 328.060 ;
        RECT 1276.570 328.000 1276.890 328.060 ;
        RECT 868.550 327.860 1276.890 328.000 ;
        RECT 868.550 327.800 868.870 327.860 ;
        RECT 1276.570 327.800 1276.890 327.860 ;
      LAYER via ;
        RECT 868.580 327.800 868.840 328.060 ;
        RECT 1276.600 327.800 1276.860 328.060 ;
      LAYER met2 ;
        RECT 869.170 510.410 869.450 514.000 ;
        RECT 868.640 510.270 869.450 510.410 ;
        RECT 868.640 328.090 868.780 510.270 ;
        RECT 869.170 510.000 869.450 510.270 ;
        RECT 868.580 327.770 868.840 328.090 ;
        RECT 1276.600 327.770 1276.860 328.090 ;
        RECT 1276.660 17.410 1276.800 327.770 ;
        RECT 1276.660 17.270 1281.400 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 882.350 334.800 882.670 334.860 ;
        RECT 1297.270 334.800 1297.590 334.860 ;
        RECT 882.350 334.660 1297.590 334.800 ;
        RECT 882.350 334.600 882.670 334.660 ;
        RECT 1297.270 334.600 1297.590 334.660 ;
      LAYER via ;
        RECT 882.380 334.600 882.640 334.860 ;
        RECT 1297.300 334.600 1297.560 334.860 ;
      LAYER met2 ;
        RECT 881.590 510.410 881.870 514.000 ;
        RECT 881.590 510.270 882.580 510.410 ;
        RECT 881.590 510.000 881.870 510.270 ;
        RECT 882.440 334.890 882.580 510.270 ;
        RECT 882.380 334.570 882.640 334.890 ;
        RECT 1297.300 334.570 1297.560 334.890 ;
        RECT 1297.360 17.410 1297.500 334.570 ;
        RECT 1297.360 17.270 1299.340 17.410 ;
        RECT 1299.200 2.400 1299.340 17.270 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 896.610 341.940 896.930 342.000 ;
        RECT 1311.070 341.940 1311.390 342.000 ;
        RECT 896.610 341.800 1311.390 341.940 ;
        RECT 896.610 341.740 896.930 341.800 ;
        RECT 1311.070 341.740 1311.390 341.800 ;
        RECT 1311.070 17.920 1311.390 17.980 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1311.070 17.780 1317.370 17.920 ;
        RECT 1311.070 17.720 1311.390 17.780 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
      LAYER via ;
        RECT 896.640 341.740 896.900 342.000 ;
        RECT 1311.100 341.740 1311.360 342.000 ;
        RECT 1311.100 17.720 1311.360 17.980 ;
        RECT 1317.080 17.720 1317.340 17.980 ;
      LAYER met2 ;
        RECT 894.010 510.410 894.290 514.000 ;
        RECT 894.010 510.270 896.840 510.410 ;
        RECT 894.010 510.000 894.290 510.270 ;
        RECT 896.700 342.030 896.840 510.270 ;
        RECT 896.640 341.710 896.900 342.030 ;
        RECT 1311.100 341.710 1311.360 342.030 ;
        RECT 1311.160 18.010 1311.300 341.710 ;
        RECT 1311.100 17.690 1311.360 18.010 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1317.140 2.400 1317.280 17.690 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.270 496.980 906.590 497.040 ;
        RECT 914.090 496.980 914.410 497.040 ;
        RECT 906.270 496.840 914.410 496.980 ;
        RECT 906.270 496.780 906.590 496.840 ;
        RECT 914.090 496.780 914.410 496.840 ;
        RECT 914.090 349.080 914.410 349.140 ;
        RECT 1331.770 349.080 1332.090 349.140 ;
        RECT 914.090 348.940 1332.090 349.080 ;
        RECT 914.090 348.880 914.410 348.940 ;
        RECT 1331.770 348.880 1332.090 348.940 ;
        RECT 1331.770 62.120 1332.090 62.180 ;
        RECT 1334.990 62.120 1335.310 62.180 ;
        RECT 1331.770 61.980 1335.310 62.120 ;
        RECT 1331.770 61.920 1332.090 61.980 ;
        RECT 1334.990 61.920 1335.310 61.980 ;
      LAYER via ;
        RECT 906.300 496.780 906.560 497.040 ;
        RECT 914.120 496.780 914.380 497.040 ;
        RECT 914.120 348.880 914.380 349.140 ;
        RECT 1331.800 348.880 1332.060 349.140 ;
        RECT 1331.800 61.920 1332.060 62.180 ;
        RECT 1335.020 61.920 1335.280 62.180 ;
      LAYER met2 ;
        RECT 906.430 510.340 906.710 514.000 ;
        RECT 906.360 510.000 906.710 510.340 ;
        RECT 906.360 497.070 906.500 510.000 ;
        RECT 906.300 496.750 906.560 497.070 ;
        RECT 914.120 496.750 914.380 497.070 ;
        RECT 914.180 349.170 914.320 496.750 ;
        RECT 914.120 348.850 914.380 349.170 ;
        RECT 1331.800 348.850 1332.060 349.170 ;
        RECT 1331.860 62.210 1332.000 348.850 ;
        RECT 1331.800 61.890 1332.060 62.210 ;
        RECT 1335.020 61.890 1335.280 62.210 ;
        RECT 1335.080 2.400 1335.220 61.890 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 461.065 427.805 461.235 448.715 ;
        RECT 461.065 338.045 461.235 403.835 ;
        RECT 460.605 241.485 460.775 289.595 ;
        RECT 690.145 186.405 690.315 234.515 ;
      LAYER mcon ;
        RECT 461.065 448.545 461.235 448.715 ;
        RECT 461.065 403.665 461.235 403.835 ;
        RECT 460.605 289.425 460.775 289.595 ;
        RECT 690.145 234.345 690.315 234.515 ;
      LAYER met1 ;
        RECT 460.530 476.580 460.850 476.640 ;
        RECT 460.530 476.440 461.680 476.580 ;
        RECT 460.530 476.380 460.850 476.440 ;
        RECT 461.540 476.300 461.680 476.440 ;
        RECT 461.450 476.040 461.770 476.300 ;
        RECT 460.990 448.700 461.310 448.760 ;
        RECT 460.795 448.560 461.310 448.700 ;
        RECT 460.990 448.500 461.310 448.560 ;
        RECT 460.990 427.960 461.310 428.020 ;
        RECT 460.795 427.820 461.310 427.960 ;
        RECT 460.990 427.760 461.310 427.820 ;
        RECT 459.610 403.820 459.930 403.880 ;
        RECT 461.005 403.820 461.295 403.865 ;
        RECT 459.610 403.680 461.295 403.820 ;
        RECT 459.610 403.620 459.930 403.680 ;
        RECT 461.005 403.635 461.295 403.680 ;
        RECT 461.005 338.200 461.295 338.245 ;
        RECT 461.450 338.200 461.770 338.260 ;
        RECT 461.005 338.060 461.770 338.200 ;
        RECT 461.005 338.015 461.295 338.060 ;
        RECT 461.450 338.000 461.770 338.060 ;
        RECT 460.545 289.580 460.835 289.625 ;
        RECT 460.990 289.580 461.310 289.640 ;
        RECT 460.545 289.440 461.310 289.580 ;
        RECT 460.545 289.395 460.835 289.440 ;
        RECT 460.990 289.380 461.310 289.440 ;
        RECT 460.530 241.640 460.850 241.700 ;
        RECT 460.335 241.500 460.850 241.640 ;
        RECT 460.530 241.440 460.850 241.500 ;
        RECT 460.530 237.900 460.850 237.960 ;
        RECT 690.070 237.900 690.390 237.960 ;
        RECT 460.530 237.760 690.390 237.900 ;
        RECT 460.530 237.700 460.850 237.760 ;
        RECT 690.070 237.700 690.390 237.760 ;
        RECT 690.070 234.500 690.390 234.560 ;
        RECT 689.875 234.360 690.390 234.500 ;
        RECT 690.070 234.300 690.390 234.360 ;
        RECT 690.070 186.560 690.390 186.620 ;
        RECT 689.875 186.420 690.390 186.560 ;
        RECT 690.070 186.360 690.390 186.420 ;
        RECT 690.070 137.940 690.390 138.000 ;
        RECT 692.370 137.940 692.690 138.000 ;
        RECT 690.070 137.800 692.690 137.940 ;
        RECT 690.070 137.740 690.390 137.800 ;
        RECT 692.370 137.740 692.690 137.800 ;
      LAYER via ;
        RECT 460.560 476.380 460.820 476.640 ;
        RECT 461.480 476.040 461.740 476.300 ;
        RECT 461.020 448.500 461.280 448.760 ;
        RECT 461.020 427.760 461.280 428.020 ;
        RECT 459.640 403.620 459.900 403.880 ;
        RECT 461.480 338.000 461.740 338.260 ;
        RECT 461.020 289.380 461.280 289.640 ;
        RECT 460.560 241.440 460.820 241.700 ;
        RECT 460.560 237.700 460.820 237.960 ;
        RECT 690.100 237.700 690.360 237.960 ;
        RECT 690.100 234.300 690.360 234.560 ;
        RECT 690.100 186.360 690.360 186.620 ;
        RECT 690.100 137.740 690.360 138.000 ;
        RECT 692.400 137.740 692.660 138.000 ;
      LAYER met2 ;
        RECT 461.150 510.410 461.430 514.000 ;
        RECT 460.620 510.270 461.430 510.410 ;
        RECT 460.620 476.670 460.760 510.270 ;
        RECT 461.150 510.000 461.430 510.270 ;
        RECT 460.560 476.350 460.820 476.670 ;
        RECT 461.480 476.010 461.740 476.330 ;
        RECT 461.540 475.730 461.680 476.010 ;
        RECT 461.080 475.590 461.680 475.730 ;
        RECT 461.080 448.790 461.220 475.590 ;
        RECT 461.020 448.470 461.280 448.790 ;
        RECT 461.020 427.730 461.280 428.050 ;
        RECT 461.080 427.565 461.220 427.730 ;
        RECT 459.630 427.195 459.910 427.565 ;
        RECT 461.010 427.195 461.290 427.565 ;
        RECT 459.700 403.910 459.840 427.195 ;
        RECT 459.640 403.590 459.900 403.910 ;
        RECT 461.480 337.970 461.740 338.290 ;
        RECT 461.540 303.010 461.680 337.970 ;
        RECT 461.080 302.870 461.680 303.010 ;
        RECT 461.080 289.670 461.220 302.870 ;
        RECT 461.020 289.350 461.280 289.670 ;
        RECT 460.560 241.410 460.820 241.730 ;
        RECT 460.620 237.990 460.760 241.410 ;
        RECT 460.560 237.670 460.820 237.990 ;
        RECT 690.100 237.670 690.360 237.990 ;
        RECT 690.160 234.590 690.300 237.670 ;
        RECT 690.100 234.270 690.360 234.590 ;
        RECT 690.100 186.330 690.360 186.650 ;
        RECT 690.160 138.030 690.300 186.330 ;
        RECT 690.100 137.710 690.360 138.030 ;
        RECT 692.400 137.710 692.660 138.030 ;
        RECT 692.460 2.400 692.600 137.710 ;
        RECT 692.250 -4.800 692.810 2.400 ;
      LAYER via2 ;
        RECT 459.630 427.240 459.910 427.520 ;
        RECT 461.010 427.240 461.290 427.520 ;
      LAYER met3 ;
        RECT 459.605 427.530 459.935 427.545 ;
        RECT 460.985 427.530 461.315 427.545 ;
        RECT 459.605 427.230 461.315 427.530 ;
        RECT 459.605 427.215 459.935 427.230 ;
        RECT 460.985 427.215 461.315 427.230 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 918.690 497.320 919.010 497.380 ;
        RECT 934.790 497.320 935.110 497.380 ;
        RECT 918.690 497.180 935.110 497.320 ;
        RECT 918.690 497.120 919.010 497.180 ;
        RECT 934.790 497.120 935.110 497.180 ;
        RECT 934.790 355.540 935.110 355.600 ;
        RECT 1352.470 355.540 1352.790 355.600 ;
        RECT 934.790 355.400 1352.790 355.540 ;
        RECT 934.790 355.340 935.110 355.400 ;
        RECT 1352.470 355.340 1352.790 355.400 ;
      LAYER via ;
        RECT 918.720 497.120 918.980 497.380 ;
        RECT 934.820 497.120 935.080 497.380 ;
        RECT 934.820 355.340 935.080 355.600 ;
        RECT 1352.500 355.340 1352.760 355.600 ;
      LAYER met2 ;
        RECT 918.850 510.340 919.130 514.000 ;
        RECT 918.780 510.000 919.130 510.340 ;
        RECT 918.780 497.410 918.920 510.000 ;
        RECT 918.720 497.090 918.980 497.410 ;
        RECT 934.820 497.090 935.080 497.410 ;
        RECT 934.880 355.630 935.020 497.090 ;
        RECT 934.820 355.310 935.080 355.630 ;
        RECT 1352.500 355.310 1352.760 355.630 ;
        RECT 1352.560 2.400 1352.700 355.310 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 930.650 362.680 930.970 362.740 ;
        RECT 1366.270 362.680 1366.590 362.740 ;
        RECT 930.650 362.540 1366.590 362.680 ;
        RECT 930.650 362.480 930.970 362.540 ;
        RECT 1366.270 362.480 1366.590 362.540 ;
      LAYER via ;
        RECT 930.680 362.480 930.940 362.740 ;
        RECT 1366.300 362.480 1366.560 362.740 ;
      LAYER met2 ;
        RECT 931.270 510.410 931.550 514.000 ;
        RECT 930.740 510.270 931.550 510.410 ;
        RECT 930.740 362.770 930.880 510.270 ;
        RECT 931.270 510.000 931.550 510.270 ;
        RECT 930.680 362.450 930.940 362.770 ;
        RECT 1366.300 362.450 1366.560 362.770 ;
        RECT 1366.360 17.410 1366.500 362.450 ;
        RECT 1366.360 17.270 1370.640 17.410 ;
        RECT 1370.500 2.400 1370.640 17.270 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.450 369.480 944.770 369.540 ;
        RECT 1386.970 369.480 1387.290 369.540 ;
        RECT 944.450 369.340 1387.290 369.480 ;
        RECT 944.450 369.280 944.770 369.340 ;
        RECT 1386.970 369.280 1387.290 369.340 ;
      LAYER via ;
        RECT 944.480 369.280 944.740 369.540 ;
        RECT 1387.000 369.280 1387.260 369.540 ;
      LAYER met2 ;
        RECT 943.690 510.410 943.970 514.000 ;
        RECT 943.690 510.270 944.680 510.410 ;
        RECT 943.690 510.000 943.970 510.270 ;
        RECT 944.540 369.570 944.680 510.270 ;
        RECT 944.480 369.250 944.740 369.570 ;
        RECT 1387.000 369.250 1387.260 369.570 ;
        RECT 1387.060 17.410 1387.200 369.250 ;
        RECT 1387.060 17.270 1388.580 17.410 ;
        RECT 1388.440 2.400 1388.580 17.270 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 958.710 376.280 959.030 376.340 ;
        RECT 1400.770 376.280 1401.090 376.340 ;
        RECT 958.710 376.140 1401.090 376.280 ;
        RECT 958.710 376.080 959.030 376.140 ;
        RECT 1400.770 376.080 1401.090 376.140 ;
      LAYER via ;
        RECT 958.740 376.080 959.000 376.340 ;
        RECT 1400.800 376.080 1401.060 376.340 ;
      LAYER met2 ;
        RECT 956.110 510.410 956.390 514.000 ;
        RECT 956.110 510.270 958.940 510.410 ;
        RECT 956.110 510.000 956.390 510.270 ;
        RECT 958.800 376.370 958.940 510.270 ;
        RECT 958.740 376.050 959.000 376.370 ;
        RECT 1400.800 376.050 1401.060 376.370 ;
        RECT 1400.860 17.410 1401.000 376.050 ;
        RECT 1400.860 17.270 1406.520 17.410 ;
        RECT 1406.380 2.400 1406.520 17.270 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 972.050 382.740 972.370 382.800 ;
        RECT 1421.470 382.740 1421.790 382.800 ;
        RECT 972.050 382.600 1421.790 382.740 ;
        RECT 972.050 382.540 972.370 382.600 ;
        RECT 1421.470 382.540 1421.790 382.600 ;
      LAYER via ;
        RECT 972.080 382.540 972.340 382.800 ;
        RECT 1421.500 382.540 1421.760 382.800 ;
      LAYER met2 ;
        RECT 968.530 510.410 968.810 514.000 ;
        RECT 968.530 510.270 972.280 510.410 ;
        RECT 968.530 510.000 968.810 510.270 ;
        RECT 972.140 382.830 972.280 510.270 ;
        RECT 972.080 382.510 972.340 382.830 ;
        RECT 1421.500 382.510 1421.760 382.830 ;
        RECT 1421.560 17.410 1421.700 382.510 ;
        RECT 1421.560 17.270 1424.000 17.410 ;
        RECT 1423.860 2.400 1424.000 17.270 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 980.330 472.500 980.650 472.560 ;
        RECT 1435.270 472.500 1435.590 472.560 ;
        RECT 980.330 472.360 1435.590 472.500 ;
        RECT 980.330 472.300 980.650 472.360 ;
        RECT 1435.270 472.300 1435.590 472.360 ;
        RECT 1435.270 7.040 1435.590 7.100 ;
        RECT 1441.710 7.040 1442.030 7.100 ;
        RECT 1435.270 6.900 1442.030 7.040 ;
        RECT 1435.270 6.840 1435.590 6.900 ;
        RECT 1441.710 6.840 1442.030 6.900 ;
      LAYER via ;
        RECT 980.360 472.300 980.620 472.560 ;
        RECT 1435.300 472.300 1435.560 472.560 ;
        RECT 1435.300 6.840 1435.560 7.100 ;
        RECT 1441.740 6.840 1442.000 7.100 ;
      LAYER met2 ;
        RECT 980.490 510.340 980.770 514.000 ;
        RECT 980.420 510.000 980.770 510.340 ;
        RECT 980.420 472.590 980.560 510.000 ;
        RECT 980.360 472.270 980.620 472.590 ;
        RECT 1435.300 472.270 1435.560 472.590 ;
        RECT 1435.360 7.130 1435.500 472.270 ;
        RECT 1435.300 6.810 1435.560 7.130 ;
        RECT 1441.740 6.810 1442.000 7.130 ;
        RECT 1441.800 2.400 1441.940 6.810 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 992.825 427.805 992.995 448.715 ;
      LAYER mcon ;
        RECT 992.825 448.545 992.995 448.715 ;
      LAYER met1 ;
        RECT 992.750 448.700 993.070 448.760 ;
        RECT 992.555 448.560 993.070 448.700 ;
        RECT 992.750 448.500 993.070 448.560 ;
        RECT 992.750 427.960 993.070 428.020 ;
        RECT 992.555 427.820 993.070 427.960 ;
        RECT 992.750 427.760 993.070 427.820 ;
        RECT 992.750 390.220 993.070 390.280 ;
        RECT 1455.970 390.220 1456.290 390.280 ;
        RECT 992.750 390.080 1456.290 390.220 ;
        RECT 992.750 390.020 993.070 390.080 ;
        RECT 1455.970 390.020 1456.290 390.080 ;
      LAYER via ;
        RECT 992.780 448.500 993.040 448.760 ;
        RECT 992.780 427.760 993.040 428.020 ;
        RECT 992.780 390.020 993.040 390.280 ;
        RECT 1456.000 390.020 1456.260 390.280 ;
      LAYER met2 ;
        RECT 992.910 510.340 993.190 514.000 ;
        RECT 992.840 510.000 993.190 510.340 ;
        RECT 992.840 448.790 992.980 510.000 ;
        RECT 992.780 448.470 993.040 448.790 ;
        RECT 992.780 427.730 993.040 428.050 ;
        RECT 992.840 390.310 992.980 427.730 ;
        RECT 992.780 389.990 993.040 390.310 ;
        RECT 1456.000 389.990 1456.260 390.310 ;
        RECT 1456.060 18.090 1456.200 389.990 ;
        RECT 1456.060 17.950 1459.880 18.090 ;
        RECT 1459.740 2.400 1459.880 17.950 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1006.550 397.020 1006.870 397.080 ;
        RECT 1476.670 397.020 1476.990 397.080 ;
        RECT 1006.550 396.880 1476.990 397.020 ;
        RECT 1006.550 396.820 1006.870 396.880 ;
        RECT 1476.670 396.820 1476.990 396.880 ;
      LAYER via ;
        RECT 1006.580 396.820 1006.840 397.080 ;
        RECT 1476.700 396.820 1476.960 397.080 ;
      LAYER met2 ;
        RECT 1005.330 510.410 1005.610 514.000 ;
        RECT 1005.330 510.270 1006.780 510.410 ;
        RECT 1005.330 510.000 1005.610 510.270 ;
        RECT 1006.640 397.110 1006.780 510.270 ;
        RECT 1006.580 396.790 1006.840 397.110 ;
        RECT 1476.700 396.790 1476.960 397.110 ;
        RECT 1476.760 17.410 1476.900 396.790 ;
        RECT 1476.760 17.270 1477.820 17.410 ;
        RECT 1477.680 2.400 1477.820 17.270 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1020.810 403.480 1021.130 403.540 ;
        RECT 1490.470 403.480 1490.790 403.540 ;
        RECT 1020.810 403.340 1490.790 403.480 ;
        RECT 1020.810 403.280 1021.130 403.340 ;
        RECT 1490.470 403.280 1490.790 403.340 ;
      LAYER via ;
        RECT 1020.840 403.280 1021.100 403.540 ;
        RECT 1490.500 403.280 1490.760 403.540 ;
      LAYER met2 ;
        RECT 1017.750 510.410 1018.030 514.000 ;
        RECT 1017.750 510.270 1021.040 510.410 ;
        RECT 1017.750 510.000 1018.030 510.270 ;
        RECT 1020.900 403.570 1021.040 510.270 ;
        RECT 1020.840 403.250 1021.100 403.570 ;
        RECT 1490.500 403.250 1490.760 403.570 ;
        RECT 1490.560 16.730 1490.700 403.250 ;
        RECT 1490.560 16.590 1495.760 16.730 ;
        RECT 1495.620 2.400 1495.760 16.590 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1030.010 496.980 1030.330 497.040 ;
        RECT 1034.150 496.980 1034.470 497.040 ;
        RECT 1030.010 496.840 1034.470 496.980 ;
        RECT 1030.010 496.780 1030.330 496.840 ;
        RECT 1034.150 496.780 1034.470 496.840 ;
        RECT 1034.150 417.420 1034.470 417.480 ;
        RECT 1511.170 417.420 1511.490 417.480 ;
        RECT 1034.150 417.280 1511.490 417.420 ;
        RECT 1034.150 417.220 1034.470 417.280 ;
        RECT 1511.170 417.220 1511.490 417.280 ;
      LAYER via ;
        RECT 1030.040 496.780 1030.300 497.040 ;
        RECT 1034.180 496.780 1034.440 497.040 ;
        RECT 1034.180 417.220 1034.440 417.480 ;
        RECT 1511.200 417.220 1511.460 417.480 ;
      LAYER met2 ;
        RECT 1030.170 510.340 1030.450 514.000 ;
        RECT 1030.100 510.000 1030.450 510.340 ;
        RECT 1030.100 497.070 1030.240 510.000 ;
        RECT 1030.040 496.750 1030.300 497.070 ;
        RECT 1034.180 496.750 1034.440 497.070 ;
        RECT 1034.240 417.510 1034.380 496.750 ;
        RECT 1034.180 417.190 1034.440 417.510 ;
        RECT 1511.200 417.190 1511.460 417.510 ;
        RECT 1511.260 16.730 1511.400 417.190 ;
        RECT 1511.260 16.590 1513.240 16.730 ;
        RECT 1513.100 2.400 1513.240 16.590 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 475.710 245.040 476.030 245.100 ;
        RECT 703.870 245.040 704.190 245.100 ;
        RECT 475.710 244.900 704.190 245.040 ;
        RECT 475.710 244.840 476.030 244.900 ;
        RECT 703.870 244.840 704.190 244.900 ;
        RECT 703.870 38.320 704.190 38.380 ;
        RECT 710.310 38.320 710.630 38.380 ;
        RECT 703.870 38.180 710.630 38.320 ;
        RECT 703.870 38.120 704.190 38.180 ;
        RECT 710.310 38.120 710.630 38.180 ;
      LAYER via ;
        RECT 475.740 244.840 476.000 245.100 ;
        RECT 703.900 244.840 704.160 245.100 ;
        RECT 703.900 38.120 704.160 38.380 ;
        RECT 710.340 38.120 710.600 38.380 ;
      LAYER met2 ;
        RECT 473.570 510.410 473.850 514.000 ;
        RECT 473.570 510.270 475.940 510.410 ;
        RECT 473.570 510.000 473.850 510.270 ;
        RECT 475.800 245.130 475.940 510.270 ;
        RECT 475.740 244.810 476.000 245.130 ;
        RECT 703.900 244.810 704.160 245.130 ;
        RECT 703.960 38.410 704.100 244.810 ;
        RECT 703.900 38.090 704.160 38.410 ;
        RECT 710.340 38.090 710.600 38.410 ;
        RECT 710.400 2.400 710.540 38.090 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1042.430 496.980 1042.750 497.040 ;
        RECT 1047.950 496.980 1048.270 497.040 ;
        RECT 1042.430 496.840 1048.270 496.980 ;
        RECT 1042.430 496.780 1042.750 496.840 ;
        RECT 1047.950 496.780 1048.270 496.840 ;
        RECT 1047.950 424.220 1048.270 424.280 ;
        RECT 1524.970 424.220 1525.290 424.280 ;
        RECT 1047.950 424.080 1525.290 424.220 ;
        RECT 1047.950 424.020 1048.270 424.080 ;
        RECT 1524.970 424.020 1525.290 424.080 ;
        RECT 1524.970 17.920 1525.290 17.980 ;
        RECT 1530.950 17.920 1531.270 17.980 ;
        RECT 1524.970 17.780 1531.270 17.920 ;
        RECT 1524.970 17.720 1525.290 17.780 ;
        RECT 1530.950 17.720 1531.270 17.780 ;
      LAYER via ;
        RECT 1042.460 496.780 1042.720 497.040 ;
        RECT 1047.980 496.780 1048.240 497.040 ;
        RECT 1047.980 424.020 1048.240 424.280 ;
        RECT 1525.000 424.020 1525.260 424.280 ;
        RECT 1525.000 17.720 1525.260 17.980 ;
        RECT 1530.980 17.720 1531.240 17.980 ;
      LAYER met2 ;
        RECT 1042.590 510.340 1042.870 514.000 ;
        RECT 1042.520 510.000 1042.870 510.340 ;
        RECT 1042.520 497.070 1042.660 510.000 ;
        RECT 1042.460 496.750 1042.720 497.070 ;
        RECT 1047.980 496.750 1048.240 497.070 ;
        RECT 1048.040 424.310 1048.180 496.750 ;
        RECT 1047.980 423.990 1048.240 424.310 ;
        RECT 1525.000 423.990 1525.260 424.310 ;
        RECT 1525.060 18.010 1525.200 423.990 ;
        RECT 1525.000 17.690 1525.260 18.010 ;
        RECT 1530.980 17.690 1531.240 18.010 ;
        RECT 1531.040 2.400 1531.180 17.690 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1055.310 431.360 1055.630 431.420 ;
        RECT 1545.670 431.360 1545.990 431.420 ;
        RECT 1055.310 431.220 1545.990 431.360 ;
        RECT 1055.310 431.160 1055.630 431.220 ;
        RECT 1545.670 431.160 1545.990 431.220 ;
        RECT 1545.670 2.960 1545.990 3.020 ;
        RECT 1548.890 2.960 1549.210 3.020 ;
        RECT 1545.670 2.820 1549.210 2.960 ;
        RECT 1545.670 2.760 1545.990 2.820 ;
        RECT 1548.890 2.760 1549.210 2.820 ;
      LAYER via ;
        RECT 1055.340 431.160 1055.600 431.420 ;
        RECT 1545.700 431.160 1545.960 431.420 ;
        RECT 1545.700 2.760 1545.960 3.020 ;
        RECT 1548.920 2.760 1549.180 3.020 ;
      LAYER met2 ;
        RECT 1055.010 510.340 1055.290 514.000 ;
        RECT 1054.940 510.000 1055.290 510.340 ;
        RECT 1054.940 497.490 1055.080 510.000 ;
        RECT 1054.940 497.350 1055.540 497.490 ;
        RECT 1055.400 431.450 1055.540 497.350 ;
        RECT 1055.340 431.130 1055.600 431.450 ;
        RECT 1545.700 431.130 1545.960 431.450 ;
        RECT 1545.760 3.050 1545.900 431.130 ;
        RECT 1545.700 2.730 1545.960 3.050 ;
        RECT 1548.920 2.730 1549.180 3.050 ;
        RECT 1548.980 2.400 1549.120 2.730 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1068.650 451.760 1068.970 451.820 ;
        RECT 1566.370 451.760 1566.690 451.820 ;
        RECT 1068.650 451.620 1566.690 451.760 ;
        RECT 1068.650 451.560 1068.970 451.620 ;
        RECT 1566.370 451.560 1566.690 451.620 ;
      LAYER via ;
        RECT 1068.680 451.560 1068.940 451.820 ;
        RECT 1566.400 451.560 1566.660 451.820 ;
      LAYER met2 ;
        RECT 1067.430 510.410 1067.710 514.000 ;
        RECT 1067.430 510.270 1068.880 510.410 ;
        RECT 1067.430 510.000 1067.710 510.270 ;
        RECT 1068.740 451.850 1068.880 510.270 ;
        RECT 1068.680 451.530 1068.940 451.850 ;
        RECT 1566.400 451.530 1566.660 451.850 ;
        RECT 1566.460 17.410 1566.600 451.530 ;
        RECT 1566.460 17.270 1567.060 17.410 ;
        RECT 1566.920 2.400 1567.060 17.270 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1082.910 458.900 1083.230 458.960 ;
        RECT 1580.170 458.900 1580.490 458.960 ;
        RECT 1082.910 458.760 1580.490 458.900 ;
        RECT 1082.910 458.700 1083.230 458.760 ;
        RECT 1580.170 458.700 1580.490 458.760 ;
      LAYER via ;
        RECT 1082.940 458.700 1083.200 458.960 ;
        RECT 1580.200 458.700 1580.460 458.960 ;
      LAYER met2 ;
        RECT 1079.850 510.410 1080.130 514.000 ;
        RECT 1079.850 510.270 1083.140 510.410 ;
        RECT 1079.850 510.000 1080.130 510.270 ;
        RECT 1083.000 458.990 1083.140 510.270 ;
        RECT 1082.940 458.670 1083.200 458.990 ;
        RECT 1580.200 458.670 1580.460 458.990 ;
        RECT 1580.260 16.730 1580.400 458.670 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1092.110 496.980 1092.430 497.040 ;
        RECT 1096.250 496.980 1096.570 497.040 ;
        RECT 1092.110 496.840 1096.570 496.980 ;
        RECT 1092.110 496.780 1092.430 496.840 ;
        RECT 1096.250 496.780 1096.570 496.840 ;
        RECT 1096.250 465.700 1096.570 465.760 ;
        RECT 1600.870 465.700 1601.190 465.760 ;
        RECT 1096.250 465.560 1601.190 465.700 ;
        RECT 1096.250 465.500 1096.570 465.560 ;
        RECT 1600.870 465.500 1601.190 465.560 ;
      LAYER via ;
        RECT 1092.140 496.780 1092.400 497.040 ;
        RECT 1096.280 496.780 1096.540 497.040 ;
        RECT 1096.280 465.500 1096.540 465.760 ;
        RECT 1600.900 465.500 1601.160 465.760 ;
      LAYER met2 ;
        RECT 1092.270 510.340 1092.550 514.000 ;
        RECT 1092.200 510.000 1092.550 510.340 ;
        RECT 1092.200 497.070 1092.340 510.000 ;
        RECT 1092.140 496.750 1092.400 497.070 ;
        RECT 1096.280 496.750 1096.540 497.070 ;
        RECT 1096.340 465.790 1096.480 496.750 ;
        RECT 1096.280 465.470 1096.540 465.790 ;
        RECT 1600.900 465.470 1601.160 465.790 ;
        RECT 1600.960 16.730 1601.100 465.470 ;
        RECT 1600.960 16.590 1602.480 16.730 ;
        RECT 1602.340 2.400 1602.480 16.590 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1104.070 496.980 1104.390 497.040 ;
        RECT 1110.510 496.980 1110.830 497.040 ;
        RECT 1104.070 496.840 1110.830 496.980 ;
        RECT 1104.070 496.780 1104.390 496.840 ;
        RECT 1110.510 496.780 1110.830 496.840 ;
        RECT 1110.510 38.320 1110.830 38.380 ;
        RECT 1620.190 38.320 1620.510 38.380 ;
        RECT 1110.510 38.180 1620.510 38.320 ;
        RECT 1110.510 38.120 1110.830 38.180 ;
        RECT 1620.190 38.120 1620.510 38.180 ;
      LAYER via ;
        RECT 1104.100 496.780 1104.360 497.040 ;
        RECT 1110.540 496.780 1110.800 497.040 ;
        RECT 1110.540 38.120 1110.800 38.380 ;
        RECT 1620.220 38.120 1620.480 38.380 ;
      LAYER met2 ;
        RECT 1104.230 510.340 1104.510 514.000 ;
        RECT 1104.160 510.000 1104.510 510.340 ;
        RECT 1104.160 497.070 1104.300 510.000 ;
        RECT 1104.100 496.750 1104.360 497.070 ;
        RECT 1110.540 496.750 1110.800 497.070 ;
        RECT 1110.600 38.410 1110.740 496.750 ;
        RECT 1110.540 38.090 1110.800 38.410 ;
        RECT 1620.220 38.090 1620.480 38.410 ;
        RECT 1620.280 2.400 1620.420 38.090 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1117.410 45.120 1117.730 45.180 ;
        RECT 1638.130 45.120 1638.450 45.180 ;
        RECT 1117.410 44.980 1638.450 45.120 ;
        RECT 1117.410 44.920 1117.730 44.980 ;
        RECT 1638.130 44.920 1638.450 44.980 ;
      LAYER via ;
        RECT 1117.440 44.920 1117.700 45.180 ;
        RECT 1638.160 44.920 1638.420 45.180 ;
      LAYER met2 ;
        RECT 1116.650 510.410 1116.930 514.000 ;
        RECT 1116.650 510.270 1117.640 510.410 ;
        RECT 1116.650 510.000 1116.930 510.270 ;
        RECT 1117.500 45.210 1117.640 510.270 ;
        RECT 1117.440 44.890 1117.700 45.210 ;
        RECT 1638.160 44.890 1638.420 45.210 ;
        RECT 1638.220 2.400 1638.360 44.890 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1128.910 479.640 1129.230 479.700 ;
        RECT 1656.070 479.640 1656.390 479.700 ;
        RECT 1128.910 479.500 1656.390 479.640 ;
        RECT 1128.910 479.440 1129.230 479.500 ;
        RECT 1656.070 479.440 1656.390 479.500 ;
      LAYER via ;
        RECT 1128.940 479.440 1129.200 479.700 ;
        RECT 1656.100 479.440 1656.360 479.700 ;
      LAYER met2 ;
        RECT 1129.070 510.340 1129.350 514.000 ;
        RECT 1129.000 510.000 1129.350 510.340 ;
        RECT 1129.000 479.730 1129.140 510.000 ;
        RECT 1128.940 479.410 1129.200 479.730 ;
        RECT 1656.100 479.410 1656.360 479.730 ;
        RECT 1656.160 2.400 1656.300 479.410 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1141.330 493.920 1141.650 493.980 ;
        RECT 1669.870 493.920 1670.190 493.980 ;
        RECT 1141.330 493.780 1670.190 493.920 ;
        RECT 1141.330 493.720 1141.650 493.780 ;
        RECT 1669.870 493.720 1670.190 493.780 ;
      LAYER via ;
        RECT 1141.360 493.720 1141.620 493.980 ;
        RECT 1669.900 493.720 1670.160 493.980 ;
      LAYER met2 ;
        RECT 1141.490 510.340 1141.770 514.000 ;
        RECT 1141.420 510.000 1141.770 510.340 ;
        RECT 1141.420 494.010 1141.560 510.000 ;
        RECT 1141.360 493.690 1141.620 494.010 ;
        RECT 1669.900 493.690 1670.160 494.010 ;
        RECT 1669.960 17.410 1670.100 493.690 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.750 486.440 1154.070 486.500 ;
        RECT 1690.570 486.440 1690.890 486.500 ;
        RECT 1153.750 486.300 1690.890 486.440 ;
        RECT 1153.750 486.240 1154.070 486.300 ;
        RECT 1690.570 486.240 1690.890 486.300 ;
      LAYER via ;
        RECT 1153.780 486.240 1154.040 486.500 ;
        RECT 1690.600 486.240 1690.860 486.500 ;
      LAYER met2 ;
        RECT 1153.910 510.340 1154.190 514.000 ;
        RECT 1153.840 510.000 1154.190 510.340 ;
        RECT 1153.840 486.530 1153.980 510.000 ;
        RECT 1153.780 486.210 1154.040 486.530 ;
        RECT 1690.600 486.210 1690.860 486.530 ;
        RECT 1690.660 17.410 1690.800 486.210 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 485.830 503.440 486.150 503.500 ;
        RECT 489.510 503.440 489.830 503.500 ;
        RECT 485.830 503.300 489.830 503.440 ;
        RECT 485.830 503.240 486.150 503.300 ;
        RECT 489.510 503.240 489.830 503.300 ;
        RECT 489.510 258.640 489.830 258.700 ;
        RECT 724.570 258.640 724.890 258.700 ;
        RECT 489.510 258.500 724.890 258.640 ;
        RECT 489.510 258.440 489.830 258.500 ;
        RECT 724.570 258.440 724.890 258.500 ;
        RECT 724.570 62.120 724.890 62.180 ;
        RECT 728.250 62.120 728.570 62.180 ;
        RECT 724.570 61.980 728.570 62.120 ;
        RECT 724.570 61.920 724.890 61.980 ;
        RECT 728.250 61.920 728.570 61.980 ;
      LAYER via ;
        RECT 485.860 503.240 486.120 503.500 ;
        RECT 489.540 503.240 489.800 503.500 ;
        RECT 489.540 258.440 489.800 258.700 ;
        RECT 724.600 258.440 724.860 258.700 ;
        RECT 724.600 61.920 724.860 62.180 ;
        RECT 728.280 61.920 728.540 62.180 ;
      LAYER met2 ;
        RECT 485.990 510.340 486.270 514.000 ;
        RECT 485.920 510.000 486.270 510.340 ;
        RECT 485.920 503.530 486.060 510.000 ;
        RECT 485.860 503.210 486.120 503.530 ;
        RECT 489.540 503.210 489.800 503.530 ;
        RECT 489.600 258.730 489.740 503.210 ;
        RECT 489.540 258.410 489.800 258.730 ;
        RECT 724.600 258.410 724.860 258.730 ;
        RECT 724.660 62.210 724.800 258.410 ;
        RECT 724.600 61.890 724.860 62.210 ;
        RECT 728.280 61.890 728.540 62.210 ;
        RECT 728.340 2.400 728.480 61.890 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1166.170 496.980 1166.490 497.040 ;
        RECT 1172.150 496.980 1172.470 497.040 ;
        RECT 1166.170 496.840 1172.470 496.980 ;
        RECT 1166.170 496.780 1166.490 496.840 ;
        RECT 1172.150 496.780 1172.470 496.840 ;
        RECT 1172.150 294.000 1172.470 294.060 ;
        RECT 1704.370 294.000 1704.690 294.060 ;
        RECT 1172.150 293.860 1704.690 294.000 ;
        RECT 1172.150 293.800 1172.470 293.860 ;
        RECT 1704.370 293.800 1704.690 293.860 ;
      LAYER via ;
        RECT 1166.200 496.780 1166.460 497.040 ;
        RECT 1172.180 496.780 1172.440 497.040 ;
        RECT 1172.180 293.800 1172.440 294.060 ;
        RECT 1704.400 293.800 1704.660 294.060 ;
      LAYER met2 ;
        RECT 1166.330 510.340 1166.610 514.000 ;
        RECT 1166.260 510.000 1166.610 510.340 ;
        RECT 1166.260 497.070 1166.400 510.000 ;
        RECT 1166.200 496.750 1166.460 497.070 ;
        RECT 1172.180 496.750 1172.440 497.070 ;
        RECT 1172.240 294.090 1172.380 496.750 ;
        RECT 1172.180 293.770 1172.440 294.090 ;
        RECT 1704.400 293.770 1704.660 294.090 ;
        RECT 1704.460 17.410 1704.600 293.770 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.510 300.460 1179.830 300.520 ;
        RECT 1725.070 300.460 1725.390 300.520 ;
        RECT 1179.510 300.320 1725.390 300.460 ;
        RECT 1179.510 300.260 1179.830 300.320 ;
        RECT 1725.070 300.260 1725.390 300.320 ;
      LAYER via ;
        RECT 1179.540 300.260 1179.800 300.520 ;
        RECT 1725.100 300.260 1725.360 300.520 ;
      LAYER met2 ;
        RECT 1178.750 510.410 1179.030 514.000 ;
        RECT 1178.750 510.270 1179.740 510.410 ;
        RECT 1178.750 510.000 1179.030 510.270 ;
        RECT 1179.600 300.550 1179.740 510.270 ;
        RECT 1179.540 300.230 1179.800 300.550 ;
        RECT 1725.100 300.230 1725.360 300.550 ;
        RECT 1725.160 17.410 1725.300 300.230 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1231.490 500.720 1231.810 500.780 ;
        RECT 1221.000 500.580 1231.810 500.720 ;
        RECT 1191.010 500.380 1191.330 500.440 ;
        RECT 1221.000 500.380 1221.140 500.580 ;
        RECT 1231.490 500.520 1231.810 500.580 ;
        RECT 1191.010 500.240 1221.140 500.380 ;
        RECT 1191.010 500.180 1191.330 500.240 ;
        RECT 1231.490 51.580 1231.810 51.640 ;
        RECT 1739.330 51.580 1739.650 51.640 ;
        RECT 1231.490 51.440 1739.650 51.580 ;
        RECT 1231.490 51.380 1231.810 51.440 ;
        RECT 1739.330 51.380 1739.650 51.440 ;
        RECT 1739.330 20.980 1739.650 21.040 ;
        RECT 1745.310 20.980 1745.630 21.040 ;
        RECT 1739.330 20.840 1745.630 20.980 ;
        RECT 1739.330 20.780 1739.650 20.840 ;
        RECT 1745.310 20.780 1745.630 20.840 ;
      LAYER via ;
        RECT 1191.040 500.180 1191.300 500.440 ;
        RECT 1231.520 500.520 1231.780 500.780 ;
        RECT 1231.520 51.380 1231.780 51.640 ;
        RECT 1739.360 51.380 1739.620 51.640 ;
        RECT 1739.360 20.780 1739.620 21.040 ;
        RECT 1745.340 20.780 1745.600 21.040 ;
      LAYER met2 ;
        RECT 1191.170 510.340 1191.450 514.000 ;
        RECT 1191.100 510.000 1191.450 510.340 ;
        RECT 1191.100 500.470 1191.240 510.000 ;
        RECT 1231.520 500.490 1231.780 500.810 ;
        RECT 1191.040 500.150 1191.300 500.470 ;
        RECT 1231.580 51.670 1231.720 500.490 ;
        RECT 1231.520 51.350 1231.780 51.670 ;
        RECT 1739.360 51.350 1739.620 51.670 ;
        RECT 1739.420 21.070 1739.560 51.350 ;
        RECT 1739.360 20.750 1739.620 21.070 ;
        RECT 1745.340 20.750 1745.600 21.070 ;
        RECT 1745.400 2.400 1745.540 20.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1203.430 500.720 1203.750 500.780 ;
        RECT 1207.110 500.720 1207.430 500.780 ;
        RECT 1203.430 500.580 1207.430 500.720 ;
        RECT 1203.430 500.520 1203.750 500.580 ;
        RECT 1207.110 500.520 1207.430 500.580 ;
        RECT 1207.110 59.060 1207.430 59.120 ;
        RECT 1759.570 59.060 1759.890 59.120 ;
        RECT 1207.110 58.920 1759.890 59.060 ;
        RECT 1207.110 58.860 1207.430 58.920 ;
        RECT 1759.570 58.860 1759.890 58.920 ;
      LAYER via ;
        RECT 1203.460 500.520 1203.720 500.780 ;
        RECT 1207.140 500.520 1207.400 500.780 ;
        RECT 1207.140 58.860 1207.400 59.120 ;
        RECT 1759.600 58.860 1759.860 59.120 ;
      LAYER met2 ;
        RECT 1203.590 510.340 1203.870 514.000 ;
        RECT 1203.520 510.000 1203.870 510.340 ;
        RECT 1203.520 500.810 1203.660 510.000 ;
        RECT 1203.460 500.490 1203.720 500.810 ;
        RECT 1207.140 500.490 1207.400 500.810 ;
        RECT 1207.200 59.150 1207.340 500.490 ;
        RECT 1207.140 58.830 1207.400 59.150 ;
        RECT 1759.600 58.830 1759.860 59.150 ;
        RECT 1759.660 17.410 1759.800 58.830 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1215.390 503.440 1215.710 503.500 ;
        RECT 1220.450 503.440 1220.770 503.500 ;
        RECT 1215.390 503.300 1220.770 503.440 ;
        RECT 1215.390 503.240 1215.710 503.300 ;
        RECT 1220.450 503.240 1220.770 503.300 ;
        RECT 1220.450 369.140 1220.770 369.200 ;
        RECT 1780.270 369.140 1780.590 369.200 ;
        RECT 1220.450 369.000 1780.590 369.140 ;
        RECT 1220.450 368.940 1220.770 369.000 ;
        RECT 1780.270 368.940 1780.590 369.000 ;
      LAYER via ;
        RECT 1215.420 503.240 1215.680 503.500 ;
        RECT 1220.480 503.240 1220.740 503.500 ;
        RECT 1220.480 368.940 1220.740 369.200 ;
        RECT 1780.300 368.940 1780.560 369.200 ;
      LAYER met2 ;
        RECT 1215.550 510.340 1215.830 514.000 ;
        RECT 1215.480 510.000 1215.830 510.340 ;
        RECT 1215.480 503.530 1215.620 510.000 ;
        RECT 1215.420 503.210 1215.680 503.530 ;
        RECT 1220.480 503.210 1220.740 503.530 ;
        RECT 1220.540 369.230 1220.680 503.210 ;
        RECT 1220.480 368.910 1220.740 369.230 ;
        RECT 1780.300 368.910 1780.560 369.230 ;
        RECT 1780.360 17.410 1780.500 368.910 ;
        RECT 1780.360 17.270 1780.960 17.410 ;
        RECT 1780.820 2.400 1780.960 17.270 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.350 375.940 1227.670 376.000 ;
        RECT 1794.070 375.940 1794.390 376.000 ;
        RECT 1227.350 375.800 1794.390 375.940 ;
        RECT 1227.350 375.740 1227.670 375.800 ;
        RECT 1794.070 375.740 1794.390 375.800 ;
      LAYER via ;
        RECT 1227.380 375.740 1227.640 376.000 ;
        RECT 1794.100 375.740 1794.360 376.000 ;
      LAYER met2 ;
        RECT 1227.970 510.410 1228.250 514.000 ;
        RECT 1227.440 510.270 1228.250 510.410 ;
        RECT 1227.440 376.030 1227.580 510.270 ;
        RECT 1227.970 510.000 1228.250 510.270 ;
        RECT 1227.380 375.710 1227.640 376.030 ;
        RECT 1794.100 375.710 1794.360 376.030 ;
        RECT 1794.160 17.410 1794.300 375.710 ;
        RECT 1794.160 17.270 1798.900 17.410 ;
        RECT 1798.760 2.400 1798.900 17.270 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 65.520 1241.930 65.580 ;
        RECT 1814.770 65.520 1815.090 65.580 ;
        RECT 1241.610 65.380 1815.090 65.520 ;
        RECT 1241.610 65.320 1241.930 65.380 ;
        RECT 1814.770 65.320 1815.090 65.380 ;
      LAYER via ;
        RECT 1241.640 65.320 1241.900 65.580 ;
        RECT 1814.800 65.320 1815.060 65.580 ;
      LAYER met2 ;
        RECT 1240.390 510.410 1240.670 514.000 ;
        RECT 1240.390 510.270 1241.840 510.410 ;
        RECT 1240.390 510.000 1240.670 510.270 ;
        RECT 1241.700 65.610 1241.840 510.270 ;
        RECT 1241.640 65.290 1241.900 65.610 ;
        RECT 1814.800 65.290 1815.060 65.610 ;
        RECT 1814.860 17.410 1815.000 65.290 ;
        RECT 1814.860 17.270 1816.840 17.410 ;
        RECT 1816.700 2.400 1816.840 17.270 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1255.410 72.320 1255.730 72.380 ;
        RECT 1829.030 72.320 1829.350 72.380 ;
        RECT 1255.410 72.180 1829.350 72.320 ;
        RECT 1255.410 72.120 1255.730 72.180 ;
        RECT 1829.030 72.120 1829.350 72.180 ;
      LAYER via ;
        RECT 1255.440 72.120 1255.700 72.380 ;
        RECT 1829.060 72.120 1829.320 72.380 ;
      LAYER met2 ;
        RECT 1252.810 510.410 1253.090 514.000 ;
        RECT 1252.810 510.270 1255.640 510.410 ;
        RECT 1252.810 510.000 1253.090 510.270 ;
        RECT 1255.500 72.410 1255.640 510.270 ;
        RECT 1255.440 72.090 1255.700 72.410 ;
        RECT 1829.060 72.090 1829.320 72.410 ;
        RECT 1829.120 17.410 1829.260 72.090 ;
        RECT 1829.120 17.270 1834.780 17.410 ;
        RECT 1834.640 2.400 1834.780 17.270 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.070 496.980 1265.390 497.040 ;
        RECT 1272.890 496.980 1273.210 497.040 ;
        RECT 1265.070 496.840 1273.210 496.980 ;
        RECT 1265.070 496.780 1265.390 496.840 ;
        RECT 1272.890 496.780 1273.210 496.840 ;
        RECT 1272.890 383.080 1273.210 383.140 ;
        RECT 1849.270 383.080 1849.590 383.140 ;
        RECT 1272.890 382.940 1849.590 383.080 ;
        RECT 1272.890 382.880 1273.210 382.940 ;
        RECT 1849.270 382.880 1849.590 382.940 ;
      LAYER via ;
        RECT 1265.100 496.780 1265.360 497.040 ;
        RECT 1272.920 496.780 1273.180 497.040 ;
        RECT 1272.920 382.880 1273.180 383.140 ;
        RECT 1849.300 382.880 1849.560 383.140 ;
      LAYER met2 ;
        RECT 1265.230 510.340 1265.510 514.000 ;
        RECT 1265.160 510.000 1265.510 510.340 ;
        RECT 1265.160 497.070 1265.300 510.000 ;
        RECT 1265.100 496.750 1265.360 497.070 ;
        RECT 1272.920 496.750 1273.180 497.070 ;
        RECT 1272.980 383.170 1273.120 496.750 ;
        RECT 1272.920 382.850 1273.180 383.170 ;
        RECT 1849.300 382.850 1849.560 383.170 ;
        RECT 1849.360 17.410 1849.500 382.850 ;
        RECT 1849.360 17.270 1852.260 17.410 ;
        RECT 1852.120 2.400 1852.260 17.270 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.490 500.720 1277.810 500.780 ;
        RECT 1307.390 500.720 1307.710 500.780 ;
        RECT 1277.490 500.580 1307.710 500.720 ;
        RECT 1277.490 500.520 1277.810 500.580 ;
        RECT 1307.390 500.520 1307.710 500.580 ;
        RECT 1307.390 79.460 1307.710 79.520 ;
        RECT 1870.430 79.460 1870.750 79.520 ;
        RECT 1307.390 79.320 1870.750 79.460 ;
        RECT 1307.390 79.260 1307.710 79.320 ;
        RECT 1870.430 79.260 1870.750 79.320 ;
      LAYER via ;
        RECT 1277.520 500.520 1277.780 500.780 ;
        RECT 1307.420 500.520 1307.680 500.780 ;
        RECT 1307.420 79.260 1307.680 79.520 ;
        RECT 1870.460 79.260 1870.720 79.520 ;
      LAYER met2 ;
        RECT 1277.650 510.340 1277.930 514.000 ;
        RECT 1277.580 510.000 1277.930 510.340 ;
        RECT 1277.580 500.810 1277.720 510.000 ;
        RECT 1277.520 500.490 1277.780 500.810 ;
        RECT 1307.420 500.490 1307.680 500.810 ;
        RECT 1307.480 79.550 1307.620 500.490 ;
        RECT 1307.420 79.230 1307.680 79.550 ;
        RECT 1870.460 79.230 1870.720 79.550 ;
        RECT 1870.520 7.210 1870.660 79.230 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 498.250 503.440 498.570 503.500 ;
        RECT 502.850 503.440 503.170 503.500 ;
        RECT 498.250 503.300 503.170 503.440 ;
        RECT 498.250 503.240 498.570 503.300 ;
        RECT 502.850 503.240 503.170 503.300 ;
        RECT 502.850 265.440 503.170 265.500 ;
        RECT 745.270 265.440 745.590 265.500 ;
        RECT 502.850 265.300 745.590 265.440 ;
        RECT 502.850 265.240 503.170 265.300 ;
        RECT 745.270 265.240 745.590 265.300 ;
      LAYER via ;
        RECT 498.280 503.240 498.540 503.500 ;
        RECT 502.880 503.240 503.140 503.500 ;
        RECT 502.880 265.240 503.140 265.500 ;
        RECT 745.300 265.240 745.560 265.500 ;
      LAYER met2 ;
        RECT 498.410 510.340 498.690 514.000 ;
        RECT 498.340 510.000 498.690 510.340 ;
        RECT 498.340 503.530 498.480 510.000 ;
        RECT 498.280 503.210 498.540 503.530 ;
        RECT 502.880 503.210 503.140 503.530 ;
        RECT 502.940 265.530 503.080 503.210 ;
        RECT 502.880 265.210 503.140 265.530 ;
        RECT 745.300 265.210 745.560 265.530 ;
        RECT 745.360 16.900 745.500 265.210 ;
        RECT 745.360 16.760 746.420 16.900 ;
        RECT 746.280 2.400 746.420 16.760 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1289.910 86.940 1290.230 87.000 ;
        RECT 1883.770 86.940 1884.090 87.000 ;
        RECT 1289.910 86.800 1884.090 86.940 ;
        RECT 1289.910 86.740 1290.230 86.800 ;
        RECT 1883.770 86.740 1884.090 86.800 ;
      LAYER via ;
        RECT 1289.940 86.740 1290.200 87.000 ;
        RECT 1883.800 86.740 1884.060 87.000 ;
      LAYER met2 ;
        RECT 1290.070 510.340 1290.350 514.000 ;
        RECT 1290.000 510.000 1290.350 510.340 ;
        RECT 1290.000 87.030 1290.140 510.000 ;
        RECT 1289.940 86.710 1290.200 87.030 ;
        RECT 1883.800 86.710 1884.060 87.030 ;
        RECT 1883.860 17.410 1884.000 86.710 ;
        RECT 1883.860 17.270 1888.140 17.410 ;
        RECT 1888.000 2.400 1888.140 17.270 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.250 389.880 1303.570 389.940 ;
        RECT 1904.470 389.880 1904.790 389.940 ;
        RECT 1303.250 389.740 1904.790 389.880 ;
        RECT 1303.250 389.680 1303.570 389.740 ;
        RECT 1904.470 389.680 1904.790 389.740 ;
      LAYER via ;
        RECT 1303.280 389.680 1303.540 389.940 ;
        RECT 1904.500 389.680 1904.760 389.940 ;
      LAYER met2 ;
        RECT 1302.490 510.410 1302.770 514.000 ;
        RECT 1302.490 510.270 1303.480 510.410 ;
        RECT 1302.490 510.000 1302.770 510.270 ;
        RECT 1303.340 389.970 1303.480 510.270 ;
        RECT 1303.280 389.650 1303.540 389.970 ;
        RECT 1904.500 389.650 1904.760 389.970 ;
        RECT 1904.560 17.410 1904.700 389.650 ;
        RECT 1904.560 17.270 1906.080 17.410 ;
        RECT 1905.940 2.400 1906.080 17.270 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.510 396.680 1317.830 396.740 ;
        RECT 1918.270 396.680 1918.590 396.740 ;
        RECT 1317.510 396.540 1918.590 396.680 ;
        RECT 1317.510 396.480 1317.830 396.540 ;
        RECT 1918.270 396.480 1918.590 396.540 ;
      LAYER via ;
        RECT 1317.540 396.480 1317.800 396.740 ;
        RECT 1918.300 396.480 1918.560 396.740 ;
      LAYER met2 ;
        RECT 1314.910 510.410 1315.190 514.000 ;
        RECT 1314.910 510.270 1317.740 510.410 ;
        RECT 1314.910 510.000 1315.190 510.270 ;
        RECT 1317.600 396.770 1317.740 510.270 ;
        RECT 1317.540 396.450 1317.800 396.770 ;
        RECT 1918.300 396.450 1918.560 396.770 ;
        RECT 1918.360 17.410 1918.500 396.450 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1326.710 502.080 1327.030 502.140 ;
        RECT 1330.850 502.080 1331.170 502.140 ;
        RECT 1326.710 501.940 1331.170 502.080 ;
        RECT 1326.710 501.880 1327.030 501.940 ;
        RECT 1330.850 501.880 1331.170 501.940 ;
        RECT 1330.850 404.160 1331.170 404.220 ;
        RECT 1938.970 404.160 1939.290 404.220 ;
        RECT 1330.850 404.020 1939.290 404.160 ;
        RECT 1330.850 403.960 1331.170 404.020 ;
        RECT 1938.970 403.960 1939.290 404.020 ;
      LAYER via ;
        RECT 1326.740 501.880 1327.000 502.140 ;
        RECT 1330.880 501.880 1331.140 502.140 ;
        RECT 1330.880 403.960 1331.140 404.220 ;
        RECT 1939.000 403.960 1939.260 404.220 ;
      LAYER met2 ;
        RECT 1326.870 510.340 1327.150 514.000 ;
        RECT 1326.800 510.000 1327.150 510.340 ;
        RECT 1326.800 502.170 1326.940 510.000 ;
        RECT 1326.740 501.850 1327.000 502.170 ;
        RECT 1330.880 501.850 1331.140 502.170 ;
        RECT 1330.940 404.250 1331.080 501.850 ;
        RECT 1330.880 403.930 1331.140 404.250 ;
        RECT 1939.000 403.930 1939.260 404.250 ;
        RECT 1939.060 17.410 1939.200 403.930 ;
        RECT 1939.060 17.270 1941.500 17.410 ;
        RECT 1941.360 2.400 1941.500 17.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1339.130 503.440 1339.450 503.500 ;
        RECT 1345.110 503.440 1345.430 503.500 ;
        RECT 1339.130 503.300 1345.430 503.440 ;
        RECT 1339.130 503.240 1339.450 503.300 ;
        RECT 1345.110 503.240 1345.430 503.300 ;
        RECT 1345.110 93.400 1345.430 93.460 ;
        RECT 1953.230 93.400 1953.550 93.460 ;
        RECT 1345.110 93.260 1953.550 93.400 ;
        RECT 1345.110 93.200 1345.430 93.260 ;
        RECT 1953.230 93.200 1953.550 93.260 ;
        RECT 1953.230 16.900 1953.550 16.960 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 1953.230 16.760 1959.530 16.900 ;
        RECT 1953.230 16.700 1953.550 16.760 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
      LAYER via ;
        RECT 1339.160 503.240 1339.420 503.500 ;
        RECT 1345.140 503.240 1345.400 503.500 ;
        RECT 1345.140 93.200 1345.400 93.460 ;
        RECT 1953.260 93.200 1953.520 93.460 ;
        RECT 1953.260 16.700 1953.520 16.960 ;
        RECT 1959.240 16.700 1959.500 16.960 ;
      LAYER met2 ;
        RECT 1339.290 510.340 1339.570 514.000 ;
        RECT 1339.220 510.000 1339.570 510.340 ;
        RECT 1339.220 503.530 1339.360 510.000 ;
        RECT 1339.160 503.210 1339.420 503.530 ;
        RECT 1345.140 503.210 1345.400 503.530 ;
        RECT 1345.200 93.490 1345.340 503.210 ;
        RECT 1345.140 93.170 1345.400 93.490 ;
        RECT 1953.260 93.170 1953.520 93.490 ;
        RECT 1953.320 16.990 1953.460 93.170 ;
        RECT 1953.260 16.670 1953.520 16.990 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 1959.300 2.400 1959.440 16.670 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 203.900 1352.330 203.960 ;
        RECT 1973.470 203.900 1973.790 203.960 ;
        RECT 1352.010 203.760 1973.790 203.900 ;
        RECT 1352.010 203.700 1352.330 203.760 ;
        RECT 1973.470 203.700 1973.790 203.760 ;
      LAYER via ;
        RECT 1352.040 203.700 1352.300 203.960 ;
        RECT 1973.500 203.700 1973.760 203.960 ;
      LAYER met2 ;
        RECT 1351.710 510.340 1351.990 514.000 ;
        RECT 1351.640 510.000 1351.990 510.340 ;
        RECT 1351.640 503.610 1351.780 510.000 ;
        RECT 1351.640 503.470 1352.240 503.610 ;
        RECT 1352.100 203.990 1352.240 503.470 ;
        RECT 1352.040 203.670 1352.300 203.990 ;
        RECT 1973.500 203.670 1973.760 203.990 ;
        RECT 1973.560 17.410 1973.700 203.670 ;
        RECT 1973.560 17.270 1977.380 17.410 ;
        RECT 1977.240 2.400 1977.380 17.270 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.350 417.760 1365.670 417.820 ;
        RECT 1994.170 417.760 1994.490 417.820 ;
        RECT 1365.350 417.620 1994.490 417.760 ;
        RECT 1365.350 417.560 1365.670 417.620 ;
        RECT 1994.170 417.560 1994.490 417.620 ;
      LAYER via ;
        RECT 1365.380 417.560 1365.640 417.820 ;
        RECT 1994.200 417.560 1994.460 417.820 ;
      LAYER met2 ;
        RECT 1364.130 510.410 1364.410 514.000 ;
        RECT 1364.130 510.270 1365.580 510.410 ;
        RECT 1364.130 510.000 1364.410 510.270 ;
        RECT 1365.440 417.850 1365.580 510.270 ;
        RECT 1365.380 417.530 1365.640 417.850 ;
        RECT 1994.200 417.530 1994.460 417.850 ;
        RECT 1994.260 17.410 1994.400 417.530 ;
        RECT 1994.260 17.270 1995.320 17.410 ;
        RECT 1995.180 2.400 1995.320 17.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1379.610 424.900 1379.930 424.960 ;
        RECT 2007.970 424.900 2008.290 424.960 ;
        RECT 1379.610 424.760 2008.290 424.900 ;
        RECT 1379.610 424.700 1379.930 424.760 ;
        RECT 2007.970 424.700 2008.290 424.760 ;
      LAYER via ;
        RECT 1379.640 424.700 1379.900 424.960 ;
        RECT 2008.000 424.700 2008.260 424.960 ;
      LAYER met2 ;
        RECT 1376.550 510.410 1376.830 514.000 ;
        RECT 1376.550 510.270 1379.840 510.410 ;
        RECT 1376.550 510.000 1376.830 510.270 ;
        RECT 1379.700 424.990 1379.840 510.270 ;
        RECT 1379.640 424.670 1379.900 424.990 ;
        RECT 2008.000 424.670 2008.260 424.990 ;
        RECT 2008.060 17.410 2008.200 424.670 ;
        RECT 2008.060 17.270 2012.800 17.410 ;
        RECT 2012.660 2.400 2012.800 17.270 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.810 473.180 1389.130 473.240 ;
        RECT 2028.670 473.180 2028.990 473.240 ;
        RECT 1388.810 473.040 2028.990 473.180 ;
        RECT 1388.810 472.980 1389.130 473.040 ;
        RECT 2028.670 472.980 2028.990 473.040 ;
      LAYER via ;
        RECT 1388.840 472.980 1389.100 473.240 ;
        RECT 2028.700 472.980 2028.960 473.240 ;
      LAYER met2 ;
        RECT 1388.970 510.340 1389.250 514.000 ;
        RECT 1388.900 510.000 1389.250 510.340 ;
        RECT 1388.900 473.270 1389.040 510.000 ;
        RECT 1388.840 472.950 1389.100 473.270 ;
        RECT 2028.700 472.950 2028.960 473.270 ;
        RECT 2028.760 17.410 2028.900 472.950 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1401.230 500.720 1401.550 500.780 ;
        RECT 1406.750 500.720 1407.070 500.780 ;
        RECT 1401.230 500.580 1407.070 500.720 ;
        RECT 1401.230 500.520 1401.550 500.580 ;
        RECT 1406.750 500.520 1407.070 500.580 ;
        RECT 1406.750 431.700 1407.070 431.760 ;
        RECT 2042.470 431.700 2042.790 431.760 ;
        RECT 1406.750 431.560 2042.790 431.700 ;
        RECT 1406.750 431.500 1407.070 431.560 ;
        RECT 2042.470 431.500 2042.790 431.560 ;
        RECT 2042.470 20.980 2042.790 21.040 ;
        RECT 2048.450 20.980 2048.770 21.040 ;
        RECT 2042.470 20.840 2048.770 20.980 ;
        RECT 2042.470 20.780 2042.790 20.840 ;
        RECT 2048.450 20.780 2048.770 20.840 ;
      LAYER via ;
        RECT 1401.260 500.520 1401.520 500.780 ;
        RECT 1406.780 500.520 1407.040 500.780 ;
        RECT 1406.780 431.500 1407.040 431.760 ;
        RECT 2042.500 431.500 2042.760 431.760 ;
        RECT 2042.500 20.780 2042.760 21.040 ;
        RECT 2048.480 20.780 2048.740 21.040 ;
      LAYER met2 ;
        RECT 1401.390 510.340 1401.670 514.000 ;
        RECT 1401.320 510.000 1401.670 510.340 ;
        RECT 1401.320 500.810 1401.460 510.000 ;
        RECT 1401.260 500.490 1401.520 500.810 ;
        RECT 1406.780 500.490 1407.040 500.810 ;
        RECT 1406.840 431.790 1406.980 500.490 ;
        RECT 1406.780 431.470 1407.040 431.790 ;
        RECT 2042.500 431.470 2042.760 431.790 ;
        RECT 2042.560 21.070 2042.700 431.470 ;
        RECT 2042.500 20.750 2042.760 21.070 ;
        RECT 2048.480 20.750 2048.740 21.070 ;
        RECT 2048.540 2.400 2048.680 20.750 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.670 503.440 510.990 503.500 ;
        RECT 516.650 503.440 516.970 503.500 ;
        RECT 510.670 503.300 516.970 503.440 ;
        RECT 510.670 503.240 510.990 503.300 ;
        RECT 516.650 503.240 516.970 503.300 ;
        RECT 516.650 279.380 516.970 279.440 ;
        RECT 759.070 279.380 759.390 279.440 ;
        RECT 516.650 279.240 759.390 279.380 ;
        RECT 516.650 279.180 516.970 279.240 ;
        RECT 759.070 279.180 759.390 279.240 ;
      LAYER via ;
        RECT 510.700 503.240 510.960 503.500 ;
        RECT 516.680 503.240 516.940 503.500 ;
        RECT 516.680 279.180 516.940 279.440 ;
        RECT 759.100 279.180 759.360 279.440 ;
      LAYER met2 ;
        RECT 510.830 510.340 511.110 514.000 ;
        RECT 510.760 510.000 511.110 510.340 ;
        RECT 510.760 503.530 510.900 510.000 ;
        RECT 510.700 503.210 510.960 503.530 ;
        RECT 516.680 503.210 516.940 503.530 ;
        RECT 516.740 279.470 516.880 503.210 ;
        RECT 516.680 279.150 516.940 279.470 ;
        RECT 759.100 279.150 759.360 279.470 ;
        RECT 759.160 17.410 759.300 279.150 ;
        RECT 759.160 17.270 763.900 17.410 ;
        RECT 763.760 2.400 763.900 17.270 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1413.650 445.640 1413.970 445.700 ;
        RECT 2063.170 445.640 2063.490 445.700 ;
        RECT 1413.650 445.500 2063.490 445.640 ;
        RECT 1413.650 445.440 1413.970 445.500 ;
        RECT 2063.170 445.440 2063.490 445.500 ;
      LAYER via ;
        RECT 1413.680 445.440 1413.940 445.700 ;
        RECT 2063.200 445.440 2063.460 445.700 ;
      LAYER met2 ;
        RECT 1413.810 510.340 1414.090 514.000 ;
        RECT 1413.740 510.000 1414.090 510.340 ;
        RECT 1413.740 445.730 1413.880 510.000 ;
        RECT 1413.680 445.410 1413.940 445.730 ;
        RECT 2063.200 445.410 2063.460 445.730 ;
        RECT 2063.260 17.410 2063.400 445.410 ;
        RECT 2063.260 17.270 2066.620 17.410 ;
        RECT 2066.480 2.400 2066.620 17.270 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1427.450 452.100 1427.770 452.160 ;
        RECT 2083.870 452.100 2084.190 452.160 ;
        RECT 1427.450 451.960 2084.190 452.100 ;
        RECT 1427.450 451.900 1427.770 451.960 ;
        RECT 2083.870 451.900 2084.190 451.960 ;
      LAYER via ;
        RECT 1427.480 451.900 1427.740 452.160 ;
        RECT 2083.900 451.900 2084.160 452.160 ;
      LAYER met2 ;
        RECT 1426.230 510.410 1426.510 514.000 ;
        RECT 1426.230 510.270 1427.680 510.410 ;
        RECT 1426.230 510.000 1426.510 510.270 ;
        RECT 1427.540 452.190 1427.680 510.270 ;
        RECT 1427.480 451.870 1427.740 452.190 ;
        RECT 2083.900 451.870 2084.160 452.190 ;
        RECT 2083.960 17.410 2084.100 451.870 ;
        RECT 2083.960 17.270 2084.560 17.410 ;
        RECT 2084.420 2.400 2084.560 17.270 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1438.030 496.980 1438.350 497.040 ;
        RECT 1441.710 496.980 1442.030 497.040 ;
        RECT 1438.030 496.840 1442.030 496.980 ;
        RECT 1438.030 496.780 1438.350 496.840 ;
        RECT 1441.710 496.780 1442.030 496.840 ;
        RECT 1441.710 148.140 1442.030 148.200 ;
        RECT 2097.670 148.140 2097.990 148.200 ;
        RECT 1441.710 148.000 2097.990 148.140 ;
        RECT 1441.710 147.940 1442.030 148.000 ;
        RECT 2097.670 147.940 2097.990 148.000 ;
      LAYER via ;
        RECT 1438.060 496.780 1438.320 497.040 ;
        RECT 1441.740 496.780 1442.000 497.040 ;
        RECT 1441.740 147.940 1442.000 148.200 ;
        RECT 2097.700 147.940 2097.960 148.200 ;
      LAYER met2 ;
        RECT 1438.190 510.340 1438.470 514.000 ;
        RECT 1438.120 510.000 1438.470 510.340 ;
        RECT 1438.120 497.070 1438.260 510.000 ;
        RECT 1438.060 496.750 1438.320 497.070 ;
        RECT 1441.740 496.750 1442.000 497.070 ;
        RECT 1441.800 148.230 1441.940 496.750 ;
        RECT 1441.740 147.910 1442.000 148.230 ;
        RECT 2097.700 147.910 2097.960 148.230 ;
        RECT 2097.760 18.090 2097.900 147.910 ;
        RECT 2097.760 17.950 2102.040 18.090 ;
        RECT 2101.900 2.400 2102.040 17.950 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1450.450 496.980 1450.770 497.040 ;
        RECT 1455.050 496.980 1455.370 497.040 ;
        RECT 1450.450 496.840 1455.370 496.980 ;
        RECT 1450.450 496.780 1450.770 496.840 ;
        RECT 1455.050 496.780 1455.370 496.840 ;
        RECT 1455.050 459.240 1455.370 459.300 ;
        RECT 2118.370 459.240 2118.690 459.300 ;
        RECT 1455.050 459.100 2118.690 459.240 ;
        RECT 1455.050 459.040 1455.370 459.100 ;
        RECT 2118.370 459.040 2118.690 459.100 ;
      LAYER via ;
        RECT 1450.480 496.780 1450.740 497.040 ;
        RECT 1455.080 496.780 1455.340 497.040 ;
        RECT 1455.080 459.040 1455.340 459.300 ;
        RECT 2118.400 459.040 2118.660 459.300 ;
      LAYER met2 ;
        RECT 1450.610 510.340 1450.890 514.000 ;
        RECT 1450.540 510.000 1450.890 510.340 ;
        RECT 1450.540 497.070 1450.680 510.000 ;
        RECT 1450.480 496.750 1450.740 497.070 ;
        RECT 1455.080 496.750 1455.340 497.070 ;
        RECT 1455.140 459.330 1455.280 496.750 ;
        RECT 1455.080 459.010 1455.340 459.330 ;
        RECT 2118.400 459.010 2118.660 459.330 ;
        RECT 2118.460 17.410 2118.600 459.010 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1462.870 500.040 1463.190 500.100 ;
        RECT 1500.590 500.040 1500.910 500.100 ;
        RECT 1462.870 499.900 1500.910 500.040 ;
        RECT 1462.870 499.840 1463.190 499.900 ;
        RECT 1500.590 499.840 1500.910 499.900 ;
        RECT 1500.590 369.480 1500.910 369.540 ;
        RECT 2132.170 369.480 2132.490 369.540 ;
        RECT 1500.590 369.340 2132.490 369.480 ;
        RECT 1500.590 369.280 1500.910 369.340 ;
        RECT 2132.170 369.280 2132.490 369.340 ;
      LAYER via ;
        RECT 1462.900 499.840 1463.160 500.100 ;
        RECT 1500.620 499.840 1500.880 500.100 ;
        RECT 1500.620 369.280 1500.880 369.540 ;
        RECT 2132.200 369.280 2132.460 369.540 ;
      LAYER met2 ;
        RECT 1463.030 510.340 1463.310 514.000 ;
        RECT 1462.960 510.000 1463.310 510.340 ;
        RECT 1462.960 500.130 1463.100 510.000 ;
        RECT 1462.900 499.810 1463.160 500.130 ;
        RECT 1500.620 499.810 1500.880 500.130 ;
        RECT 1500.680 369.570 1500.820 499.810 ;
        RECT 1500.620 369.250 1500.880 369.570 ;
        RECT 2132.200 369.250 2132.460 369.570 ;
        RECT 2132.260 17.410 2132.400 369.250 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1475.290 466.040 1475.610 466.100 ;
        RECT 2152.870 466.040 2153.190 466.100 ;
        RECT 1475.290 465.900 2153.190 466.040 ;
        RECT 1475.290 465.840 1475.610 465.900 ;
        RECT 2152.870 465.840 2153.190 465.900 ;
      LAYER via ;
        RECT 1475.320 465.840 1475.580 466.100 ;
        RECT 2152.900 465.840 2153.160 466.100 ;
      LAYER met2 ;
        RECT 1475.450 510.340 1475.730 514.000 ;
        RECT 1475.380 510.000 1475.730 510.340 ;
        RECT 1475.380 466.130 1475.520 510.000 ;
        RECT 1475.320 465.810 1475.580 466.130 ;
        RECT 2152.900 465.810 2153.160 466.130 ;
        RECT 2152.960 17.410 2153.100 465.810 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1490.010 24.040 1490.330 24.100 ;
        RECT 2173.110 24.040 2173.430 24.100 ;
        RECT 1490.010 23.900 2173.430 24.040 ;
        RECT 1490.010 23.840 1490.330 23.900 ;
        RECT 2173.110 23.840 2173.430 23.900 ;
      LAYER via ;
        RECT 1490.040 23.840 1490.300 24.100 ;
        RECT 2173.140 23.840 2173.400 24.100 ;
      LAYER met2 ;
        RECT 1487.870 510.410 1488.150 514.000 ;
        RECT 1487.870 510.270 1490.240 510.410 ;
        RECT 1487.870 510.000 1488.150 510.270 ;
        RECT 1490.100 24.130 1490.240 510.270 ;
        RECT 1490.040 23.810 1490.300 24.130 ;
        RECT 2173.140 23.810 2173.400 24.130 ;
        RECT 2173.200 2.400 2173.340 23.810 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1503.810 376.280 1504.130 376.340 ;
        RECT 2187.370 376.280 2187.690 376.340 ;
        RECT 1503.810 376.140 2187.690 376.280 ;
        RECT 1503.810 376.080 1504.130 376.140 ;
        RECT 2187.370 376.080 2187.690 376.140 ;
      LAYER via ;
        RECT 1503.840 376.080 1504.100 376.340 ;
        RECT 2187.400 376.080 2187.660 376.340 ;
      LAYER met2 ;
        RECT 1500.290 510.410 1500.570 514.000 ;
        RECT 1500.290 510.270 1504.040 510.410 ;
        RECT 1500.290 510.000 1500.570 510.270 ;
        RECT 1503.900 376.370 1504.040 510.270 ;
        RECT 1503.840 376.050 1504.100 376.370 ;
        RECT 2187.400 376.050 2187.660 376.370 ;
        RECT 2187.460 17.410 2187.600 376.050 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1512.550 497.320 1512.870 497.380 ;
        RECT 1521.290 497.320 1521.610 497.380 ;
        RECT 1512.550 497.180 1521.610 497.320 ;
        RECT 1512.550 497.120 1512.870 497.180 ;
        RECT 1521.290 497.120 1521.610 497.180 ;
        RECT 1521.290 382.740 1521.610 382.800 ;
        RECT 2208.070 382.740 2208.390 382.800 ;
        RECT 1521.290 382.600 2208.390 382.740 ;
        RECT 1521.290 382.540 1521.610 382.600 ;
        RECT 2208.070 382.540 2208.390 382.600 ;
      LAYER via ;
        RECT 1512.580 497.120 1512.840 497.380 ;
        RECT 1521.320 497.120 1521.580 497.380 ;
        RECT 1521.320 382.540 1521.580 382.800 ;
        RECT 2208.100 382.540 2208.360 382.800 ;
      LAYER met2 ;
        RECT 1512.710 510.340 1512.990 514.000 ;
        RECT 1512.640 510.000 1512.990 510.340 ;
        RECT 1512.640 497.410 1512.780 510.000 ;
        RECT 1512.580 497.090 1512.840 497.410 ;
        RECT 1521.320 497.090 1521.580 497.410 ;
        RECT 1521.380 382.830 1521.520 497.090 ;
        RECT 1521.320 382.510 1521.580 382.830 ;
        RECT 2208.100 382.510 2208.360 382.830 ;
        RECT 2208.160 17.410 2208.300 382.510 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.970 479.980 1525.290 480.040 ;
        RECT 2221.870 479.980 2222.190 480.040 ;
        RECT 1524.970 479.840 2222.190 479.980 ;
        RECT 1524.970 479.780 1525.290 479.840 ;
        RECT 2221.870 479.780 2222.190 479.840 ;
      LAYER via ;
        RECT 1525.000 479.780 1525.260 480.040 ;
        RECT 2221.900 479.780 2222.160 480.040 ;
      LAYER met2 ;
        RECT 1525.130 510.340 1525.410 514.000 ;
        RECT 1525.060 510.000 1525.410 510.340 ;
        RECT 1525.060 480.070 1525.200 510.000 ;
        RECT 1525.000 479.750 1525.260 480.070 ;
        RECT 2221.900 479.750 2222.160 480.070 ;
        RECT 2221.960 17.410 2222.100 479.750 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 523.165 386.665 523.335 410.635 ;
        RECT 522.705 338.045 522.875 386.155 ;
      LAYER mcon ;
        RECT 523.165 410.465 523.335 410.635 ;
        RECT 522.705 385.985 522.875 386.155 ;
      LAYER met1 ;
        RECT 523.090 435.100 523.410 435.160 ;
        RECT 523.550 435.100 523.870 435.160 ;
        RECT 523.090 434.960 523.870 435.100 ;
        RECT 523.090 434.900 523.410 434.960 ;
        RECT 523.550 434.900 523.870 434.960 ;
        RECT 523.090 410.620 523.410 410.680 ;
        RECT 522.895 410.480 523.410 410.620 ;
        RECT 523.090 410.420 523.410 410.480 ;
        RECT 523.090 386.820 523.410 386.880 ;
        RECT 522.895 386.680 523.410 386.820 ;
        RECT 523.090 386.620 523.410 386.680 ;
        RECT 522.630 386.140 522.950 386.200 ;
        RECT 522.435 386.000 522.950 386.140 ;
        RECT 522.630 385.940 522.950 386.000 ;
        RECT 522.645 338.200 522.935 338.245 ;
        RECT 523.090 338.200 523.410 338.260 ;
        RECT 522.645 338.060 523.410 338.200 ;
        RECT 522.645 338.015 522.935 338.060 ;
        RECT 523.090 338.000 523.410 338.060 ;
        RECT 523.090 304.200 523.410 304.260 ;
        RECT 522.720 304.060 523.410 304.200 ;
        RECT 522.720 303.580 522.860 304.060 ;
        RECT 523.090 304.000 523.410 304.060 ;
        RECT 522.630 303.320 522.950 303.580 ;
        RECT 522.630 286.180 522.950 286.240 ;
        RECT 779.770 286.180 780.090 286.240 ;
        RECT 522.630 286.040 780.090 286.180 ;
        RECT 522.630 285.980 522.950 286.040 ;
        RECT 779.770 285.980 780.090 286.040 ;
      LAYER via ;
        RECT 523.120 434.900 523.380 435.160 ;
        RECT 523.580 434.900 523.840 435.160 ;
        RECT 523.120 410.420 523.380 410.680 ;
        RECT 523.120 386.620 523.380 386.880 ;
        RECT 522.660 385.940 522.920 386.200 ;
        RECT 523.120 338.000 523.380 338.260 ;
        RECT 523.120 304.000 523.380 304.260 ;
        RECT 522.660 303.320 522.920 303.580 ;
        RECT 522.660 285.980 522.920 286.240 ;
        RECT 779.800 285.980 780.060 286.240 ;
      LAYER met2 ;
        RECT 523.250 510.410 523.530 514.000 ;
        RECT 522.720 510.270 523.530 510.410 ;
        RECT 522.720 483.325 522.860 510.270 ;
        RECT 523.250 510.000 523.530 510.270 ;
        RECT 522.650 482.955 522.930 483.325 ;
        RECT 523.570 482.955 523.850 483.325 ;
        RECT 523.640 435.190 523.780 482.955 ;
        RECT 523.120 434.870 523.380 435.190 ;
        RECT 523.580 434.870 523.840 435.190 ;
        RECT 523.180 410.710 523.320 434.870 ;
        RECT 523.120 410.390 523.380 410.710 ;
        RECT 523.120 386.650 523.380 386.910 ;
        RECT 522.720 386.590 523.380 386.650 ;
        RECT 522.720 386.510 523.320 386.590 ;
        RECT 522.720 386.230 522.860 386.510 ;
        RECT 522.660 385.910 522.920 386.230 ;
        RECT 523.120 337.970 523.380 338.290 ;
        RECT 523.180 304.290 523.320 337.970 ;
        RECT 523.120 303.970 523.380 304.290 ;
        RECT 522.660 303.290 522.920 303.610 ;
        RECT 522.720 286.270 522.860 303.290 ;
        RECT 522.660 285.950 522.920 286.270 ;
        RECT 779.800 285.950 780.060 286.270 ;
        RECT 779.860 17.410 780.000 285.950 ;
        RECT 779.860 17.270 781.840 17.410 ;
        RECT 781.700 2.400 781.840 17.270 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 522.650 483.000 522.930 483.280 ;
        RECT 523.570 483.000 523.850 483.280 ;
      LAYER met3 ;
        RECT 522.625 483.290 522.955 483.305 ;
        RECT 523.545 483.290 523.875 483.305 ;
        RECT 522.625 482.990 523.875 483.290 ;
        RECT 522.625 482.975 522.955 482.990 ;
        RECT 523.545 482.975 523.875 482.990 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1538.310 390.220 1538.630 390.280 ;
        RECT 2242.570 390.220 2242.890 390.280 ;
        RECT 1538.310 390.080 2242.890 390.220 ;
        RECT 1538.310 390.020 1538.630 390.080 ;
        RECT 2242.570 390.020 2242.890 390.080 ;
      LAYER via ;
        RECT 1538.340 390.020 1538.600 390.280 ;
        RECT 2242.600 390.020 2242.860 390.280 ;
      LAYER met2 ;
        RECT 1537.550 510.410 1537.830 514.000 ;
        RECT 1537.550 510.270 1538.540 510.410 ;
        RECT 1537.550 510.000 1537.830 510.270 ;
        RECT 1538.400 390.310 1538.540 510.270 ;
        RECT 1538.340 389.990 1538.600 390.310 ;
        RECT 2242.600 389.990 2242.860 390.310 ;
        RECT 2242.660 17.410 2242.800 389.990 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1549.350 500.040 1549.670 500.100 ;
        RECT 1721.390 500.040 1721.710 500.100 ;
        RECT 1549.350 499.900 1721.710 500.040 ;
        RECT 1549.350 499.840 1549.670 499.900 ;
        RECT 1721.390 499.840 1721.710 499.900 ;
        RECT 1721.390 80.140 1721.710 80.200 ;
        RECT 2256.830 80.140 2257.150 80.200 ;
        RECT 1721.390 80.000 2257.150 80.140 ;
        RECT 1721.390 79.940 1721.710 80.000 ;
        RECT 2256.830 79.940 2257.150 80.000 ;
      LAYER via ;
        RECT 1549.380 499.840 1549.640 500.100 ;
        RECT 1721.420 499.840 1721.680 500.100 ;
        RECT 1721.420 79.940 1721.680 80.200 ;
        RECT 2256.860 79.940 2257.120 80.200 ;
      LAYER met2 ;
        RECT 1549.510 510.340 1549.790 514.000 ;
        RECT 1549.440 510.000 1549.790 510.340 ;
        RECT 1549.440 500.130 1549.580 510.000 ;
        RECT 1549.380 499.810 1549.640 500.130 ;
        RECT 1721.420 499.810 1721.680 500.130 ;
        RECT 1721.480 80.230 1721.620 499.810 ;
        RECT 1721.420 79.910 1721.680 80.230 ;
        RECT 2256.860 79.910 2257.120 80.230 ;
        RECT 2256.920 17.410 2257.060 79.910 ;
        RECT 2256.920 17.270 2262.580 17.410 ;
        RECT 2262.440 2.400 2262.580 17.270 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1561.770 486.780 1562.090 486.840 ;
        RECT 2277.070 486.780 2277.390 486.840 ;
        RECT 1561.770 486.640 2277.390 486.780 ;
        RECT 1561.770 486.580 1562.090 486.640 ;
        RECT 2277.070 486.580 2277.390 486.640 ;
      LAYER via ;
        RECT 1561.800 486.580 1562.060 486.840 ;
        RECT 2277.100 486.580 2277.360 486.840 ;
      LAYER met2 ;
        RECT 1561.930 510.340 1562.210 514.000 ;
        RECT 1561.860 510.000 1562.210 510.340 ;
        RECT 1561.860 486.870 1562.000 510.000 ;
        RECT 1561.800 486.550 1562.060 486.870 ;
        RECT 2277.100 486.550 2277.360 486.870 ;
        RECT 2277.160 17.410 2277.300 486.550 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1574.190 496.980 1574.510 497.040 ;
        RECT 1579.250 496.980 1579.570 497.040 ;
        RECT 1574.190 496.840 1579.570 496.980 ;
        RECT 1574.190 496.780 1574.510 496.840 ;
        RECT 1579.250 496.780 1579.570 496.840 ;
        RECT 1579.250 410.960 1579.570 411.020 ;
        RECT 2298.230 410.960 2298.550 411.020 ;
        RECT 1579.250 410.820 2298.550 410.960 ;
        RECT 1579.250 410.760 1579.570 410.820 ;
        RECT 2298.230 410.760 2298.550 410.820 ;
      LAYER via ;
        RECT 1574.220 496.780 1574.480 497.040 ;
        RECT 1579.280 496.780 1579.540 497.040 ;
        RECT 1579.280 410.760 1579.540 411.020 ;
        RECT 2298.260 410.760 2298.520 411.020 ;
      LAYER met2 ;
        RECT 1574.350 510.340 1574.630 514.000 ;
        RECT 1574.280 510.000 1574.630 510.340 ;
        RECT 1574.280 497.070 1574.420 510.000 ;
        RECT 1574.220 496.750 1574.480 497.070 ;
        RECT 1579.280 496.750 1579.540 497.070 ;
        RECT 1579.340 411.050 1579.480 496.750 ;
        RECT 1579.280 410.730 1579.540 411.050 ;
        RECT 2298.260 410.730 2298.520 411.050 ;
        RECT 2298.320 2.400 2298.460 410.730 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 493.580 1586.930 493.640 ;
        RECT 2311.570 493.580 2311.890 493.640 ;
        RECT 1586.610 493.440 2311.890 493.580 ;
        RECT 1586.610 493.380 1586.930 493.440 ;
        RECT 2311.570 493.380 2311.890 493.440 ;
      LAYER via ;
        RECT 1586.640 493.380 1586.900 493.640 ;
        RECT 2311.600 493.380 2311.860 493.640 ;
      LAYER met2 ;
        RECT 1586.770 510.340 1587.050 514.000 ;
        RECT 1586.700 510.000 1587.050 510.340 ;
        RECT 1586.700 493.670 1586.840 510.000 ;
        RECT 1586.640 493.350 1586.900 493.670 ;
        RECT 2311.600 493.350 2311.860 493.670 ;
        RECT 2311.660 17.410 2311.800 493.350 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.410 99.860 1600.730 99.920 ;
        RECT 2332.270 99.860 2332.590 99.920 ;
        RECT 1600.410 99.720 2332.590 99.860 ;
        RECT 1600.410 99.660 1600.730 99.720 ;
        RECT 2332.270 99.660 2332.590 99.720 ;
      LAYER via ;
        RECT 1600.440 99.660 1600.700 99.920 ;
        RECT 2332.300 99.660 2332.560 99.920 ;
      LAYER met2 ;
        RECT 1599.190 510.410 1599.470 514.000 ;
        RECT 1599.190 510.270 1600.640 510.410 ;
        RECT 1599.190 510.000 1599.470 510.270 ;
        RECT 1600.500 99.950 1600.640 510.270 ;
        RECT 1600.440 99.630 1600.700 99.950 ;
        RECT 2332.300 99.630 2332.560 99.950 ;
        RECT 2332.360 17.410 2332.500 99.630 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1614.210 306.920 1614.530 306.980 ;
        RECT 2346.070 306.920 2346.390 306.980 ;
        RECT 1614.210 306.780 2346.390 306.920 ;
        RECT 1614.210 306.720 1614.530 306.780 ;
        RECT 2346.070 306.720 2346.390 306.780 ;
      LAYER via ;
        RECT 1614.240 306.720 1614.500 306.980 ;
        RECT 2346.100 306.720 2346.360 306.980 ;
      LAYER met2 ;
        RECT 1611.610 510.410 1611.890 514.000 ;
        RECT 1611.610 510.270 1614.440 510.410 ;
        RECT 1611.610 510.000 1611.890 510.270 ;
        RECT 1614.300 307.010 1614.440 510.270 ;
        RECT 1614.240 306.690 1614.500 307.010 ;
        RECT 2346.100 306.690 2346.360 307.010 ;
        RECT 2346.160 17.410 2346.300 306.690 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1623.870 496.980 1624.190 497.040 ;
        RECT 1631.690 496.980 1632.010 497.040 ;
        RECT 1623.870 496.840 1632.010 496.980 ;
        RECT 1623.870 496.780 1624.190 496.840 ;
        RECT 1631.690 496.780 1632.010 496.840 ;
        RECT 1631.690 107.000 1632.010 107.060 ;
        RECT 2366.770 107.000 2367.090 107.060 ;
        RECT 1631.690 106.860 2367.090 107.000 ;
        RECT 1631.690 106.800 1632.010 106.860 ;
        RECT 2366.770 106.800 2367.090 106.860 ;
      LAYER via ;
        RECT 1623.900 496.780 1624.160 497.040 ;
        RECT 1631.720 496.780 1631.980 497.040 ;
        RECT 1631.720 106.800 1631.980 107.060 ;
        RECT 2366.800 106.800 2367.060 107.060 ;
      LAYER met2 ;
        RECT 1624.030 510.340 1624.310 514.000 ;
        RECT 1623.960 510.000 1624.310 510.340 ;
        RECT 1623.960 497.070 1624.100 510.000 ;
        RECT 1623.900 496.750 1624.160 497.070 ;
        RECT 1631.720 496.750 1631.980 497.070 ;
        RECT 1631.780 107.090 1631.920 496.750 ;
        RECT 1631.720 106.770 1631.980 107.090 ;
        RECT 2366.800 106.770 2367.060 107.090 ;
        RECT 2366.860 17.410 2367.000 106.770 ;
        RECT 2366.860 17.270 2369.760 17.410 ;
        RECT 2369.620 2.400 2369.760 17.270 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1636.290 496.980 1636.610 497.040 ;
        RECT 1641.350 496.980 1641.670 497.040 ;
        RECT 1636.290 496.840 1641.670 496.980 ;
        RECT 1636.290 496.780 1636.610 496.840 ;
        RECT 1641.350 496.780 1641.670 496.840 ;
        RECT 1641.350 182.820 1641.670 182.880 ;
        RECT 2387.930 182.820 2388.250 182.880 ;
        RECT 1641.350 182.680 2388.250 182.820 ;
        RECT 1641.350 182.620 1641.670 182.680 ;
        RECT 2387.930 182.620 2388.250 182.680 ;
      LAYER via ;
        RECT 1636.320 496.780 1636.580 497.040 ;
        RECT 1641.380 496.780 1641.640 497.040 ;
        RECT 1641.380 182.620 1641.640 182.880 ;
        RECT 2387.960 182.620 2388.220 182.880 ;
      LAYER met2 ;
        RECT 1636.450 510.340 1636.730 514.000 ;
        RECT 1636.380 510.000 1636.730 510.340 ;
        RECT 1636.380 497.070 1636.520 510.000 ;
        RECT 1636.320 496.750 1636.580 497.070 ;
        RECT 1641.380 496.750 1641.640 497.070 ;
        RECT 1641.440 182.910 1641.580 496.750 ;
        RECT 1641.380 182.590 1641.640 182.910 ;
        RECT 2387.960 182.590 2388.220 182.910 ;
        RECT 2388.020 17.410 2388.160 182.590 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1648.710 397.020 1649.030 397.080 ;
        RECT 2401.270 397.020 2401.590 397.080 ;
        RECT 1648.710 396.880 2401.590 397.020 ;
        RECT 1648.710 396.820 1649.030 396.880 ;
        RECT 2401.270 396.820 2401.590 396.880 ;
      LAYER via ;
        RECT 1648.740 396.820 1649.000 397.080 ;
        RECT 2401.300 396.820 2401.560 397.080 ;
      LAYER met2 ;
        RECT 1648.870 510.340 1649.150 514.000 ;
        RECT 1648.800 510.000 1649.150 510.340 ;
        RECT 1648.800 397.110 1648.940 510.000 ;
        RECT 1648.740 396.790 1649.000 397.110 ;
        RECT 2401.300 396.790 2401.560 397.110 ;
        RECT 2401.360 17.410 2401.500 396.790 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 293.320 538.130 293.380 ;
        RECT 793.570 293.320 793.890 293.380 ;
        RECT 537.810 293.180 793.890 293.320 ;
        RECT 537.810 293.120 538.130 293.180 ;
        RECT 793.570 293.120 793.890 293.180 ;
        RECT 793.570 17.580 793.890 17.640 ;
        RECT 799.550 17.580 799.870 17.640 ;
        RECT 793.570 17.440 799.870 17.580 ;
        RECT 793.570 17.380 793.890 17.440 ;
        RECT 799.550 17.380 799.870 17.440 ;
      LAYER via ;
        RECT 537.840 293.120 538.100 293.380 ;
        RECT 793.600 293.120 793.860 293.380 ;
        RECT 793.600 17.380 793.860 17.640 ;
        RECT 799.580 17.380 799.840 17.640 ;
      LAYER met2 ;
        RECT 535.210 510.410 535.490 514.000 ;
        RECT 535.210 510.270 538.040 510.410 ;
        RECT 535.210 510.000 535.490 510.270 ;
        RECT 537.900 293.410 538.040 510.270 ;
        RECT 537.840 293.090 538.100 293.410 ;
        RECT 793.600 293.090 793.860 293.410 ;
        RECT 793.660 17.670 793.800 293.090 ;
        RECT 793.600 17.350 793.860 17.670 ;
        RECT 799.580 17.350 799.840 17.670 ;
        RECT 799.640 2.400 799.780 17.350 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.870 500.040 428.190 500.100 ;
        RECT 534.590 500.040 534.910 500.100 ;
        RECT 427.870 499.900 534.910 500.040 ;
        RECT 427.870 499.840 428.190 499.900 ;
        RECT 534.590 499.840 534.910 499.900 ;
        RECT 534.590 65.860 534.910 65.920 ;
        RECT 641.770 65.860 642.090 65.920 ;
        RECT 534.590 65.720 642.090 65.860 ;
        RECT 534.590 65.660 534.910 65.720 ;
        RECT 641.770 65.660 642.090 65.720 ;
        RECT 641.770 2.960 642.090 3.020 ;
        RECT 644.990 2.960 645.310 3.020 ;
        RECT 641.770 2.820 645.310 2.960 ;
        RECT 641.770 2.760 642.090 2.820 ;
        RECT 644.990 2.760 645.310 2.820 ;
      LAYER via ;
        RECT 427.900 499.840 428.160 500.100 ;
        RECT 534.620 499.840 534.880 500.100 ;
        RECT 534.620 65.660 534.880 65.920 ;
        RECT 641.800 65.660 642.060 65.920 ;
        RECT 641.800 2.760 642.060 3.020 ;
        RECT 645.020 2.760 645.280 3.020 ;
      LAYER met2 ;
        RECT 428.030 510.340 428.310 514.000 ;
        RECT 427.960 510.000 428.310 510.340 ;
        RECT 427.960 500.130 428.100 510.000 ;
        RECT 427.900 499.810 428.160 500.130 ;
        RECT 534.620 499.810 534.880 500.130 ;
        RECT 534.680 65.950 534.820 499.810 ;
        RECT 534.620 65.630 534.880 65.950 ;
        RECT 641.800 65.630 642.060 65.950 ;
        RECT 641.860 3.050 642.000 65.630 ;
        RECT 641.800 2.730 642.060 3.050 ;
        RECT 645.020 2.730 645.280 3.050 ;
        RECT 645.080 2.400 645.220 2.730 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1664.810 496.980 1665.130 497.040 ;
        RECT 1668.950 496.980 1669.270 497.040 ;
        RECT 1664.810 496.840 1669.270 496.980 ;
        RECT 1664.810 496.780 1665.130 496.840 ;
        RECT 1668.950 496.780 1669.270 496.840 ;
        RECT 1668.950 72.660 1669.270 72.720 ;
        RECT 2429.330 72.660 2429.650 72.720 ;
        RECT 1668.950 72.520 2429.650 72.660 ;
        RECT 1668.950 72.460 1669.270 72.520 ;
        RECT 2429.330 72.460 2429.650 72.520 ;
      LAYER via ;
        RECT 1664.840 496.780 1665.100 497.040 ;
        RECT 1668.980 496.780 1669.240 497.040 ;
        RECT 1668.980 72.460 1669.240 72.720 ;
        RECT 2429.360 72.460 2429.620 72.720 ;
      LAYER met2 ;
        RECT 1664.970 510.340 1665.250 514.000 ;
        RECT 1664.900 510.000 1665.250 510.340 ;
        RECT 1664.900 497.070 1665.040 510.000 ;
        RECT 1664.840 496.750 1665.100 497.070 ;
        RECT 1668.980 496.750 1669.240 497.070 ;
        RECT 1669.040 72.750 1669.180 496.750 ;
        RECT 1668.980 72.430 1669.240 72.750 ;
        RECT 2429.360 72.430 2429.620 72.750 ;
        RECT 2429.420 37.130 2429.560 72.430 ;
        RECT 2428.960 36.990 2429.560 37.130 ;
        RECT 2428.960 2.400 2429.100 36.990 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1677.230 500.720 1677.550 500.780 ;
        RECT 1776.590 500.720 1776.910 500.780 ;
        RECT 1677.230 500.580 1776.910 500.720 ;
        RECT 1677.230 500.520 1677.550 500.580 ;
        RECT 1776.590 500.520 1776.910 500.580 ;
        RECT 1776.590 300.460 1776.910 300.520 ;
        RECT 2442.670 300.460 2442.990 300.520 ;
        RECT 1776.590 300.320 2442.990 300.460 ;
        RECT 1776.590 300.260 1776.910 300.320 ;
        RECT 2442.670 300.260 2442.990 300.320 ;
        RECT 2442.670 62.120 2442.990 62.180 ;
        RECT 2446.810 62.120 2447.130 62.180 ;
        RECT 2442.670 61.980 2447.130 62.120 ;
        RECT 2442.670 61.920 2442.990 61.980 ;
        RECT 2446.810 61.920 2447.130 61.980 ;
      LAYER via ;
        RECT 1677.260 500.520 1677.520 500.780 ;
        RECT 1776.620 500.520 1776.880 500.780 ;
        RECT 1776.620 300.260 1776.880 300.520 ;
        RECT 2442.700 300.260 2442.960 300.520 ;
        RECT 2442.700 61.920 2442.960 62.180 ;
        RECT 2446.840 61.920 2447.100 62.180 ;
      LAYER met2 ;
        RECT 1677.390 510.340 1677.670 514.000 ;
        RECT 1677.320 510.000 1677.670 510.340 ;
        RECT 1677.320 500.810 1677.460 510.000 ;
        RECT 1677.260 500.490 1677.520 500.810 ;
        RECT 1776.620 500.490 1776.880 500.810 ;
        RECT 1776.680 300.550 1776.820 500.490 ;
        RECT 1776.620 300.230 1776.880 300.550 ;
        RECT 2442.700 300.230 2442.960 300.550 ;
        RECT 2442.760 62.210 2442.900 300.230 ;
        RECT 2442.700 61.890 2442.960 62.210 ;
        RECT 2446.840 61.890 2447.100 62.210 ;
        RECT 2446.900 2.400 2447.040 61.890 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2463.445 48.365 2463.615 96.475 ;
      LAYER mcon ;
        RECT 2463.445 96.305 2463.615 96.475 ;
      LAYER met1 ;
        RECT 1690.110 113.800 1690.430 113.860 ;
        RECT 2463.370 113.800 2463.690 113.860 ;
        RECT 1690.110 113.660 2463.690 113.800 ;
        RECT 1690.110 113.600 1690.430 113.660 ;
        RECT 2463.370 113.600 2463.690 113.660 ;
        RECT 2463.370 96.460 2463.690 96.520 ;
        RECT 2463.370 96.320 2463.885 96.460 ;
        RECT 2463.370 96.260 2463.690 96.320 ;
        RECT 2463.385 48.520 2463.675 48.565 ;
        RECT 2464.750 48.520 2465.070 48.580 ;
        RECT 2463.385 48.380 2465.070 48.520 ;
        RECT 2463.385 48.335 2463.675 48.380 ;
        RECT 2464.750 48.320 2465.070 48.380 ;
      LAYER via ;
        RECT 1690.140 113.600 1690.400 113.860 ;
        RECT 2463.400 113.600 2463.660 113.860 ;
        RECT 2463.400 96.260 2463.660 96.520 ;
        RECT 2464.780 48.320 2465.040 48.580 ;
      LAYER met2 ;
        RECT 1689.810 510.340 1690.090 514.000 ;
        RECT 1689.740 510.000 1690.090 510.340 ;
        RECT 1689.740 497.490 1689.880 510.000 ;
        RECT 1689.740 497.350 1690.340 497.490 ;
        RECT 1690.200 113.890 1690.340 497.350 ;
        RECT 1690.140 113.570 1690.400 113.890 ;
        RECT 2463.400 113.570 2463.660 113.890 ;
        RECT 2463.460 96.550 2463.600 113.570 ;
        RECT 2463.400 96.230 2463.660 96.550 ;
        RECT 2464.780 48.290 2465.040 48.610 ;
        RECT 2464.840 2.400 2464.980 48.290 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 293.320 1703.770 293.380 ;
        RECT 2477.170 293.320 2477.490 293.380 ;
        RECT 1703.450 293.180 2477.490 293.320 ;
        RECT 1703.450 293.120 1703.770 293.180 ;
        RECT 2477.170 293.120 2477.490 293.180 ;
      LAYER via ;
        RECT 1703.480 293.120 1703.740 293.380 ;
        RECT 2477.200 293.120 2477.460 293.380 ;
      LAYER met2 ;
        RECT 1702.230 510.410 1702.510 514.000 ;
        RECT 1702.230 510.270 1703.680 510.410 ;
        RECT 1702.230 510.000 1702.510 510.270 ;
        RECT 1703.540 293.410 1703.680 510.270 ;
        RECT 1703.480 293.090 1703.740 293.410 ;
        RECT 2477.200 293.090 2477.460 293.410 ;
        RECT 2477.260 17.410 2477.400 293.090 ;
        RECT 2477.260 17.270 2482.920 17.410 ;
        RECT 2482.780 2.400 2482.920 17.270 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 120.600 1718.030 120.660 ;
        RECT 2497.870 120.600 2498.190 120.660 ;
        RECT 1717.710 120.460 2498.190 120.600 ;
        RECT 1717.710 120.400 1718.030 120.460 ;
        RECT 2497.870 120.400 2498.190 120.460 ;
      LAYER via ;
        RECT 1717.740 120.400 1718.000 120.660 ;
        RECT 2497.900 120.400 2498.160 120.660 ;
      LAYER met2 ;
        RECT 1714.650 510.410 1714.930 514.000 ;
        RECT 1714.650 510.270 1717.940 510.410 ;
        RECT 1714.650 510.000 1714.930 510.270 ;
        RECT 1717.800 120.690 1717.940 510.270 ;
        RECT 1717.740 120.370 1718.000 120.690 ;
        RECT 2497.900 120.370 2498.160 120.690 ;
        RECT 2497.960 17.410 2498.100 120.370 ;
        RECT 2497.960 17.270 2500.860 17.410 ;
        RECT 2500.720 2.400 2500.860 17.270 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1726.910 503.440 1727.230 503.500 ;
        RECT 1731.510 503.440 1731.830 503.500 ;
        RECT 1726.910 503.300 1731.830 503.440 ;
        RECT 1726.910 503.240 1727.230 503.300 ;
        RECT 1731.510 503.240 1731.830 503.300 ;
        RECT 1731.510 196.760 1731.830 196.820 ;
        RECT 2512.130 196.760 2512.450 196.820 ;
        RECT 1731.510 196.620 2512.450 196.760 ;
        RECT 1731.510 196.560 1731.830 196.620 ;
        RECT 2512.130 196.560 2512.450 196.620 ;
        RECT 2512.130 17.920 2512.450 17.980 ;
        RECT 2518.110 17.920 2518.430 17.980 ;
        RECT 2512.130 17.780 2518.430 17.920 ;
        RECT 2512.130 17.720 2512.450 17.780 ;
        RECT 2518.110 17.720 2518.430 17.780 ;
      LAYER via ;
        RECT 1726.940 503.240 1727.200 503.500 ;
        RECT 1731.540 503.240 1731.800 503.500 ;
        RECT 1731.540 196.560 1731.800 196.820 ;
        RECT 2512.160 196.560 2512.420 196.820 ;
        RECT 2512.160 17.720 2512.420 17.980 ;
        RECT 2518.140 17.720 2518.400 17.980 ;
      LAYER met2 ;
        RECT 1727.070 510.340 1727.350 514.000 ;
        RECT 1727.000 510.000 1727.350 510.340 ;
        RECT 1727.000 503.530 1727.140 510.000 ;
        RECT 1726.940 503.210 1727.200 503.530 ;
        RECT 1731.540 503.210 1731.800 503.530 ;
        RECT 1731.600 196.850 1731.740 503.210 ;
        RECT 1731.540 196.530 1731.800 196.850 ;
        RECT 2512.160 196.530 2512.420 196.850 ;
        RECT 2512.220 18.010 2512.360 196.530 ;
        RECT 2512.160 17.690 2512.420 18.010 ;
        RECT 2518.140 17.690 2518.400 18.010 ;
        RECT 2518.200 2.400 2518.340 17.690 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 503.440 1739.650 503.500 ;
        RECT 1744.850 503.440 1745.170 503.500 ;
        RECT 1739.330 503.300 1745.170 503.440 ;
        RECT 1739.330 503.240 1739.650 503.300 ;
        RECT 1744.850 503.240 1745.170 503.300 ;
        RECT 1744.850 189.620 1745.170 189.680 ;
        RECT 2532.370 189.620 2532.690 189.680 ;
        RECT 1744.850 189.480 2532.690 189.620 ;
        RECT 1744.850 189.420 1745.170 189.480 ;
        RECT 2532.370 189.420 2532.690 189.480 ;
        RECT 2532.370 62.120 2532.690 62.180 ;
        RECT 2536.050 62.120 2536.370 62.180 ;
        RECT 2532.370 61.980 2536.370 62.120 ;
        RECT 2532.370 61.920 2532.690 61.980 ;
        RECT 2536.050 61.920 2536.370 61.980 ;
      LAYER via ;
        RECT 1739.360 503.240 1739.620 503.500 ;
        RECT 1744.880 503.240 1745.140 503.500 ;
        RECT 1744.880 189.420 1745.140 189.680 ;
        RECT 2532.400 189.420 2532.660 189.680 ;
        RECT 2532.400 61.920 2532.660 62.180 ;
        RECT 2536.080 61.920 2536.340 62.180 ;
      LAYER met2 ;
        RECT 1739.490 510.340 1739.770 514.000 ;
        RECT 1739.420 510.000 1739.770 510.340 ;
        RECT 1739.420 503.530 1739.560 510.000 ;
        RECT 1739.360 503.210 1739.620 503.530 ;
        RECT 1744.880 503.210 1745.140 503.530 ;
        RECT 1744.940 189.710 1745.080 503.210 ;
        RECT 1744.880 189.390 1745.140 189.710 ;
        RECT 2532.400 189.390 2532.660 189.710 ;
        RECT 2532.460 62.210 2532.600 189.390 ;
        RECT 2532.400 61.890 2532.660 62.210 ;
        RECT 2536.080 61.890 2536.340 62.210 ;
        RECT 2536.140 2.400 2536.280 61.890 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2553.145 48.365 2553.315 96.475 ;
      LAYER mcon ;
        RECT 2553.145 96.305 2553.315 96.475 ;
      LAYER met1 ;
        RECT 1752.210 127.740 1752.530 127.800 ;
        RECT 2553.530 127.740 2553.850 127.800 ;
        RECT 1752.210 127.600 2553.850 127.740 ;
        RECT 1752.210 127.540 1752.530 127.600 ;
        RECT 2553.530 127.540 2553.850 127.600 ;
        RECT 2553.070 96.460 2553.390 96.520 ;
        RECT 2552.875 96.320 2553.390 96.460 ;
        RECT 2553.070 96.260 2553.390 96.320 ;
        RECT 2553.085 48.520 2553.375 48.565 ;
        RECT 2553.990 48.520 2554.310 48.580 ;
        RECT 2553.085 48.380 2554.310 48.520 ;
        RECT 2553.085 48.335 2553.375 48.380 ;
        RECT 2553.990 48.320 2554.310 48.380 ;
      LAYER via ;
        RECT 1752.240 127.540 1752.500 127.800 ;
        RECT 2553.560 127.540 2553.820 127.800 ;
        RECT 2553.100 96.260 2553.360 96.520 ;
        RECT 2554.020 48.320 2554.280 48.580 ;
      LAYER met2 ;
        RECT 1751.910 510.340 1752.190 514.000 ;
        RECT 1751.840 510.000 1752.190 510.340 ;
        RECT 1751.840 504.290 1751.980 510.000 ;
        RECT 1751.840 504.150 1752.440 504.290 ;
        RECT 1752.300 127.830 1752.440 504.150 ;
        RECT 1752.240 127.510 1752.500 127.830 ;
        RECT 2553.560 127.510 2553.820 127.830 ;
        RECT 2553.620 96.970 2553.760 127.510 ;
        RECT 2553.160 96.830 2553.760 96.970 ;
        RECT 2553.160 96.550 2553.300 96.830 ;
        RECT 2553.100 96.230 2553.360 96.550 ;
        RECT 2554.020 48.290 2554.280 48.610 ;
        RECT 2554.080 2.400 2554.220 48.290 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 134.540 1766.330 134.600 ;
        RECT 2566.870 134.540 2567.190 134.600 ;
        RECT 1766.010 134.400 2567.190 134.540 ;
        RECT 1766.010 134.340 1766.330 134.400 ;
        RECT 2566.870 134.340 2567.190 134.400 ;
        RECT 2566.870 62.120 2567.190 62.180 ;
        RECT 2571.930 62.120 2572.250 62.180 ;
        RECT 2566.870 61.980 2572.250 62.120 ;
        RECT 2566.870 61.920 2567.190 61.980 ;
        RECT 2571.930 61.920 2572.250 61.980 ;
      LAYER via ;
        RECT 1766.040 134.340 1766.300 134.600 ;
        RECT 2566.900 134.340 2567.160 134.600 ;
        RECT 2566.900 61.920 2567.160 62.180 ;
        RECT 2571.960 61.920 2572.220 62.180 ;
      LAYER met2 ;
        RECT 1764.330 510.410 1764.610 514.000 ;
        RECT 1764.330 510.270 1766.240 510.410 ;
        RECT 1764.330 510.000 1764.610 510.270 ;
        RECT 1766.100 134.630 1766.240 510.270 ;
        RECT 1766.040 134.310 1766.300 134.630 ;
        RECT 2566.900 134.310 2567.160 134.630 ;
        RECT 2566.960 62.210 2567.100 134.310 ;
        RECT 2566.900 61.890 2567.160 62.210 ;
        RECT 2571.960 61.890 2572.220 62.210 ;
        RECT 2572.020 2.400 2572.160 61.890 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2589.485 2.805 2589.655 48.195 ;
      LAYER mcon ;
        RECT 2589.485 48.025 2589.655 48.195 ;
      LAYER met1 ;
        RECT 1779.810 210.360 1780.130 210.420 ;
        RECT 2587.570 210.360 2587.890 210.420 ;
        RECT 1779.810 210.220 2587.890 210.360 ;
        RECT 1779.810 210.160 1780.130 210.220 ;
        RECT 2587.570 210.160 2587.890 210.220 ;
        RECT 2587.570 62.260 2587.890 62.520 ;
        RECT 2587.660 61.780 2587.800 62.260 ;
        RECT 2589.410 61.780 2589.730 61.840 ;
        RECT 2587.660 61.640 2589.730 61.780 ;
        RECT 2589.410 61.580 2589.730 61.640 ;
        RECT 2589.410 48.180 2589.730 48.240 ;
        RECT 2589.215 48.040 2589.730 48.180 ;
        RECT 2589.410 47.980 2589.730 48.040 ;
        RECT 2589.410 2.960 2589.730 3.020 ;
        RECT 2589.215 2.820 2589.730 2.960 ;
        RECT 2589.410 2.760 2589.730 2.820 ;
      LAYER via ;
        RECT 1779.840 210.160 1780.100 210.420 ;
        RECT 2587.600 210.160 2587.860 210.420 ;
        RECT 2587.600 62.260 2587.860 62.520 ;
        RECT 2589.440 61.580 2589.700 61.840 ;
        RECT 2589.440 47.980 2589.700 48.240 ;
        RECT 2589.440 2.760 2589.700 3.020 ;
      LAYER met2 ;
        RECT 1776.290 510.410 1776.570 514.000 ;
        RECT 1776.290 510.270 1780.040 510.410 ;
        RECT 1776.290 510.000 1776.570 510.270 ;
        RECT 1779.900 210.450 1780.040 510.270 ;
        RECT 1779.840 210.130 1780.100 210.450 ;
        RECT 2587.600 210.130 2587.860 210.450 ;
        RECT 2587.660 62.550 2587.800 210.130 ;
        RECT 2587.600 62.230 2587.860 62.550 ;
        RECT 2589.440 61.550 2589.700 61.870 ;
        RECT 2589.500 48.270 2589.640 61.550 ;
        RECT 2589.440 47.950 2589.700 48.270 ;
        RECT 2589.440 2.730 2589.700 3.050 ;
        RECT 2589.500 2.400 2589.640 2.730 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 306.920 551.930 306.980 ;
        RECT 821.170 306.920 821.490 306.980 ;
        RECT 551.610 306.780 821.490 306.920 ;
        RECT 551.610 306.720 551.930 306.780 ;
        RECT 821.170 306.720 821.490 306.780 ;
      LAYER via ;
        RECT 551.640 306.720 551.900 306.980 ;
        RECT 821.200 306.720 821.460 306.980 ;
      LAYER met2 ;
        RECT 551.770 510.340 552.050 514.000 ;
        RECT 551.700 510.000 552.050 510.340 ;
        RECT 551.700 307.010 551.840 510.000 ;
        RECT 551.640 306.690 551.900 307.010 ;
        RECT 821.200 306.690 821.460 307.010 ;
        RECT 821.260 17.410 821.400 306.690 ;
        RECT 821.260 17.270 823.700 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1788.550 496.980 1788.870 497.040 ;
        RECT 1793.610 496.980 1793.930 497.040 ;
        RECT 1788.550 496.840 1793.930 496.980 ;
        RECT 1788.550 496.780 1788.870 496.840 ;
        RECT 1793.610 496.780 1793.930 496.840 ;
        RECT 1793.610 30.840 1793.930 30.900 ;
        RECT 2607.350 30.840 2607.670 30.900 ;
        RECT 1793.610 30.700 2607.670 30.840 ;
        RECT 1793.610 30.640 1793.930 30.700 ;
        RECT 2607.350 30.640 2607.670 30.700 ;
      LAYER via ;
        RECT 1788.580 496.780 1788.840 497.040 ;
        RECT 1793.640 496.780 1793.900 497.040 ;
        RECT 1793.640 30.640 1793.900 30.900 ;
        RECT 2607.380 30.640 2607.640 30.900 ;
      LAYER met2 ;
        RECT 1788.710 510.340 1788.990 514.000 ;
        RECT 1788.640 510.000 1788.990 510.340 ;
        RECT 1788.640 497.070 1788.780 510.000 ;
        RECT 1788.580 496.750 1788.840 497.070 ;
        RECT 1793.640 496.750 1793.900 497.070 ;
        RECT 1793.700 30.930 1793.840 496.750 ;
        RECT 1793.640 30.610 1793.900 30.930 ;
        RECT 2607.380 30.610 2607.640 30.930 ;
        RECT 2607.440 2.400 2607.580 30.610 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.970 496.980 1801.290 497.040 ;
        RECT 1807.410 496.980 1807.730 497.040 ;
        RECT 1800.970 496.840 1807.730 496.980 ;
        RECT 1800.970 496.780 1801.290 496.840 ;
        RECT 1807.410 496.780 1807.730 496.840 ;
        RECT 1807.410 141.340 1807.730 141.400 ;
        RECT 2622.530 141.340 2622.850 141.400 ;
        RECT 1807.410 141.200 2622.850 141.340 ;
        RECT 1807.410 141.140 1807.730 141.200 ;
        RECT 2622.530 141.140 2622.850 141.200 ;
        RECT 2622.070 62.260 2622.390 62.520 ;
        RECT 2622.160 61.780 2622.300 62.260 ;
        RECT 2625.290 61.780 2625.610 61.840 ;
        RECT 2622.160 61.640 2625.610 61.780 ;
        RECT 2625.290 61.580 2625.610 61.640 ;
        RECT 2625.290 47.980 2625.610 48.240 ;
        RECT 2625.380 47.560 2625.520 47.980 ;
        RECT 2625.290 47.300 2625.610 47.560 ;
      LAYER via ;
        RECT 1801.000 496.780 1801.260 497.040 ;
        RECT 1807.440 496.780 1807.700 497.040 ;
        RECT 1807.440 141.140 1807.700 141.400 ;
        RECT 2622.560 141.140 2622.820 141.400 ;
        RECT 2622.100 62.260 2622.360 62.520 ;
        RECT 2625.320 61.580 2625.580 61.840 ;
        RECT 2625.320 47.980 2625.580 48.240 ;
        RECT 2625.320 47.300 2625.580 47.560 ;
      LAYER met2 ;
        RECT 1801.130 510.340 1801.410 514.000 ;
        RECT 1801.060 510.000 1801.410 510.340 ;
        RECT 1801.060 497.070 1801.200 510.000 ;
        RECT 1801.000 496.750 1801.260 497.070 ;
        RECT 1807.440 496.750 1807.700 497.070 ;
        RECT 1807.500 141.430 1807.640 496.750 ;
        RECT 1807.440 141.110 1807.700 141.430 ;
        RECT 2622.560 141.110 2622.820 141.430 ;
        RECT 2622.620 96.970 2622.760 141.110 ;
        RECT 2622.160 96.830 2622.760 96.970 ;
        RECT 2622.160 62.550 2622.300 96.830 ;
        RECT 2622.100 62.230 2622.360 62.550 ;
        RECT 2625.320 61.550 2625.580 61.870 ;
        RECT 2625.380 48.270 2625.520 61.550 ;
        RECT 2625.320 47.950 2625.580 48.270 ;
        RECT 2625.320 47.270 2625.580 47.590 ;
        RECT 2625.380 2.400 2625.520 47.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 37.980 1814.630 38.040 ;
        RECT 1814.310 37.840 2628.740 37.980 ;
        RECT 1814.310 37.780 1814.630 37.840 ;
        RECT 2628.600 37.640 2628.740 37.840 ;
        RECT 2643.230 37.640 2643.550 37.700 ;
        RECT 2628.600 37.500 2643.550 37.640 ;
        RECT 2643.230 37.440 2643.550 37.500 ;
      LAYER via ;
        RECT 1814.340 37.780 1814.600 38.040 ;
        RECT 2643.260 37.440 2643.520 37.700 ;
      LAYER met2 ;
        RECT 1813.550 510.410 1813.830 514.000 ;
        RECT 1813.550 510.270 1814.540 510.410 ;
        RECT 1813.550 510.000 1813.830 510.270 ;
        RECT 1814.400 38.070 1814.540 510.270 ;
        RECT 1814.340 37.750 1814.600 38.070 ;
        RECT 2643.260 37.410 2643.520 37.730 ;
        RECT 2643.320 2.400 2643.460 37.410 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 217.160 1828.430 217.220 ;
        RECT 2656.570 217.160 2656.890 217.220 ;
        RECT 1828.110 217.020 2656.890 217.160 ;
        RECT 1828.110 216.960 1828.430 217.020 ;
        RECT 2656.570 216.960 2656.890 217.020 ;
        RECT 2656.570 62.120 2656.890 62.180 ;
        RECT 2661.170 62.120 2661.490 62.180 ;
        RECT 2656.570 61.980 2661.490 62.120 ;
        RECT 2656.570 61.920 2656.890 61.980 ;
        RECT 2661.170 61.920 2661.490 61.980 ;
      LAYER via ;
        RECT 1828.140 216.960 1828.400 217.220 ;
        RECT 2656.600 216.960 2656.860 217.220 ;
        RECT 2656.600 61.920 2656.860 62.180 ;
        RECT 2661.200 61.920 2661.460 62.180 ;
      LAYER met2 ;
        RECT 1825.970 510.410 1826.250 514.000 ;
        RECT 1825.970 510.270 1828.340 510.410 ;
        RECT 1825.970 510.000 1826.250 510.270 ;
        RECT 1828.200 217.250 1828.340 510.270 ;
        RECT 1828.140 216.930 1828.400 217.250 ;
        RECT 2656.600 216.930 2656.860 217.250 ;
        RECT 2656.660 62.210 2656.800 216.930 ;
        RECT 2656.600 61.890 2656.860 62.210 ;
        RECT 2661.200 61.890 2661.460 62.210 ;
        RECT 2661.260 2.400 2661.400 61.890 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1838.230 496.980 1838.550 497.040 ;
        RECT 1841.910 496.980 1842.230 497.040 ;
        RECT 1838.230 496.840 1842.230 496.980 ;
        RECT 1838.230 496.780 1838.550 496.840 ;
        RECT 1841.910 496.780 1842.230 496.840 ;
        RECT 1841.910 224.300 1842.230 224.360 ;
        RECT 2677.270 224.300 2677.590 224.360 ;
        RECT 1841.910 224.160 2677.590 224.300 ;
        RECT 1841.910 224.100 1842.230 224.160 ;
        RECT 2677.270 224.100 2677.590 224.160 ;
      LAYER via ;
        RECT 1838.260 496.780 1838.520 497.040 ;
        RECT 1841.940 496.780 1842.200 497.040 ;
        RECT 1841.940 224.100 1842.200 224.360 ;
        RECT 2677.300 224.100 2677.560 224.360 ;
      LAYER met2 ;
        RECT 1838.390 510.340 1838.670 514.000 ;
        RECT 1838.320 510.000 1838.670 510.340 ;
        RECT 1838.320 497.070 1838.460 510.000 ;
        RECT 1838.260 496.750 1838.520 497.070 ;
        RECT 1841.940 496.750 1842.200 497.070 ;
        RECT 1842.000 224.390 1842.140 496.750 ;
        RECT 1841.940 224.070 1842.200 224.390 ;
        RECT 2677.300 224.070 2677.560 224.390 ;
        RECT 2677.360 17.410 2677.500 224.070 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1850.650 503.440 1850.970 503.500 ;
        RECT 1855.710 503.440 1856.030 503.500 ;
        RECT 1850.650 503.300 1856.030 503.440 ;
        RECT 1850.650 503.240 1850.970 503.300 ;
        RECT 1855.710 503.240 1856.030 503.300 ;
        RECT 1855.710 231.100 1856.030 231.160 ;
        RECT 2691.070 231.100 2691.390 231.160 ;
        RECT 1855.710 230.960 2691.390 231.100 ;
        RECT 1855.710 230.900 1856.030 230.960 ;
        RECT 2691.070 230.900 2691.390 230.960 ;
      LAYER via ;
        RECT 1850.680 503.240 1850.940 503.500 ;
        RECT 1855.740 503.240 1856.000 503.500 ;
        RECT 1855.740 230.900 1856.000 231.160 ;
        RECT 2691.100 230.900 2691.360 231.160 ;
      LAYER met2 ;
        RECT 1850.810 510.340 1851.090 514.000 ;
        RECT 1850.740 510.000 1851.090 510.340 ;
        RECT 1850.740 503.530 1850.880 510.000 ;
        RECT 1850.680 503.210 1850.940 503.530 ;
        RECT 1855.740 503.210 1856.000 503.530 ;
        RECT 1855.800 231.190 1855.940 503.210 ;
        RECT 1855.740 230.870 1856.000 231.190 ;
        RECT 2691.100 230.870 2691.360 231.190 ;
        RECT 2691.160 16.730 2691.300 230.870 ;
        RECT 2691.160 16.590 2696.820 16.730 ;
        RECT 2696.680 2.400 2696.820 16.590 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1863.070 500.720 1863.390 500.780 ;
        RECT 1869.050 500.720 1869.370 500.780 ;
        RECT 1863.070 500.580 1869.370 500.720 ;
        RECT 1863.070 500.520 1863.390 500.580 ;
        RECT 1869.050 500.520 1869.370 500.580 ;
        RECT 1869.050 237.900 1869.370 237.960 ;
        RECT 2711.770 237.900 2712.090 237.960 ;
        RECT 1869.050 237.760 2712.090 237.900 ;
        RECT 1869.050 237.700 1869.370 237.760 ;
        RECT 2711.770 237.700 2712.090 237.760 ;
      LAYER via ;
        RECT 1863.100 500.520 1863.360 500.780 ;
        RECT 1869.080 500.520 1869.340 500.780 ;
        RECT 1869.080 237.700 1869.340 237.960 ;
        RECT 2711.800 237.700 2712.060 237.960 ;
      LAYER met2 ;
        RECT 1863.230 510.340 1863.510 514.000 ;
        RECT 1863.160 510.000 1863.510 510.340 ;
        RECT 1863.160 500.810 1863.300 510.000 ;
        RECT 1863.100 500.490 1863.360 500.810 ;
        RECT 1869.080 500.490 1869.340 500.810 ;
        RECT 1869.140 237.990 1869.280 500.490 ;
        RECT 1869.080 237.670 1869.340 237.990 ;
        RECT 2711.800 237.670 2712.060 237.990 ;
        RECT 2711.860 16.730 2712.000 237.670 ;
        RECT 2711.860 16.590 2714.760 16.730 ;
        RECT 2714.620 2.400 2714.760 16.590 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 44.780 1876.730 44.840 ;
        RECT 2732.930 44.780 2733.250 44.840 ;
        RECT 1876.410 44.640 2733.250 44.780 ;
        RECT 1876.410 44.580 1876.730 44.640 ;
        RECT 2732.930 44.580 2733.250 44.640 ;
      LAYER via ;
        RECT 1876.440 44.580 1876.700 44.840 ;
        RECT 2732.960 44.580 2733.220 44.840 ;
      LAYER met2 ;
        RECT 1875.650 510.410 1875.930 514.000 ;
        RECT 1875.650 510.270 1876.640 510.410 ;
        RECT 1875.650 510.000 1875.930 510.270 ;
        RECT 1876.500 44.870 1876.640 510.270 ;
        RECT 1876.440 44.550 1876.700 44.870 ;
        RECT 2732.960 44.550 2733.220 44.870 ;
        RECT 2733.020 37.130 2733.160 44.550 ;
        RECT 2732.560 36.990 2733.160 37.130 ;
        RECT 2732.560 2.400 2732.700 36.990 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2750.485 2.805 2750.655 48.195 ;
      LAYER mcon ;
        RECT 2750.485 48.025 2750.655 48.195 ;
      LAYER met1 ;
        RECT 1890.210 245.040 1890.530 245.100 ;
        RECT 2746.270 245.040 2746.590 245.100 ;
        RECT 1890.210 244.900 2746.590 245.040 ;
        RECT 1890.210 244.840 1890.530 244.900 ;
        RECT 2746.270 244.840 2746.590 244.900 ;
        RECT 2746.270 62.120 2746.590 62.180 ;
        RECT 2750.410 62.120 2750.730 62.180 ;
        RECT 2746.270 61.980 2750.730 62.120 ;
        RECT 2746.270 61.920 2746.590 61.980 ;
        RECT 2750.410 61.920 2750.730 61.980 ;
        RECT 2750.410 48.180 2750.730 48.240 ;
        RECT 2750.215 48.040 2750.730 48.180 ;
        RECT 2750.410 47.980 2750.730 48.040 ;
        RECT 2750.410 2.960 2750.730 3.020 ;
        RECT 2750.215 2.820 2750.730 2.960 ;
        RECT 2750.410 2.760 2750.730 2.820 ;
      LAYER via ;
        RECT 1890.240 244.840 1890.500 245.100 ;
        RECT 2746.300 244.840 2746.560 245.100 ;
        RECT 2746.300 61.920 2746.560 62.180 ;
        RECT 2750.440 61.920 2750.700 62.180 ;
        RECT 2750.440 47.980 2750.700 48.240 ;
        RECT 2750.440 2.760 2750.700 3.020 ;
      LAYER met2 ;
        RECT 1888.070 510.410 1888.350 514.000 ;
        RECT 1888.070 510.270 1890.440 510.410 ;
        RECT 1888.070 510.000 1888.350 510.270 ;
        RECT 1890.300 245.130 1890.440 510.270 ;
        RECT 1890.240 244.810 1890.500 245.130 ;
        RECT 2746.300 244.810 2746.560 245.130 ;
        RECT 2746.360 62.210 2746.500 244.810 ;
        RECT 2746.300 61.890 2746.560 62.210 ;
        RECT 2750.440 61.890 2750.700 62.210 ;
        RECT 2750.500 48.270 2750.640 61.890 ;
        RECT 2750.440 47.950 2750.700 48.270 ;
        RECT 2750.440 2.730 2750.700 3.050 ;
        RECT 2750.500 2.400 2750.640 2.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2767.045 48.365 2767.215 96.475 ;
      LAYER mcon ;
        RECT 2767.045 96.305 2767.215 96.475 ;
      LAYER met1 ;
        RECT 1899.870 496.980 1900.190 497.040 ;
        RECT 1903.550 496.980 1903.870 497.040 ;
        RECT 1899.870 496.840 1903.870 496.980 ;
        RECT 1899.870 496.780 1900.190 496.840 ;
        RECT 1903.550 496.780 1903.870 496.840 ;
        RECT 1903.550 155.280 1903.870 155.340 ;
        RECT 2766.970 155.280 2767.290 155.340 ;
        RECT 1903.550 155.140 2767.290 155.280 ;
        RECT 1903.550 155.080 1903.870 155.140 ;
        RECT 2766.970 155.080 2767.290 155.140 ;
        RECT 2766.970 96.460 2767.290 96.520 ;
        RECT 2766.775 96.320 2767.290 96.460 ;
        RECT 2766.970 96.260 2767.290 96.320 ;
        RECT 2766.985 48.520 2767.275 48.565 ;
        RECT 2767.890 48.520 2768.210 48.580 ;
        RECT 2766.985 48.380 2768.210 48.520 ;
        RECT 2766.985 48.335 2767.275 48.380 ;
        RECT 2767.890 48.320 2768.210 48.380 ;
      LAYER via ;
        RECT 1899.900 496.780 1900.160 497.040 ;
        RECT 1903.580 496.780 1903.840 497.040 ;
        RECT 1903.580 155.080 1903.840 155.340 ;
        RECT 2767.000 155.080 2767.260 155.340 ;
        RECT 2767.000 96.260 2767.260 96.520 ;
        RECT 2767.920 48.320 2768.180 48.580 ;
      LAYER met2 ;
        RECT 1900.030 510.340 1900.310 514.000 ;
        RECT 1899.960 510.000 1900.310 510.340 ;
        RECT 1899.960 497.070 1900.100 510.000 ;
        RECT 1899.900 496.750 1900.160 497.070 ;
        RECT 1903.580 496.750 1903.840 497.070 ;
        RECT 1903.640 155.370 1903.780 496.750 ;
        RECT 1903.580 155.050 1903.840 155.370 ;
        RECT 2767.000 155.050 2767.260 155.370 ;
        RECT 2767.060 96.550 2767.200 155.050 ;
        RECT 2767.000 96.230 2767.260 96.550 ;
        RECT 2767.920 48.290 2768.180 48.610 ;
        RECT 2767.980 2.400 2768.120 48.290 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 314.060 565.730 314.120 ;
        RECT 834.970 314.060 835.290 314.120 ;
        RECT 565.410 313.920 835.290 314.060 ;
        RECT 565.410 313.860 565.730 313.920 ;
        RECT 834.970 313.860 835.290 313.920 ;
        RECT 834.970 17.580 835.290 17.640 ;
        RECT 840.950 17.580 841.270 17.640 ;
        RECT 834.970 17.440 841.270 17.580 ;
        RECT 834.970 17.380 835.290 17.440 ;
        RECT 840.950 17.380 841.270 17.440 ;
      LAYER via ;
        RECT 565.440 313.860 565.700 314.120 ;
        RECT 835.000 313.860 835.260 314.120 ;
        RECT 835.000 17.380 835.260 17.640 ;
        RECT 840.980 17.380 841.240 17.640 ;
      LAYER met2 ;
        RECT 564.190 510.410 564.470 514.000 ;
        RECT 564.190 510.270 565.640 510.410 ;
        RECT 564.190 510.000 564.470 510.270 ;
        RECT 565.500 314.150 565.640 510.270 ;
        RECT 565.440 313.830 565.700 314.150 ;
        RECT 835.000 313.830 835.260 314.150 ;
        RECT 835.060 17.670 835.200 313.830 ;
        RECT 835.000 17.350 835.260 17.670 ;
        RECT 840.980 17.350 841.240 17.670 ;
        RECT 841.040 2.400 841.180 17.350 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1912.290 496.980 1912.610 497.040 ;
        RECT 1917.810 496.980 1918.130 497.040 ;
        RECT 1912.290 496.840 1918.130 496.980 ;
        RECT 1912.290 496.780 1912.610 496.840 ;
        RECT 1917.810 496.780 1918.130 496.840 ;
        RECT 1917.810 51.580 1918.130 51.640 ;
        RECT 2785.830 51.580 2786.150 51.640 ;
        RECT 1917.810 51.440 2786.150 51.580 ;
        RECT 1917.810 51.380 1918.130 51.440 ;
        RECT 2785.830 51.380 2786.150 51.440 ;
      LAYER via ;
        RECT 1912.320 496.780 1912.580 497.040 ;
        RECT 1917.840 496.780 1918.100 497.040 ;
        RECT 1917.840 51.380 1918.100 51.640 ;
        RECT 2785.860 51.380 2786.120 51.640 ;
      LAYER met2 ;
        RECT 1912.450 510.340 1912.730 514.000 ;
        RECT 1912.380 510.000 1912.730 510.340 ;
        RECT 1912.380 497.070 1912.520 510.000 ;
        RECT 1912.320 496.750 1912.580 497.070 ;
        RECT 1917.840 496.750 1918.100 497.070 ;
        RECT 1917.900 51.670 1918.040 496.750 ;
        RECT 1917.840 51.350 1918.100 51.670 ;
        RECT 2785.860 51.350 2786.120 51.670 ;
        RECT 2785.920 2.400 2786.060 51.350 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.710 162.080 1925.030 162.140 ;
        RECT 2801.470 162.080 2801.790 162.140 ;
        RECT 1924.710 161.940 2801.790 162.080 ;
        RECT 1924.710 161.880 1925.030 161.940 ;
        RECT 2801.470 161.880 2801.790 161.940 ;
        RECT 2801.470 96.460 2801.790 96.520 ;
        RECT 2803.770 96.460 2804.090 96.520 ;
        RECT 2801.470 96.320 2804.090 96.460 ;
        RECT 2801.470 96.260 2801.790 96.320 ;
        RECT 2803.770 96.260 2804.090 96.320 ;
      LAYER via ;
        RECT 1924.740 161.880 1925.000 162.140 ;
        RECT 2801.500 161.880 2801.760 162.140 ;
        RECT 2801.500 96.260 2801.760 96.520 ;
        RECT 2803.800 96.260 2804.060 96.520 ;
      LAYER met2 ;
        RECT 1924.870 510.340 1925.150 514.000 ;
        RECT 1924.800 510.000 1925.150 510.340 ;
        RECT 1924.800 162.170 1924.940 510.000 ;
        RECT 1924.740 161.850 1925.000 162.170 ;
        RECT 2801.500 161.850 2801.760 162.170 ;
        RECT 2801.560 96.550 2801.700 161.850 ;
        RECT 2801.500 96.230 2801.760 96.550 ;
        RECT 2803.800 96.230 2804.060 96.550 ;
        RECT 2803.860 2.400 2804.000 96.230 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 168.880 1938.830 168.940 ;
        RECT 2815.730 168.880 2816.050 168.940 ;
        RECT 1938.510 168.740 2816.050 168.880 ;
        RECT 1938.510 168.680 1938.830 168.740 ;
        RECT 2815.730 168.680 2816.050 168.740 ;
        RECT 2815.730 37.980 2816.050 38.040 ;
        RECT 2821.710 37.980 2822.030 38.040 ;
        RECT 2815.730 37.840 2822.030 37.980 ;
        RECT 2815.730 37.780 2816.050 37.840 ;
        RECT 2821.710 37.780 2822.030 37.840 ;
      LAYER via ;
        RECT 1938.540 168.680 1938.800 168.940 ;
        RECT 2815.760 168.680 2816.020 168.940 ;
        RECT 2815.760 37.780 2816.020 38.040 ;
        RECT 2821.740 37.780 2822.000 38.040 ;
      LAYER met2 ;
        RECT 1937.290 510.410 1937.570 514.000 ;
        RECT 1937.290 510.270 1938.740 510.410 ;
        RECT 1937.290 510.000 1937.570 510.270 ;
        RECT 1938.600 168.970 1938.740 510.270 ;
        RECT 1938.540 168.650 1938.800 168.970 ;
        RECT 2815.760 168.650 2816.020 168.970 ;
        RECT 2815.820 38.070 2815.960 168.650 ;
        RECT 2815.760 37.750 2816.020 38.070 ;
        RECT 2821.740 37.750 2822.000 38.070 ;
        RECT 2821.800 2.400 2821.940 37.750 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 58.720 1952.630 58.780 ;
        RECT 2839.190 58.720 2839.510 58.780 ;
        RECT 1952.310 58.580 2839.510 58.720 ;
        RECT 1952.310 58.520 1952.630 58.580 ;
        RECT 2839.190 58.520 2839.510 58.580 ;
      LAYER via ;
        RECT 1952.340 58.520 1952.600 58.780 ;
        RECT 2839.220 58.520 2839.480 58.780 ;
      LAYER met2 ;
        RECT 1949.710 510.410 1949.990 514.000 ;
        RECT 1949.710 510.270 1952.540 510.410 ;
        RECT 1949.710 510.000 1949.990 510.270 ;
        RECT 1952.400 58.810 1952.540 510.270 ;
        RECT 1952.340 58.490 1952.600 58.810 ;
        RECT 2839.220 58.490 2839.480 58.810 ;
        RECT 2839.280 2.400 2839.420 58.490 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1961.970 500.720 1962.290 500.780 ;
        RECT 2231.990 500.720 2232.310 500.780 ;
        RECT 1961.970 500.580 2232.310 500.720 ;
        RECT 1961.970 500.520 1962.290 500.580 ;
        RECT 2231.990 500.520 2232.310 500.580 ;
        RECT 2231.990 100.200 2232.310 100.260 ;
        RECT 2857.130 100.200 2857.450 100.260 ;
        RECT 2231.990 100.060 2857.450 100.200 ;
        RECT 2231.990 100.000 2232.310 100.060 ;
        RECT 2857.130 100.000 2857.450 100.060 ;
      LAYER via ;
        RECT 1962.000 500.520 1962.260 500.780 ;
        RECT 2232.020 500.520 2232.280 500.780 ;
        RECT 2232.020 100.000 2232.280 100.260 ;
        RECT 2857.160 100.000 2857.420 100.260 ;
      LAYER met2 ;
        RECT 1962.130 510.340 1962.410 514.000 ;
        RECT 1962.060 510.000 1962.410 510.340 ;
        RECT 1962.060 500.810 1962.200 510.000 ;
        RECT 1962.000 500.490 1962.260 500.810 ;
        RECT 2232.020 500.490 2232.280 500.810 ;
        RECT 2232.080 100.290 2232.220 500.490 ;
        RECT 2232.020 99.970 2232.280 100.290 ;
        RECT 2857.160 99.970 2857.420 100.290 ;
        RECT 2857.220 2.400 2857.360 99.970 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1974.390 472.500 1974.710 472.560 ;
        RECT 2870.470 472.500 2870.790 472.560 ;
        RECT 1974.390 472.360 2870.790 472.500 ;
        RECT 1974.390 472.300 1974.710 472.360 ;
        RECT 2870.470 472.300 2870.790 472.360 ;
      LAYER via ;
        RECT 1974.420 472.300 1974.680 472.560 ;
        RECT 2870.500 472.300 2870.760 472.560 ;
      LAYER met2 ;
        RECT 1974.550 510.340 1974.830 514.000 ;
        RECT 1974.480 510.000 1974.830 510.340 ;
        RECT 1974.480 472.590 1974.620 510.000 ;
        RECT 1974.420 472.270 1974.680 472.590 ;
        RECT 2870.500 472.270 2870.760 472.590 ;
        RECT 2870.560 18.090 2870.700 472.270 ;
        RECT 2870.560 17.950 2875.300 18.090 ;
        RECT 2875.160 2.400 2875.300 17.950 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2839.265 193.205 2839.435 241.315 ;
        RECT 2840.185 89.845 2840.355 137.955 ;
      LAYER mcon ;
        RECT 2839.265 241.145 2839.435 241.315 ;
        RECT 2840.185 137.785 2840.355 137.955 ;
      LAYER met1 ;
        RECT 1986.810 251.840 1987.130 251.900 ;
        RECT 2839.650 251.840 2839.970 251.900 ;
        RECT 1986.810 251.700 2839.970 251.840 ;
        RECT 1986.810 251.640 1987.130 251.700 ;
        RECT 2839.650 251.640 2839.970 251.700 ;
        RECT 2839.205 241.300 2839.495 241.345 ;
        RECT 2839.650 241.300 2839.970 241.360 ;
        RECT 2839.205 241.160 2839.970 241.300 ;
        RECT 2839.205 241.115 2839.495 241.160 ;
        RECT 2839.650 241.100 2839.970 241.160 ;
        RECT 2839.190 193.360 2839.510 193.420 ;
        RECT 2838.995 193.220 2839.510 193.360 ;
        RECT 2839.190 193.160 2839.510 193.220 ;
        RECT 2839.190 158.680 2839.510 158.740 ;
        RECT 2840.110 158.680 2840.430 158.740 ;
        RECT 2839.190 158.540 2840.430 158.680 ;
        RECT 2839.190 158.480 2839.510 158.540 ;
        RECT 2840.110 158.480 2840.430 158.540 ;
        RECT 2840.110 137.940 2840.430 138.000 ;
        RECT 2839.915 137.800 2840.430 137.940 ;
        RECT 2840.110 137.740 2840.430 137.800 ;
        RECT 2840.110 90.000 2840.430 90.060 ;
        RECT 2839.915 89.860 2840.430 90.000 ;
        RECT 2840.110 89.800 2840.430 89.860 ;
        RECT 2841.030 17.920 2841.350 17.980 ;
        RECT 2841.030 17.780 2863.800 17.920 ;
        RECT 2841.030 17.720 2841.350 17.780 ;
        RECT 2863.660 17.580 2863.800 17.780 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2863.660 17.440 2893.330 17.580 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 1986.840 251.640 1987.100 251.900 ;
        RECT 2839.680 251.640 2839.940 251.900 ;
        RECT 2839.680 241.100 2839.940 241.360 ;
        RECT 2839.220 193.160 2839.480 193.420 ;
        RECT 2839.220 158.480 2839.480 158.740 ;
        RECT 2840.140 158.480 2840.400 158.740 ;
        RECT 2840.140 137.740 2840.400 138.000 ;
        RECT 2840.140 89.800 2840.400 90.060 ;
        RECT 2841.060 17.720 2841.320 17.980 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 1986.970 510.340 1987.250 514.000 ;
        RECT 1986.900 510.000 1987.250 510.340 ;
        RECT 1986.900 251.930 1987.040 510.000 ;
        RECT 1986.840 251.610 1987.100 251.930 ;
        RECT 2839.680 251.610 2839.940 251.930 ;
        RECT 2839.740 241.390 2839.880 251.610 ;
        RECT 2839.680 241.070 2839.940 241.390 ;
        RECT 2839.220 193.130 2839.480 193.450 ;
        RECT 2839.280 158.770 2839.420 193.130 ;
        RECT 2839.220 158.450 2839.480 158.770 ;
        RECT 2840.140 158.450 2840.400 158.770 ;
        RECT 2840.200 138.030 2840.340 158.450 ;
        RECT 2840.140 137.710 2840.400 138.030 ;
        RECT 2840.140 89.770 2840.400 90.090 ;
        RECT 2840.200 41.325 2840.340 89.770 ;
        RECT 2840.130 40.955 2840.410 41.325 ;
        RECT 2841.050 40.275 2841.330 40.645 ;
        RECT 2841.120 18.010 2841.260 40.275 ;
        RECT 2841.060 17.690 2841.320 18.010 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 2840.130 41.000 2840.410 41.280 ;
        RECT 2841.050 40.320 2841.330 40.600 ;
      LAYER met3 ;
        RECT 2840.105 41.290 2840.435 41.305 ;
        RECT 2839.430 40.990 2840.435 41.290 ;
        RECT 2839.430 40.610 2839.730 40.990 ;
        RECT 2840.105 40.975 2840.435 40.990 ;
        RECT 2841.025 40.610 2841.355 40.625 ;
        RECT 2839.430 40.310 2841.355 40.610 ;
        RECT 2841.025 40.295 2841.355 40.310 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2432.625 17.085 2432.795 36.635 ;
        RECT 2497.945 16.405 2498.115 17.255 ;
        RECT 2545.785 16.405 2545.955 17.595 ;
        RECT 2559.585 17.425 2560.215 17.595 ;
        RECT 2560.045 17.085 2560.215 17.425 ;
        RECT 2594.545 17.085 2594.715 17.935 ;
        RECT 2642.385 17.085 2642.555 17.935 ;
        RECT 2795.105 16.405 2795.275 17.595 ;
      LAYER mcon ;
        RECT 2432.625 36.465 2432.795 36.635 ;
        RECT 2594.545 17.765 2594.715 17.935 ;
        RECT 2545.785 17.425 2545.955 17.595 ;
        RECT 2497.945 17.085 2498.115 17.255 ;
        RECT 2642.385 17.765 2642.555 17.935 ;
        RECT 2795.105 17.425 2795.275 17.595 ;
      LAYER met1 ;
        RECT 2000.150 417.760 2000.470 417.820 ;
        RECT 2411.390 417.760 2411.710 417.820 ;
        RECT 2000.150 417.620 2411.710 417.760 ;
        RECT 2000.150 417.560 2000.470 417.620 ;
        RECT 2411.390 417.560 2411.710 417.620 ;
        RECT 2410.930 36.620 2411.250 36.680 ;
        RECT 2432.565 36.620 2432.855 36.665 ;
        RECT 2410.930 36.480 2432.855 36.620 ;
        RECT 2410.930 36.420 2411.250 36.480 ;
        RECT 2432.565 36.435 2432.855 36.480 ;
        RECT 2594.485 17.920 2594.775 17.965 ;
        RECT 2642.325 17.920 2642.615 17.965 ;
        RECT 2594.485 17.780 2642.615 17.920 ;
        RECT 2594.485 17.735 2594.775 17.780 ;
        RECT 2642.325 17.735 2642.615 17.780 ;
        RECT 2545.725 17.580 2546.015 17.625 ;
        RECT 2559.525 17.580 2559.815 17.625 ;
        RECT 2795.045 17.580 2795.335 17.625 ;
        RECT 2545.725 17.440 2559.815 17.580 ;
        RECT 2545.725 17.395 2546.015 17.440 ;
        RECT 2559.525 17.395 2559.815 17.440 ;
        RECT 2649.300 17.440 2795.335 17.580 ;
        RECT 2432.565 17.240 2432.855 17.285 ;
        RECT 2497.885 17.240 2498.175 17.285 ;
        RECT 2432.565 17.100 2498.175 17.240 ;
        RECT 2432.565 17.055 2432.855 17.100 ;
        RECT 2497.885 17.055 2498.175 17.100 ;
        RECT 2559.985 17.240 2560.275 17.285 ;
        RECT 2594.485 17.240 2594.775 17.285 ;
        RECT 2559.985 17.100 2594.775 17.240 ;
        RECT 2559.985 17.055 2560.275 17.100 ;
        RECT 2594.485 17.055 2594.775 17.100 ;
        RECT 2642.325 17.240 2642.615 17.285 ;
        RECT 2649.300 17.240 2649.440 17.440 ;
        RECT 2795.045 17.395 2795.335 17.440 ;
        RECT 2642.325 17.100 2649.440 17.240 ;
        RECT 2642.325 17.055 2642.615 17.100 ;
        RECT 2497.885 16.560 2498.175 16.605 ;
        RECT 2545.725 16.560 2546.015 16.605 ;
        RECT 2497.885 16.420 2546.015 16.560 ;
        RECT 2497.885 16.375 2498.175 16.420 ;
        RECT 2545.725 16.375 2546.015 16.420 ;
        RECT 2795.045 16.560 2795.335 16.605 ;
        RECT 2910.950 16.560 2911.270 16.620 ;
        RECT 2795.045 16.420 2911.270 16.560 ;
        RECT 2795.045 16.375 2795.335 16.420 ;
        RECT 2910.950 16.360 2911.270 16.420 ;
      LAYER via ;
        RECT 2000.180 417.560 2000.440 417.820 ;
        RECT 2411.420 417.560 2411.680 417.820 ;
        RECT 2410.960 36.420 2411.220 36.680 ;
        RECT 2910.980 16.360 2911.240 16.620 ;
      LAYER met2 ;
        RECT 1999.390 510.410 1999.670 514.000 ;
        RECT 1999.390 510.270 2000.380 510.410 ;
        RECT 1999.390 510.000 1999.670 510.270 ;
        RECT 2000.240 417.850 2000.380 510.270 ;
        RECT 2000.180 417.530 2000.440 417.850 ;
        RECT 2411.420 417.530 2411.680 417.850 ;
        RECT 2411.480 45.970 2411.620 417.530 ;
        RECT 2411.020 45.830 2411.620 45.970 ;
        RECT 2411.020 36.710 2411.160 45.830 ;
        RECT 2410.960 36.390 2411.220 36.710 ;
        RECT 2910.980 16.330 2911.240 16.650 ;
        RECT 2911.040 2.400 2911.180 16.330 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.210 320.860 579.530 320.920 ;
        RECT 855.670 320.860 855.990 320.920 ;
        RECT 579.210 320.720 855.990 320.860 ;
        RECT 579.210 320.660 579.530 320.720 ;
        RECT 855.670 320.660 855.990 320.720 ;
      LAYER via ;
        RECT 579.240 320.660 579.500 320.920 ;
        RECT 855.700 320.660 855.960 320.920 ;
      LAYER met2 ;
        RECT 576.610 510.410 576.890 514.000 ;
        RECT 576.610 510.270 579.440 510.410 ;
        RECT 576.610 510.000 576.890 510.270 ;
        RECT 579.300 320.950 579.440 510.270 ;
        RECT 579.240 320.630 579.500 320.950 ;
        RECT 855.700 320.630 855.960 320.950 ;
        RECT 855.760 17.410 855.900 320.630 ;
        RECT 855.760 17.270 859.120 17.410 ;
        RECT 858.980 2.400 859.120 17.270 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 588.870 496.980 589.190 497.040 ;
        RECT 592.550 496.980 592.870 497.040 ;
        RECT 588.870 496.840 592.870 496.980 ;
        RECT 588.870 496.780 589.190 496.840 ;
        RECT 592.550 496.780 592.870 496.840 ;
        RECT 592.550 334.460 592.870 334.520 ;
        RECT 876.370 334.460 876.690 334.520 ;
        RECT 592.550 334.320 876.690 334.460 ;
        RECT 592.550 334.260 592.870 334.320 ;
        RECT 876.370 334.260 876.690 334.320 ;
      LAYER via ;
        RECT 588.900 496.780 589.160 497.040 ;
        RECT 592.580 496.780 592.840 497.040 ;
        RECT 592.580 334.260 592.840 334.520 ;
        RECT 876.400 334.260 876.660 334.520 ;
      LAYER met2 ;
        RECT 589.030 510.340 589.310 514.000 ;
        RECT 588.960 510.000 589.310 510.340 ;
        RECT 588.960 497.070 589.100 510.000 ;
        RECT 588.900 496.750 589.160 497.070 ;
        RECT 592.580 496.750 592.840 497.070 ;
        RECT 592.640 334.550 592.780 496.750 ;
        RECT 592.580 334.230 592.840 334.550 ;
        RECT 876.400 334.230 876.660 334.550 ;
        RECT 876.460 17.410 876.600 334.230 ;
        RECT 876.460 17.270 877.060 17.410 ;
        RECT 876.920 2.400 877.060 17.270 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 601.290 496.980 601.610 497.040 ;
        RECT 606.350 496.980 606.670 497.040 ;
        RECT 601.290 496.840 606.670 496.980 ;
        RECT 601.290 496.780 601.610 496.840 ;
        RECT 606.350 496.780 606.670 496.840 ;
        RECT 606.350 341.600 606.670 341.660 ;
        RECT 890.170 341.600 890.490 341.660 ;
        RECT 606.350 341.460 890.490 341.600 ;
        RECT 606.350 341.400 606.670 341.460 ;
        RECT 890.170 341.400 890.490 341.460 ;
      LAYER via ;
        RECT 601.320 496.780 601.580 497.040 ;
        RECT 606.380 496.780 606.640 497.040 ;
        RECT 606.380 341.400 606.640 341.660 ;
        RECT 890.200 341.400 890.460 341.660 ;
      LAYER met2 ;
        RECT 601.450 510.340 601.730 514.000 ;
        RECT 601.380 510.000 601.730 510.340 ;
        RECT 601.380 497.070 601.520 510.000 ;
        RECT 601.320 496.750 601.580 497.070 ;
        RECT 606.380 496.750 606.640 497.070 ;
        RECT 606.440 341.690 606.580 496.750 ;
        RECT 606.380 341.370 606.640 341.690 ;
        RECT 890.200 341.370 890.460 341.690 ;
        RECT 890.260 18.090 890.400 341.370 ;
        RECT 890.260 17.950 895.000 18.090 ;
        RECT 894.860 2.400 895.000 17.950 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.250 348.400 613.570 348.460 ;
        RECT 910.870 348.400 911.190 348.460 ;
        RECT 613.250 348.260 911.190 348.400 ;
        RECT 613.250 348.200 613.570 348.260 ;
        RECT 910.870 348.200 911.190 348.260 ;
      LAYER via ;
        RECT 613.280 348.200 613.540 348.460 ;
        RECT 910.900 348.200 911.160 348.460 ;
      LAYER met2 ;
        RECT 613.870 510.410 614.150 514.000 ;
        RECT 613.340 510.270 614.150 510.410 ;
        RECT 613.340 348.490 613.480 510.270 ;
        RECT 613.870 510.000 614.150 510.270 ;
        RECT 613.280 348.170 613.540 348.490 ;
        RECT 910.900 348.170 911.160 348.490 ;
        RECT 910.960 17.410 911.100 348.170 ;
        RECT 910.960 17.270 912.940 17.410 ;
        RECT 912.800 2.400 912.940 17.270 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 355.200 627.370 355.260 ;
        RECT 924.670 355.200 924.990 355.260 ;
        RECT 627.050 355.060 924.990 355.200 ;
        RECT 627.050 355.000 627.370 355.060 ;
        RECT 924.670 355.000 924.990 355.060 ;
      LAYER via ;
        RECT 627.080 355.000 627.340 355.260 ;
        RECT 924.700 355.000 924.960 355.260 ;
      LAYER met2 ;
        RECT 626.290 510.410 626.570 514.000 ;
        RECT 626.290 510.270 627.280 510.410 ;
        RECT 626.290 510.000 626.570 510.270 ;
        RECT 627.140 355.290 627.280 510.270 ;
        RECT 627.080 354.970 627.340 355.290 ;
        RECT 924.700 354.970 924.960 355.290 ;
        RECT 924.760 17.410 924.900 354.970 ;
        RECT 924.760 17.270 930.420 17.410 ;
        RECT 930.280 2.400 930.420 17.270 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 641.310 375.940 641.630 376.000 ;
        RECT 945.370 375.940 945.690 376.000 ;
        RECT 641.310 375.800 945.690 375.940 ;
        RECT 641.310 375.740 641.630 375.800 ;
        RECT 945.370 375.740 945.690 375.800 ;
      LAYER via ;
        RECT 641.340 375.740 641.600 376.000 ;
        RECT 945.400 375.740 945.660 376.000 ;
      LAYER met2 ;
        RECT 638.710 510.410 638.990 514.000 ;
        RECT 638.710 510.270 641.540 510.410 ;
        RECT 638.710 510.000 638.990 510.270 ;
        RECT 641.400 376.030 641.540 510.270 ;
        RECT 641.340 375.710 641.600 376.030 ;
        RECT 945.400 375.710 945.660 376.030 ;
        RECT 945.460 17.410 945.600 375.710 ;
        RECT 945.460 17.270 948.360 17.410 ;
        RECT 948.220 2.400 948.360 17.270 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.510 496.980 650.830 497.040 ;
        RECT 655.110 496.980 655.430 497.040 ;
        RECT 650.510 496.840 655.430 496.980 ;
        RECT 650.510 496.780 650.830 496.840 ;
        RECT 655.110 496.780 655.430 496.840 ;
        RECT 655.110 382.740 655.430 382.800 ;
        RECT 966.070 382.740 966.390 382.800 ;
        RECT 655.110 382.600 966.390 382.740 ;
        RECT 655.110 382.540 655.430 382.600 ;
        RECT 966.070 382.540 966.390 382.600 ;
      LAYER via ;
        RECT 650.540 496.780 650.800 497.040 ;
        RECT 655.140 496.780 655.400 497.040 ;
        RECT 655.140 382.540 655.400 382.800 ;
        RECT 966.100 382.540 966.360 382.800 ;
      LAYER met2 ;
        RECT 650.670 510.340 650.950 514.000 ;
        RECT 650.600 510.000 650.950 510.340 ;
        RECT 650.600 497.070 650.740 510.000 ;
        RECT 650.540 496.750 650.800 497.070 ;
        RECT 655.140 496.750 655.400 497.070 ;
        RECT 655.200 382.830 655.340 496.750 ;
        RECT 655.140 382.510 655.400 382.830 ;
        RECT 966.100 382.510 966.360 382.830 ;
        RECT 966.160 2.400 966.300 382.510 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 496.980 663.250 497.040 ;
        RECT 668.910 496.980 669.230 497.040 ;
        RECT 662.930 496.840 669.230 496.980 ;
        RECT 662.930 496.780 663.250 496.840 ;
        RECT 668.910 496.780 669.230 496.840 ;
        RECT 668.910 389.880 669.230 389.940 ;
        RECT 979.870 389.880 980.190 389.940 ;
        RECT 668.910 389.740 980.190 389.880 ;
        RECT 668.910 389.680 669.230 389.740 ;
        RECT 979.870 389.680 980.190 389.740 ;
        RECT 979.870 62.120 980.190 62.180 ;
        RECT 984.010 62.120 984.330 62.180 ;
        RECT 979.870 61.980 984.330 62.120 ;
        RECT 979.870 61.920 980.190 61.980 ;
        RECT 984.010 61.920 984.330 61.980 ;
      LAYER via ;
        RECT 662.960 496.780 663.220 497.040 ;
        RECT 668.940 496.780 669.200 497.040 ;
        RECT 668.940 389.680 669.200 389.940 ;
        RECT 979.900 389.680 980.160 389.940 ;
        RECT 979.900 61.920 980.160 62.180 ;
        RECT 984.040 61.920 984.300 62.180 ;
      LAYER met2 ;
        RECT 663.090 510.340 663.370 514.000 ;
        RECT 663.020 510.000 663.370 510.340 ;
        RECT 663.020 497.070 663.160 510.000 ;
        RECT 662.960 496.750 663.220 497.070 ;
        RECT 668.940 496.750 669.200 497.070 ;
        RECT 669.000 389.970 669.140 496.750 ;
        RECT 668.940 389.650 669.200 389.970 ;
        RECT 979.900 389.650 980.160 389.970 ;
        RECT 979.960 62.210 980.100 389.650 ;
        RECT 979.900 61.890 980.160 62.210 ;
        RECT 984.040 61.890 984.300 62.210 ;
        RECT 984.100 2.400 984.240 61.890 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 19.960 441.530 20.020 ;
        RECT 662.930 19.960 663.250 20.020 ;
        RECT 441.210 19.820 663.250 19.960 ;
        RECT 441.210 19.760 441.530 19.820 ;
        RECT 662.930 19.760 663.250 19.820 ;
      LAYER via ;
        RECT 441.240 19.760 441.500 20.020 ;
        RECT 662.960 19.760 663.220 20.020 ;
      LAYER met2 ;
        RECT 440.450 510.410 440.730 514.000 ;
        RECT 440.450 510.270 441.440 510.410 ;
        RECT 440.450 510.000 440.730 510.270 ;
        RECT 441.300 20.050 441.440 510.270 ;
        RECT 441.240 19.730 441.500 20.050 ;
        RECT 662.960 19.730 663.220 20.050 ;
        RECT 663.020 2.400 663.160 19.730 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1000.645 282.965 1000.815 331.075 ;
        RECT 1000.645 186.405 1000.815 234.515 ;
        RECT 1000.645 48.365 1000.815 114.155 ;
      LAYER mcon ;
        RECT 1000.645 330.905 1000.815 331.075 ;
        RECT 1000.645 234.345 1000.815 234.515 ;
        RECT 1000.645 113.985 1000.815 114.155 ;
      LAYER met1 ;
        RECT 675.350 396.680 675.670 396.740 ;
        RECT 1000.570 396.680 1000.890 396.740 ;
        RECT 675.350 396.540 1000.890 396.680 ;
        RECT 675.350 396.480 675.670 396.540 ;
        RECT 1000.570 396.480 1000.890 396.540 ;
        RECT 1000.570 331.060 1000.890 331.120 ;
        RECT 1000.375 330.920 1000.890 331.060 ;
        RECT 1000.570 330.860 1000.890 330.920 ;
        RECT 1000.570 283.120 1000.890 283.180 ;
        RECT 1000.375 282.980 1000.890 283.120 ;
        RECT 1000.570 282.920 1000.890 282.980 ;
        RECT 1000.570 234.500 1000.890 234.560 ;
        RECT 1000.375 234.360 1000.890 234.500 ;
        RECT 1000.570 234.300 1000.890 234.360 ;
        RECT 1000.570 186.560 1000.890 186.620 ;
        RECT 1000.375 186.420 1000.890 186.560 ;
        RECT 1000.570 186.360 1000.890 186.420 ;
        RECT 1000.570 114.140 1000.890 114.200 ;
        RECT 1000.375 114.000 1000.890 114.140 ;
        RECT 1000.570 113.940 1000.890 114.000 ;
        RECT 1000.585 48.520 1000.875 48.565 ;
        RECT 1001.950 48.520 1002.270 48.580 ;
        RECT 1000.585 48.380 1002.270 48.520 ;
        RECT 1000.585 48.335 1000.875 48.380 ;
        RECT 1001.950 48.320 1002.270 48.380 ;
        RECT 1001.950 2.960 1002.270 3.020 ;
        RECT 1002.410 2.960 1002.730 3.020 ;
        RECT 1001.950 2.820 1002.730 2.960 ;
        RECT 1001.950 2.760 1002.270 2.820 ;
        RECT 1002.410 2.760 1002.730 2.820 ;
      LAYER via ;
        RECT 675.380 396.480 675.640 396.740 ;
        RECT 1000.600 396.480 1000.860 396.740 ;
        RECT 1000.600 330.860 1000.860 331.120 ;
        RECT 1000.600 282.920 1000.860 283.180 ;
        RECT 1000.600 234.300 1000.860 234.560 ;
        RECT 1000.600 186.360 1000.860 186.620 ;
        RECT 1000.600 113.940 1000.860 114.200 ;
        RECT 1001.980 48.320 1002.240 48.580 ;
        RECT 1001.980 2.760 1002.240 3.020 ;
        RECT 1002.440 2.760 1002.700 3.020 ;
      LAYER met2 ;
        RECT 675.510 510.340 675.790 514.000 ;
        RECT 675.440 510.000 675.790 510.340 ;
        RECT 675.440 396.770 675.580 510.000 ;
        RECT 675.380 396.450 675.640 396.770 ;
        RECT 1000.600 396.450 1000.860 396.770 ;
        RECT 1000.660 331.150 1000.800 396.450 ;
        RECT 1000.600 330.830 1000.860 331.150 ;
        RECT 1000.600 282.890 1000.860 283.210 ;
        RECT 1000.660 234.590 1000.800 282.890 ;
        RECT 1000.600 234.270 1000.860 234.590 ;
        RECT 1000.600 186.330 1000.860 186.650 ;
        RECT 1000.660 114.230 1000.800 186.330 ;
        RECT 1000.600 113.910 1000.860 114.230 ;
        RECT 1001.980 48.290 1002.240 48.610 ;
        RECT 1002.040 48.010 1002.180 48.290 ;
        RECT 1002.040 47.870 1002.640 48.010 ;
        RECT 1002.500 3.050 1002.640 47.870 ;
        RECT 1001.980 2.730 1002.240 3.050 ;
        RECT 1002.440 2.730 1002.700 3.050 ;
        RECT 1002.040 2.400 1002.180 2.730 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.150 403.480 689.470 403.540 ;
        RECT 1014.370 403.480 1014.690 403.540 ;
        RECT 689.150 403.340 1014.690 403.480 ;
        RECT 689.150 403.280 689.470 403.340 ;
        RECT 1014.370 403.280 1014.690 403.340 ;
        RECT 1014.370 62.120 1014.690 62.180 ;
        RECT 1019.430 62.120 1019.750 62.180 ;
        RECT 1014.370 61.980 1019.750 62.120 ;
        RECT 1014.370 61.920 1014.690 61.980 ;
        RECT 1019.430 61.920 1019.750 61.980 ;
      LAYER via ;
        RECT 689.180 403.280 689.440 403.540 ;
        RECT 1014.400 403.280 1014.660 403.540 ;
        RECT 1014.400 61.920 1014.660 62.180 ;
        RECT 1019.460 61.920 1019.720 62.180 ;
      LAYER met2 ;
        RECT 687.930 510.410 688.210 514.000 ;
        RECT 687.930 510.270 689.380 510.410 ;
        RECT 687.930 510.000 688.210 510.270 ;
        RECT 689.240 403.570 689.380 510.270 ;
        RECT 689.180 403.250 689.440 403.570 ;
        RECT 1014.400 403.250 1014.660 403.570 ;
        RECT 1014.460 62.210 1014.600 403.250 ;
        RECT 1014.400 61.890 1014.660 62.210 ;
        RECT 1019.460 61.890 1019.720 62.210 ;
        RECT 1019.520 2.400 1019.660 61.890 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 410.960 703.730 411.020 ;
        RECT 1035.070 410.960 1035.390 411.020 ;
        RECT 703.410 410.820 1035.390 410.960 ;
        RECT 703.410 410.760 703.730 410.820 ;
        RECT 1035.070 410.760 1035.390 410.820 ;
      LAYER via ;
        RECT 703.440 410.760 703.700 411.020 ;
        RECT 1035.100 410.760 1035.360 411.020 ;
      LAYER met2 ;
        RECT 700.350 510.410 700.630 514.000 ;
        RECT 700.350 510.270 703.640 510.410 ;
        RECT 700.350 510.000 700.630 510.270 ;
        RECT 703.500 411.050 703.640 510.270 ;
        RECT 703.440 410.730 703.700 411.050 ;
        RECT 1035.100 410.730 1035.360 411.050 ;
        RECT 1035.160 16.730 1035.300 410.730 ;
        RECT 1035.160 16.590 1037.600 16.730 ;
        RECT 1037.460 2.400 1037.600 16.590 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 712.610 496.980 712.930 497.040 ;
        RECT 716.750 496.980 717.070 497.040 ;
        RECT 712.610 496.840 717.070 496.980 ;
        RECT 712.610 496.780 712.930 496.840 ;
        RECT 716.750 496.780 717.070 496.840 ;
        RECT 716.750 431.360 717.070 431.420 ;
        RECT 1048.870 431.360 1049.190 431.420 ;
        RECT 716.750 431.220 1049.190 431.360 ;
        RECT 716.750 431.160 717.070 431.220 ;
        RECT 1048.870 431.160 1049.190 431.220 ;
        RECT 1048.870 17.580 1049.190 17.640 ;
        RECT 1055.310 17.580 1055.630 17.640 ;
        RECT 1048.870 17.440 1055.630 17.580 ;
        RECT 1048.870 17.380 1049.190 17.440 ;
        RECT 1055.310 17.380 1055.630 17.440 ;
      LAYER via ;
        RECT 712.640 496.780 712.900 497.040 ;
        RECT 716.780 496.780 717.040 497.040 ;
        RECT 716.780 431.160 717.040 431.420 ;
        RECT 1048.900 431.160 1049.160 431.420 ;
        RECT 1048.900 17.380 1049.160 17.640 ;
        RECT 1055.340 17.380 1055.600 17.640 ;
      LAYER met2 ;
        RECT 712.770 510.340 713.050 514.000 ;
        RECT 712.700 510.000 713.050 510.340 ;
        RECT 712.700 497.070 712.840 510.000 ;
        RECT 712.640 496.750 712.900 497.070 ;
        RECT 716.780 496.750 717.040 497.070 ;
        RECT 716.840 431.450 716.980 496.750 ;
        RECT 716.780 431.130 717.040 431.450 ;
        RECT 1048.900 431.130 1049.160 431.450 ;
        RECT 1048.960 17.670 1049.100 431.130 ;
        RECT 1048.900 17.350 1049.160 17.670 ;
        RECT 1055.340 17.350 1055.600 17.670 ;
        RECT 1055.400 2.400 1055.540 17.350 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 725.030 496.980 725.350 497.040 ;
        RECT 730.550 496.980 730.870 497.040 ;
        RECT 725.030 496.840 730.870 496.980 ;
        RECT 725.030 496.780 725.350 496.840 ;
        RECT 730.550 496.780 730.870 496.840 ;
        RECT 730.550 438.500 730.870 438.560 ;
        RECT 1069.570 438.500 1069.890 438.560 ;
        RECT 730.550 438.360 1069.890 438.500 ;
        RECT 730.550 438.300 730.870 438.360 ;
        RECT 1069.570 438.300 1069.890 438.360 ;
      LAYER via ;
        RECT 725.060 496.780 725.320 497.040 ;
        RECT 730.580 496.780 730.840 497.040 ;
        RECT 730.580 438.300 730.840 438.560 ;
        RECT 1069.600 438.300 1069.860 438.560 ;
      LAYER met2 ;
        RECT 725.190 510.340 725.470 514.000 ;
        RECT 725.120 510.000 725.470 510.340 ;
        RECT 725.120 497.070 725.260 510.000 ;
        RECT 725.060 496.750 725.320 497.070 ;
        RECT 730.580 496.750 730.840 497.070 ;
        RECT 730.640 438.590 730.780 496.750 ;
        RECT 730.580 438.270 730.840 438.590 ;
        RECT 1069.600 438.270 1069.860 438.590 ;
        RECT 1069.660 17.410 1069.800 438.270 ;
        RECT 1069.660 17.270 1073.480 17.410 ;
        RECT 1073.340 2.400 1073.480 17.270 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.450 465.700 737.770 465.760 ;
        RECT 1090.270 465.700 1090.590 465.760 ;
        RECT 737.450 465.560 1090.590 465.700 ;
        RECT 737.450 465.500 737.770 465.560 ;
        RECT 1090.270 465.500 1090.590 465.560 ;
      LAYER via ;
        RECT 737.480 465.500 737.740 465.760 ;
        RECT 1090.300 465.500 1090.560 465.760 ;
      LAYER met2 ;
        RECT 737.610 510.340 737.890 514.000 ;
        RECT 737.540 510.000 737.890 510.340 ;
        RECT 737.540 465.790 737.680 510.000 ;
        RECT 737.480 465.470 737.740 465.790 ;
        RECT 1090.300 465.470 1090.560 465.790 ;
        RECT 1090.360 17.410 1090.500 465.470 ;
        RECT 1090.360 17.270 1090.960 17.410 ;
        RECT 1090.820 2.400 1090.960 17.270 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 749.870 479.640 750.190 479.700 ;
        RECT 1104.070 479.640 1104.390 479.700 ;
        RECT 749.870 479.500 1104.390 479.640 ;
        RECT 749.870 479.440 750.190 479.500 ;
        RECT 1104.070 479.440 1104.390 479.500 ;
      LAYER via ;
        RECT 749.900 479.440 750.160 479.700 ;
        RECT 1104.100 479.440 1104.360 479.700 ;
      LAYER met2 ;
        RECT 750.030 510.340 750.310 514.000 ;
        RECT 749.960 510.000 750.310 510.340 ;
        RECT 749.960 479.730 750.100 510.000 ;
        RECT 749.900 479.410 750.160 479.730 ;
        RECT 1104.100 479.410 1104.360 479.730 ;
        RECT 1104.160 17.410 1104.300 479.410 ;
        RECT 1104.160 17.270 1108.900 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 761.830 500.720 762.150 500.780 ;
        RECT 765.510 500.720 765.830 500.780 ;
        RECT 761.830 500.580 765.830 500.720 ;
        RECT 761.830 500.520 762.150 500.580 ;
        RECT 765.510 500.520 765.830 500.580 ;
        RECT 765.510 459.240 765.830 459.300 ;
        RECT 1124.770 459.240 1125.090 459.300 ;
        RECT 765.510 459.100 1125.090 459.240 ;
        RECT 765.510 459.040 765.830 459.100 ;
        RECT 1124.770 459.040 1125.090 459.100 ;
      LAYER via ;
        RECT 761.860 500.520 762.120 500.780 ;
        RECT 765.540 500.520 765.800 500.780 ;
        RECT 765.540 459.040 765.800 459.300 ;
        RECT 1124.800 459.040 1125.060 459.300 ;
      LAYER met2 ;
        RECT 761.990 510.340 762.270 514.000 ;
        RECT 761.920 510.000 762.270 510.340 ;
        RECT 761.920 500.810 762.060 510.000 ;
        RECT 761.860 500.490 762.120 500.810 ;
        RECT 765.540 500.490 765.800 500.810 ;
        RECT 765.600 459.330 765.740 500.490 ;
        RECT 765.540 459.010 765.800 459.330 ;
        RECT 1124.800 459.010 1125.060 459.330 ;
        RECT 1124.860 17.410 1125.000 459.010 ;
        RECT 1124.860 17.270 1126.840 17.410 ;
        RECT 1126.700 2.400 1126.840 17.270 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 774.250 503.440 774.570 503.500 ;
        RECT 778.850 503.440 779.170 503.500 ;
        RECT 774.250 503.300 779.170 503.440 ;
        RECT 774.250 503.240 774.570 503.300 ;
        RECT 778.850 503.240 779.170 503.300 ;
        RECT 778.850 452.100 779.170 452.160 ;
        RECT 1138.570 452.100 1138.890 452.160 ;
        RECT 778.850 451.960 1138.890 452.100 ;
        RECT 778.850 451.900 779.170 451.960 ;
        RECT 1138.570 451.900 1138.890 451.960 ;
        RECT 1138.570 17.920 1138.890 17.980 ;
        RECT 1144.550 17.920 1144.870 17.980 ;
        RECT 1138.570 17.780 1144.870 17.920 ;
        RECT 1138.570 17.720 1138.890 17.780 ;
        RECT 1144.550 17.720 1144.870 17.780 ;
      LAYER via ;
        RECT 774.280 503.240 774.540 503.500 ;
        RECT 778.880 503.240 779.140 503.500 ;
        RECT 778.880 451.900 779.140 452.160 ;
        RECT 1138.600 451.900 1138.860 452.160 ;
        RECT 1138.600 17.720 1138.860 17.980 ;
        RECT 1144.580 17.720 1144.840 17.980 ;
      LAYER met2 ;
        RECT 774.410 510.340 774.690 514.000 ;
        RECT 774.340 510.000 774.690 510.340 ;
        RECT 774.340 503.530 774.480 510.000 ;
        RECT 774.280 503.210 774.540 503.530 ;
        RECT 778.880 503.210 779.140 503.530 ;
        RECT 778.940 452.190 779.080 503.210 ;
        RECT 778.880 451.870 779.140 452.190 ;
        RECT 1138.600 451.870 1138.860 452.190 ;
        RECT 1138.660 18.010 1138.800 451.870 ;
        RECT 1138.600 17.690 1138.860 18.010 ;
        RECT 1144.580 17.690 1144.840 18.010 ;
        RECT 1144.640 2.400 1144.780 17.690 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 786.670 496.980 786.990 497.040 ;
        RECT 792.650 496.980 792.970 497.040 ;
        RECT 786.670 496.840 792.970 496.980 ;
        RECT 786.670 496.780 786.990 496.840 ;
        RECT 792.650 496.780 792.970 496.840 ;
        RECT 792.650 445.300 792.970 445.360 ;
        RECT 1159.270 445.300 1159.590 445.360 ;
        RECT 792.650 445.160 1159.590 445.300 ;
        RECT 792.650 445.100 792.970 445.160 ;
        RECT 1159.270 445.100 1159.590 445.160 ;
      LAYER via ;
        RECT 786.700 496.780 786.960 497.040 ;
        RECT 792.680 496.780 792.940 497.040 ;
        RECT 792.680 445.100 792.940 445.360 ;
        RECT 1159.300 445.100 1159.560 445.360 ;
      LAYER met2 ;
        RECT 786.830 510.340 787.110 514.000 ;
        RECT 786.760 510.000 787.110 510.340 ;
        RECT 786.760 497.070 786.900 510.000 ;
        RECT 786.700 496.750 786.960 497.070 ;
        RECT 792.680 496.750 792.940 497.070 ;
        RECT 792.740 445.390 792.880 496.750 ;
        RECT 792.680 445.070 792.940 445.390 ;
        RECT 1159.300 445.070 1159.560 445.390 ;
        RECT 1159.360 17.410 1159.500 445.070 ;
        RECT 1159.360 17.270 1162.720 17.410 ;
        RECT 1162.580 2.400 1162.720 17.270 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 19.620 455.330 19.680 ;
        RECT 680.410 19.620 680.730 19.680 ;
        RECT 455.010 19.480 680.730 19.620 ;
        RECT 455.010 19.420 455.330 19.480 ;
        RECT 680.410 19.420 680.730 19.480 ;
      LAYER via ;
        RECT 455.040 19.420 455.300 19.680 ;
        RECT 680.440 19.420 680.700 19.680 ;
      LAYER met2 ;
        RECT 452.870 510.410 453.150 514.000 ;
        RECT 452.870 510.270 455.240 510.410 ;
        RECT 452.870 510.000 453.150 510.270 ;
        RECT 455.100 19.710 455.240 510.270 ;
        RECT 455.040 19.390 455.300 19.710 ;
        RECT 680.440 19.390 680.700 19.710 ;
        RECT 680.500 2.400 680.640 19.390 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 800.010 210.360 800.330 210.420 ;
        RECT 1179.970 210.360 1180.290 210.420 ;
        RECT 800.010 210.220 1180.290 210.360 ;
        RECT 800.010 210.160 800.330 210.220 ;
        RECT 1179.970 210.160 1180.290 210.220 ;
      LAYER via ;
        RECT 800.040 210.160 800.300 210.420 ;
        RECT 1180.000 210.160 1180.260 210.420 ;
      LAYER met2 ;
        RECT 799.250 510.410 799.530 514.000 ;
        RECT 799.250 510.270 800.240 510.410 ;
        RECT 799.250 510.000 799.530 510.270 ;
        RECT 800.100 210.450 800.240 510.270 ;
        RECT 800.040 210.130 800.300 210.450 ;
        RECT 1180.000 210.130 1180.260 210.450 ;
        RECT 1180.060 2.400 1180.200 210.130 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 813.810 190.300 814.130 190.360 ;
        RECT 1193.770 190.300 1194.090 190.360 ;
        RECT 813.810 190.160 1194.090 190.300 ;
        RECT 813.810 190.100 814.130 190.160 ;
        RECT 1193.770 190.100 1194.090 190.160 ;
      LAYER via ;
        RECT 813.840 190.100 814.100 190.360 ;
        RECT 1193.800 190.100 1194.060 190.360 ;
      LAYER met2 ;
        RECT 811.670 510.410 811.950 514.000 ;
        RECT 811.670 510.270 814.040 510.410 ;
        RECT 811.670 510.000 811.950 510.270 ;
        RECT 813.900 190.390 814.040 510.270 ;
        RECT 813.840 190.070 814.100 190.390 ;
        RECT 1193.800 190.070 1194.060 190.390 ;
        RECT 1193.860 17.410 1194.000 190.070 ;
        RECT 1193.860 17.270 1198.140 17.410 ;
        RECT 1198.000 2.400 1198.140 17.270 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 823.930 497.320 824.250 497.380 ;
        RECT 845.090 497.320 845.410 497.380 ;
        RECT 823.930 497.180 845.410 497.320 ;
        RECT 823.930 497.120 824.250 497.180 ;
        RECT 845.090 497.120 845.410 497.180 ;
        RECT 845.090 231.100 845.410 231.160 ;
        RECT 1214.470 231.100 1214.790 231.160 ;
        RECT 845.090 230.960 1214.790 231.100 ;
        RECT 845.090 230.900 845.410 230.960 ;
        RECT 1214.470 230.900 1214.790 230.960 ;
      LAYER via ;
        RECT 823.960 497.120 824.220 497.380 ;
        RECT 845.120 497.120 845.380 497.380 ;
        RECT 845.120 230.900 845.380 231.160 ;
        RECT 1214.500 230.900 1214.760 231.160 ;
      LAYER met2 ;
        RECT 824.090 510.340 824.370 514.000 ;
        RECT 824.020 510.000 824.370 510.340 ;
        RECT 824.020 497.410 824.160 510.000 ;
        RECT 823.960 497.090 824.220 497.410 ;
        RECT 845.120 497.090 845.380 497.410 ;
        RECT 845.180 231.190 845.320 497.090 ;
        RECT 845.120 230.870 845.380 231.190 ;
        RECT 1214.500 230.870 1214.760 231.190 ;
        RECT 1214.560 17.410 1214.700 230.870 ;
        RECT 1214.560 17.270 1216.080 17.410 ;
        RECT 1215.940 2.400 1216.080 17.270 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 836.350 496.980 836.670 497.040 ;
        RECT 840.950 496.980 841.270 497.040 ;
        RECT 836.350 496.840 841.270 496.980 ;
        RECT 836.350 496.780 836.670 496.840 ;
        RECT 840.950 496.780 841.270 496.840 ;
        RECT 840.950 217.500 841.270 217.560 ;
        RECT 1228.270 217.500 1228.590 217.560 ;
        RECT 840.950 217.360 1228.590 217.500 ;
        RECT 840.950 217.300 841.270 217.360 ;
        RECT 1228.270 217.300 1228.590 217.360 ;
      LAYER via ;
        RECT 836.380 496.780 836.640 497.040 ;
        RECT 840.980 496.780 841.240 497.040 ;
        RECT 840.980 217.300 841.240 217.560 ;
        RECT 1228.300 217.300 1228.560 217.560 ;
      LAYER met2 ;
        RECT 836.510 510.340 836.790 514.000 ;
        RECT 836.440 510.000 836.790 510.340 ;
        RECT 836.440 497.070 836.580 510.000 ;
        RECT 836.380 496.750 836.640 497.070 ;
        RECT 840.980 496.750 841.240 497.070 ;
        RECT 841.040 217.590 841.180 496.750 ;
        RECT 840.980 217.270 841.240 217.590 ;
        RECT 1228.300 217.270 1228.560 217.590 ;
        RECT 1228.360 17.410 1228.500 217.270 ;
        RECT 1228.360 17.270 1234.020 17.410 ;
        RECT 1233.880 2.400 1234.020 17.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.770 496.980 849.090 497.040 ;
        RECT 854.750 496.980 855.070 497.040 ;
        RECT 848.770 496.840 855.070 496.980 ;
        RECT 848.770 496.780 849.090 496.840 ;
        RECT 854.750 496.780 855.070 496.840 ;
        RECT 854.750 238.240 855.070 238.300 ;
        RECT 1248.970 238.240 1249.290 238.300 ;
        RECT 854.750 238.100 1249.290 238.240 ;
        RECT 854.750 238.040 855.070 238.100 ;
        RECT 1248.970 238.040 1249.290 238.100 ;
      LAYER via ;
        RECT 848.800 496.780 849.060 497.040 ;
        RECT 854.780 496.780 855.040 497.040 ;
        RECT 854.780 238.040 855.040 238.300 ;
        RECT 1249.000 238.040 1249.260 238.300 ;
      LAYER met2 ;
        RECT 848.930 510.340 849.210 514.000 ;
        RECT 848.860 510.000 849.210 510.340 ;
        RECT 848.860 497.070 849.000 510.000 ;
        RECT 848.800 496.750 849.060 497.070 ;
        RECT 854.780 496.750 855.040 497.070 ;
        RECT 854.840 238.330 854.980 496.750 ;
        RECT 854.780 238.010 855.040 238.330 ;
        RECT 1249.000 238.010 1249.260 238.330 ;
        RECT 1249.060 17.410 1249.200 238.010 ;
        RECT 1249.060 17.270 1251.960 17.410 ;
        RECT 1251.820 2.400 1251.960 17.270 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 990.065 476.085 990.235 500.395 ;
        RECT 990.065 427.805 990.235 475.575 ;
        RECT 990.065 379.525 990.235 401.115 ;
        RECT 990.525 96.645 990.695 144.755 ;
      LAYER mcon ;
        RECT 990.065 500.225 990.235 500.395 ;
        RECT 990.065 475.405 990.235 475.575 ;
        RECT 990.065 400.945 990.235 401.115 ;
        RECT 990.525 144.585 990.695 144.755 ;
      LAYER met1 ;
        RECT 861.190 500.380 861.510 500.440 ;
        RECT 990.005 500.380 990.295 500.425 ;
        RECT 861.190 500.240 990.295 500.380 ;
        RECT 861.190 500.180 861.510 500.240 ;
        RECT 990.005 500.195 990.295 500.240 ;
        RECT 989.990 476.240 990.310 476.300 ;
        RECT 989.795 476.100 990.310 476.240 ;
        RECT 989.990 476.040 990.310 476.100 ;
        RECT 989.990 475.560 990.310 475.620 ;
        RECT 989.795 475.420 990.310 475.560 ;
        RECT 989.990 475.360 990.310 475.420 ;
        RECT 990.005 427.960 990.295 428.005 ;
        RECT 990.450 427.960 990.770 428.020 ;
        RECT 990.005 427.820 990.770 427.960 ;
        RECT 990.005 427.775 990.295 427.820 ;
        RECT 990.450 427.760 990.770 427.820 ;
        RECT 990.005 401.100 990.295 401.145 ;
        RECT 990.450 401.100 990.770 401.160 ;
        RECT 990.005 400.960 990.770 401.100 ;
        RECT 990.005 400.915 990.295 400.960 ;
        RECT 990.450 400.900 990.770 400.960 ;
        RECT 989.990 379.680 990.310 379.740 ;
        RECT 989.795 379.540 990.310 379.680 ;
        RECT 989.990 379.480 990.310 379.540 ;
        RECT 988.610 289.920 988.930 289.980 ;
        RECT 989.990 289.920 990.310 289.980 ;
        RECT 988.610 289.780 990.310 289.920 ;
        RECT 988.610 289.720 988.930 289.780 ;
        RECT 989.990 289.720 990.310 289.780 ;
        RECT 989.990 158.680 990.310 158.740 ;
        RECT 990.910 158.680 991.230 158.740 ;
        RECT 989.990 158.540 991.230 158.680 ;
        RECT 989.990 158.480 990.310 158.540 ;
        RECT 990.910 158.480 991.230 158.540 ;
        RECT 990.465 144.740 990.755 144.785 ;
        RECT 990.910 144.740 991.230 144.800 ;
        RECT 990.465 144.600 991.230 144.740 ;
        RECT 990.465 144.555 990.755 144.600 ;
        RECT 990.910 144.540 991.230 144.600 ;
        RECT 990.450 96.800 990.770 96.860 ;
        RECT 990.255 96.660 990.770 96.800 ;
        RECT 990.450 96.600 990.770 96.660 ;
        RECT 990.910 24.380 991.230 24.440 ;
        RECT 1269.210 24.380 1269.530 24.440 ;
        RECT 990.910 24.240 1269.530 24.380 ;
        RECT 990.910 24.180 991.230 24.240 ;
        RECT 1269.210 24.180 1269.530 24.240 ;
      LAYER via ;
        RECT 861.220 500.180 861.480 500.440 ;
        RECT 990.020 476.040 990.280 476.300 ;
        RECT 990.020 475.360 990.280 475.620 ;
        RECT 990.480 427.760 990.740 428.020 ;
        RECT 990.480 400.900 990.740 401.160 ;
        RECT 990.020 379.480 990.280 379.740 ;
        RECT 988.640 289.720 988.900 289.980 ;
        RECT 990.020 289.720 990.280 289.980 ;
        RECT 990.020 158.480 990.280 158.740 ;
        RECT 990.940 158.480 991.200 158.740 ;
        RECT 990.940 144.540 991.200 144.800 ;
        RECT 990.480 96.600 990.740 96.860 ;
        RECT 990.940 24.180 991.200 24.440 ;
        RECT 1269.240 24.180 1269.500 24.440 ;
      LAYER met2 ;
        RECT 861.350 510.340 861.630 514.000 ;
        RECT 861.280 510.000 861.630 510.340 ;
        RECT 861.280 500.470 861.420 510.000 ;
        RECT 861.220 500.150 861.480 500.470 ;
        RECT 990.020 476.010 990.280 476.330 ;
        RECT 990.080 475.650 990.220 476.010 ;
        RECT 990.020 475.330 990.280 475.650 ;
        RECT 990.480 427.730 990.740 428.050 ;
        RECT 990.540 401.190 990.680 427.730 ;
        RECT 990.480 400.870 990.740 401.190 ;
        RECT 990.020 379.450 990.280 379.770 ;
        RECT 990.080 337.805 990.220 379.450 ;
        RECT 988.630 337.435 988.910 337.805 ;
        RECT 990.010 337.435 990.290 337.805 ;
        RECT 988.700 290.010 988.840 337.435 ;
        RECT 988.640 289.690 988.900 290.010 ;
        RECT 990.020 289.690 990.280 290.010 ;
        RECT 990.080 158.770 990.220 289.690 ;
        RECT 990.020 158.450 990.280 158.770 ;
        RECT 990.940 158.450 991.200 158.770 ;
        RECT 991.000 144.830 991.140 158.450 ;
        RECT 990.940 144.510 991.200 144.830 ;
        RECT 990.480 96.570 990.740 96.890 ;
        RECT 990.540 62.290 990.680 96.570 ;
        RECT 990.540 62.150 991.140 62.290 ;
        RECT 991.000 24.470 991.140 62.150 ;
        RECT 990.940 24.150 991.200 24.470 ;
        RECT 1269.240 24.150 1269.500 24.470 ;
        RECT 1269.300 2.400 1269.440 24.150 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 988.630 337.480 988.910 337.760 ;
        RECT 990.010 337.480 990.290 337.760 ;
      LAYER met3 ;
        RECT 988.605 337.770 988.935 337.785 ;
        RECT 989.985 337.770 990.315 337.785 ;
        RECT 988.605 337.470 990.315 337.770 ;
        RECT 988.605 337.455 988.935 337.470 ;
        RECT 989.985 337.455 990.315 337.470 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 875.910 410.620 876.230 410.680 ;
        RECT 1283.470 410.620 1283.790 410.680 ;
        RECT 875.910 410.480 1283.790 410.620 ;
        RECT 875.910 410.420 876.230 410.480 ;
        RECT 1283.470 410.420 1283.790 410.480 ;
      LAYER via ;
        RECT 875.940 410.420 876.200 410.680 ;
        RECT 1283.500 410.420 1283.760 410.680 ;
      LAYER met2 ;
        RECT 873.310 510.410 873.590 514.000 ;
        RECT 873.310 510.270 876.140 510.410 ;
        RECT 873.310 510.000 873.590 510.270 ;
        RECT 876.000 410.710 876.140 510.270 ;
        RECT 875.940 410.390 876.200 410.710 ;
        RECT 1283.500 410.390 1283.760 410.710 ;
        RECT 1283.560 17.410 1283.700 410.390 ;
        RECT 1283.560 17.270 1287.380 17.410 ;
        RECT 1287.240 2.400 1287.380 17.270 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 889.250 251.840 889.570 251.900 ;
        RECT 1304.170 251.840 1304.490 251.900 ;
        RECT 889.250 251.700 1304.490 251.840 ;
        RECT 889.250 251.640 889.570 251.700 ;
        RECT 1304.170 251.640 1304.490 251.700 ;
      LAYER via ;
        RECT 889.280 251.640 889.540 251.900 ;
        RECT 1304.200 251.640 1304.460 251.900 ;
      LAYER met2 ;
        RECT 885.730 510.410 886.010 514.000 ;
        RECT 885.730 510.270 889.480 510.410 ;
        RECT 885.730 510.000 886.010 510.270 ;
        RECT 889.340 251.930 889.480 510.270 ;
        RECT 889.280 251.610 889.540 251.930 ;
        RECT 1304.200 251.610 1304.460 251.930 ;
        RECT 1304.260 17.410 1304.400 251.610 ;
        RECT 1304.260 17.270 1305.320 17.410 ;
        RECT 1305.180 2.400 1305.320 17.270 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.990 496.980 898.310 497.040 ;
        RECT 903.510 496.980 903.830 497.040 ;
        RECT 897.990 496.840 903.830 496.980 ;
        RECT 897.990 496.780 898.310 496.840 ;
        RECT 903.510 496.780 903.830 496.840 ;
        RECT 903.510 258.980 903.830 259.040 ;
        RECT 1317.970 258.980 1318.290 259.040 ;
        RECT 903.510 258.840 1318.290 258.980 ;
        RECT 903.510 258.780 903.830 258.840 ;
        RECT 1317.970 258.780 1318.290 258.840 ;
        RECT 1317.970 62.120 1318.290 62.180 ;
        RECT 1323.030 62.120 1323.350 62.180 ;
        RECT 1317.970 61.980 1323.350 62.120 ;
        RECT 1317.970 61.920 1318.290 61.980 ;
        RECT 1323.030 61.920 1323.350 61.980 ;
      LAYER via ;
        RECT 898.020 496.780 898.280 497.040 ;
        RECT 903.540 496.780 903.800 497.040 ;
        RECT 903.540 258.780 903.800 259.040 ;
        RECT 1318.000 258.780 1318.260 259.040 ;
        RECT 1318.000 61.920 1318.260 62.180 ;
        RECT 1323.060 61.920 1323.320 62.180 ;
      LAYER met2 ;
        RECT 898.150 510.340 898.430 514.000 ;
        RECT 898.080 510.000 898.430 510.340 ;
        RECT 898.080 497.070 898.220 510.000 ;
        RECT 898.020 496.750 898.280 497.070 ;
        RECT 903.540 496.750 903.800 497.070 ;
        RECT 903.600 259.070 903.740 496.750 ;
        RECT 903.540 258.750 903.800 259.070 ;
        RECT 1318.000 258.750 1318.260 259.070 ;
        RECT 1318.060 62.210 1318.200 258.750 ;
        RECT 1318.000 61.890 1318.260 62.210 ;
        RECT 1323.060 61.890 1323.320 62.210 ;
        RECT 1323.120 2.400 1323.260 61.890 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1338.745 234.685 1338.915 265.795 ;
        RECT 1338.745 48.365 1338.915 113.475 ;
      LAYER mcon ;
        RECT 1338.745 265.625 1338.915 265.795 ;
        RECT 1338.745 113.305 1338.915 113.475 ;
      LAYER met1 ;
        RECT 910.410 265.780 910.730 265.840 ;
        RECT 1338.685 265.780 1338.975 265.825 ;
        RECT 910.410 265.640 1338.975 265.780 ;
        RECT 910.410 265.580 910.730 265.640 ;
        RECT 1338.685 265.595 1338.975 265.640 ;
        RECT 1338.670 234.840 1338.990 234.900 ;
        RECT 1338.475 234.700 1338.990 234.840 ;
        RECT 1338.670 234.640 1338.990 234.700 ;
        RECT 1338.670 113.460 1338.990 113.520 ;
        RECT 1338.475 113.320 1338.990 113.460 ;
        RECT 1338.670 113.260 1338.990 113.320 ;
        RECT 1338.685 48.520 1338.975 48.565 ;
        RECT 1340.510 48.520 1340.830 48.580 ;
        RECT 1338.685 48.380 1340.830 48.520 ;
        RECT 1338.685 48.335 1338.975 48.380 ;
        RECT 1340.510 48.320 1340.830 48.380 ;
      LAYER via ;
        RECT 910.440 265.580 910.700 265.840 ;
        RECT 1338.700 234.640 1338.960 234.900 ;
        RECT 1338.700 113.260 1338.960 113.520 ;
        RECT 1340.540 48.320 1340.800 48.580 ;
      LAYER met2 ;
        RECT 910.570 510.340 910.850 514.000 ;
        RECT 910.500 510.000 910.850 510.340 ;
        RECT 910.500 265.870 910.640 510.000 ;
        RECT 910.440 265.550 910.700 265.870 ;
        RECT 1338.700 234.610 1338.960 234.930 ;
        RECT 1338.760 113.550 1338.900 234.610 ;
        RECT 1338.700 113.230 1338.960 113.550 ;
        RECT 1340.540 48.290 1340.800 48.610 ;
        RECT 1340.600 2.400 1340.740 48.290 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 468.810 19.280 469.130 19.340 ;
        RECT 698.350 19.280 698.670 19.340 ;
        RECT 468.810 19.140 698.670 19.280 ;
        RECT 468.810 19.080 469.130 19.140 ;
        RECT 698.350 19.080 698.670 19.140 ;
      LAYER via ;
        RECT 468.840 19.080 469.100 19.340 ;
        RECT 698.380 19.080 698.640 19.340 ;
      LAYER met2 ;
        RECT 465.290 510.410 465.570 514.000 ;
        RECT 465.290 510.270 469.040 510.410 ;
        RECT 465.290 510.000 465.570 510.270 ;
        RECT 468.900 19.370 469.040 510.270 ;
        RECT 468.840 19.050 469.100 19.370 ;
        RECT 698.380 19.050 698.640 19.370 ;
        RECT 698.440 2.400 698.580 19.050 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 924.210 197.100 924.530 197.160 ;
        RECT 1352.930 197.100 1353.250 197.160 ;
        RECT 924.210 196.960 1353.250 197.100 ;
        RECT 924.210 196.900 924.530 196.960 ;
        RECT 1352.930 196.900 1353.250 196.960 ;
        RECT 1352.930 62.120 1353.250 62.180 ;
        RECT 1358.450 62.120 1358.770 62.180 ;
        RECT 1352.930 61.980 1358.770 62.120 ;
        RECT 1352.930 61.920 1353.250 61.980 ;
        RECT 1358.450 61.920 1358.770 61.980 ;
      LAYER via ;
        RECT 924.240 196.900 924.500 197.160 ;
        RECT 1352.960 196.900 1353.220 197.160 ;
        RECT 1352.960 61.920 1353.220 62.180 ;
        RECT 1358.480 61.920 1358.740 62.180 ;
      LAYER met2 ;
        RECT 922.990 510.410 923.270 514.000 ;
        RECT 922.990 510.270 924.440 510.410 ;
        RECT 922.990 510.000 923.270 510.270 ;
        RECT 924.300 197.190 924.440 510.270 ;
        RECT 924.240 196.870 924.500 197.190 ;
        RECT 1352.960 196.870 1353.220 197.190 ;
        RECT 1353.020 62.210 1353.160 196.870 ;
        RECT 1352.960 61.890 1353.220 62.210 ;
        RECT 1358.480 61.890 1358.740 62.210 ;
        RECT 1358.540 2.400 1358.680 61.890 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.010 438.160 938.330 438.220 ;
        RECT 1373.170 438.160 1373.490 438.220 ;
        RECT 938.010 438.020 1373.490 438.160 ;
        RECT 938.010 437.960 938.330 438.020 ;
        RECT 1373.170 437.960 1373.490 438.020 ;
      LAYER via ;
        RECT 938.040 437.960 938.300 438.220 ;
        RECT 1373.200 437.960 1373.460 438.220 ;
      LAYER met2 ;
        RECT 935.410 510.410 935.690 514.000 ;
        RECT 935.410 510.270 938.240 510.410 ;
        RECT 935.410 510.000 935.690 510.270 ;
        RECT 938.100 438.250 938.240 510.270 ;
        RECT 938.040 437.930 938.300 438.250 ;
        RECT 1373.200 437.930 1373.460 438.250 ;
        RECT 1373.260 17.410 1373.400 437.930 ;
        RECT 1373.260 17.270 1376.620 17.410 ;
        RECT 1376.480 2.400 1376.620 17.270 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 947.670 496.980 947.990 497.040 ;
        RECT 955.490 496.980 955.810 497.040 ;
        RECT 947.670 496.840 955.810 496.980 ;
        RECT 947.670 496.780 947.990 496.840 ;
        RECT 955.490 496.780 955.810 496.840 ;
        RECT 955.490 279.720 955.810 279.780 ;
        RECT 1393.870 279.720 1394.190 279.780 ;
        RECT 955.490 279.580 1394.190 279.720 ;
        RECT 955.490 279.520 955.810 279.580 ;
        RECT 1393.870 279.520 1394.190 279.580 ;
      LAYER via ;
        RECT 947.700 496.780 947.960 497.040 ;
        RECT 955.520 496.780 955.780 497.040 ;
        RECT 955.520 279.520 955.780 279.780 ;
        RECT 1393.900 279.520 1394.160 279.780 ;
      LAYER met2 ;
        RECT 947.830 510.340 948.110 514.000 ;
        RECT 947.760 510.000 948.110 510.340 ;
        RECT 947.760 497.070 947.900 510.000 ;
        RECT 947.700 496.750 947.960 497.070 ;
        RECT 955.520 496.750 955.780 497.070 ;
        RECT 955.580 279.810 955.720 496.750 ;
        RECT 955.520 279.490 955.780 279.810 ;
        RECT 1393.900 279.490 1394.160 279.810 ;
        RECT 1393.960 17.410 1394.100 279.490 ;
        RECT 1393.960 17.270 1394.560 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 960.090 496.980 960.410 497.040 ;
        RECT 965.150 496.980 965.470 497.040 ;
        RECT 960.090 496.840 965.470 496.980 ;
        RECT 960.090 496.780 960.410 496.840 ;
        RECT 965.150 496.780 965.470 496.840 ;
        RECT 965.150 286.520 965.470 286.580 ;
        RECT 1407.670 286.520 1407.990 286.580 ;
        RECT 965.150 286.380 1407.990 286.520 ;
        RECT 965.150 286.320 965.470 286.380 ;
        RECT 1407.670 286.320 1407.990 286.380 ;
      LAYER via ;
        RECT 960.120 496.780 960.380 497.040 ;
        RECT 965.180 496.780 965.440 497.040 ;
        RECT 965.180 286.320 965.440 286.580 ;
        RECT 1407.700 286.320 1407.960 286.580 ;
      LAYER met2 ;
        RECT 960.250 510.340 960.530 514.000 ;
        RECT 960.180 510.000 960.530 510.340 ;
        RECT 960.180 497.070 960.320 510.000 ;
        RECT 960.120 496.750 960.380 497.070 ;
        RECT 965.180 496.750 965.440 497.070 ;
        RECT 965.240 286.610 965.380 496.750 ;
        RECT 965.180 286.290 965.440 286.610 ;
        RECT 1407.700 286.290 1407.960 286.610 ;
        RECT 1407.760 17.410 1407.900 286.290 ;
        RECT 1407.760 17.270 1412.500 17.410 ;
        RECT 1412.360 2.400 1412.500 17.270 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 272.580 972.830 272.640 ;
        RECT 1428.370 272.580 1428.690 272.640 ;
        RECT 972.510 272.440 1428.690 272.580 ;
        RECT 972.510 272.380 972.830 272.440 ;
        RECT 1428.370 272.380 1428.690 272.440 ;
      LAYER via ;
        RECT 972.540 272.380 972.800 272.640 ;
        RECT 1428.400 272.380 1428.660 272.640 ;
      LAYER met2 ;
        RECT 972.670 510.340 972.950 514.000 ;
        RECT 972.600 510.000 972.950 510.340 ;
        RECT 972.600 272.670 972.740 510.000 ;
        RECT 972.540 272.350 972.800 272.670 ;
        RECT 1428.400 272.350 1428.660 272.670 ;
        RECT 1428.460 17.410 1428.600 272.350 ;
        RECT 1428.460 17.270 1429.980 17.410 ;
        RECT 1429.840 2.400 1429.980 17.270 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.310 245.380 986.630 245.440 ;
        RECT 1442.170 245.380 1442.490 245.440 ;
        RECT 986.310 245.240 1442.490 245.380 ;
        RECT 986.310 245.180 986.630 245.240 ;
        RECT 1442.170 245.180 1442.490 245.240 ;
      LAYER via ;
        RECT 986.340 245.180 986.600 245.440 ;
        RECT 1442.200 245.180 1442.460 245.440 ;
      LAYER met2 ;
        RECT 984.630 510.410 984.910 514.000 ;
        RECT 984.630 510.270 986.540 510.410 ;
        RECT 984.630 510.000 984.910 510.270 ;
        RECT 986.400 245.470 986.540 510.270 ;
        RECT 986.340 245.150 986.600 245.470 ;
        RECT 1442.200 245.150 1442.460 245.470 ;
        RECT 1442.260 17.410 1442.400 245.150 ;
        RECT 1442.260 17.270 1447.920 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.110 306.920 1000.430 306.980 ;
        RECT 1462.870 306.920 1463.190 306.980 ;
        RECT 1000.110 306.780 1463.190 306.920 ;
        RECT 1000.110 306.720 1000.430 306.780 ;
        RECT 1462.870 306.720 1463.190 306.780 ;
      LAYER via ;
        RECT 1000.140 306.720 1000.400 306.980 ;
        RECT 1462.900 306.720 1463.160 306.980 ;
      LAYER met2 ;
        RECT 997.050 510.410 997.330 514.000 ;
        RECT 997.050 510.270 1000.340 510.410 ;
        RECT 997.050 510.000 997.330 510.270 ;
        RECT 1000.200 307.010 1000.340 510.270 ;
        RECT 1000.140 306.690 1000.400 307.010 ;
        RECT 1462.900 306.690 1463.160 307.010 ;
        RECT 1462.960 17.410 1463.100 306.690 ;
        RECT 1462.960 17.270 1465.860 17.410 ;
        RECT 1465.720 2.400 1465.860 17.270 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1009.310 503.440 1009.630 503.500 ;
        RECT 1013.910 503.440 1014.230 503.500 ;
        RECT 1009.310 503.300 1014.230 503.440 ;
        RECT 1009.310 503.240 1009.630 503.300 ;
        RECT 1013.910 503.240 1014.230 503.300 ;
        RECT 1013.910 314.400 1014.230 314.460 ;
        RECT 1483.570 314.400 1483.890 314.460 ;
        RECT 1013.910 314.260 1483.890 314.400 ;
        RECT 1013.910 314.200 1014.230 314.260 ;
        RECT 1483.570 314.200 1483.890 314.260 ;
      LAYER via ;
        RECT 1009.340 503.240 1009.600 503.500 ;
        RECT 1013.940 503.240 1014.200 503.500 ;
        RECT 1013.940 314.200 1014.200 314.460 ;
        RECT 1483.600 314.200 1483.860 314.460 ;
      LAYER met2 ;
        RECT 1009.470 510.340 1009.750 514.000 ;
        RECT 1009.400 510.000 1009.750 510.340 ;
        RECT 1009.400 503.530 1009.540 510.000 ;
        RECT 1009.340 503.210 1009.600 503.530 ;
        RECT 1013.940 503.210 1014.200 503.530 ;
        RECT 1014.000 314.490 1014.140 503.210 ;
        RECT 1013.940 314.170 1014.200 314.490 ;
        RECT 1483.600 314.170 1483.860 314.490 ;
        RECT 1483.660 2.400 1483.800 314.170 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.730 503.440 1022.050 503.500 ;
        RECT 1027.250 503.440 1027.570 503.500 ;
        RECT 1021.730 503.300 1027.570 503.440 ;
        RECT 1021.730 503.240 1022.050 503.300 ;
        RECT 1027.250 503.240 1027.570 503.300 ;
        RECT 1027.250 321.200 1027.570 321.260 ;
        RECT 1497.370 321.200 1497.690 321.260 ;
        RECT 1027.250 321.060 1497.690 321.200 ;
        RECT 1027.250 321.000 1027.570 321.060 ;
        RECT 1497.370 321.000 1497.690 321.060 ;
      LAYER via ;
        RECT 1021.760 503.240 1022.020 503.500 ;
        RECT 1027.280 503.240 1027.540 503.500 ;
        RECT 1027.280 321.000 1027.540 321.260 ;
        RECT 1497.400 321.000 1497.660 321.260 ;
      LAYER met2 ;
        RECT 1021.890 510.340 1022.170 514.000 ;
        RECT 1021.820 510.000 1022.170 510.340 ;
        RECT 1021.820 503.530 1021.960 510.000 ;
        RECT 1021.760 503.210 1022.020 503.530 ;
        RECT 1027.280 503.210 1027.540 503.530 ;
        RECT 1027.340 321.290 1027.480 503.210 ;
        RECT 1027.280 320.970 1027.540 321.290 ;
        RECT 1497.400 320.970 1497.660 321.290 ;
        RECT 1497.460 16.730 1497.600 320.970 ;
        RECT 1497.460 16.590 1501.740 16.730 ;
        RECT 1501.600 2.400 1501.740 16.590 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 327.660 1034.930 327.720 ;
        RECT 1518.070 327.660 1518.390 327.720 ;
        RECT 1034.610 327.520 1518.390 327.660 ;
        RECT 1034.610 327.460 1034.930 327.520 ;
        RECT 1518.070 327.460 1518.390 327.520 ;
      LAYER via ;
        RECT 1034.640 327.460 1034.900 327.720 ;
        RECT 1518.100 327.460 1518.360 327.720 ;
      LAYER met2 ;
        RECT 1034.310 510.340 1034.590 514.000 ;
        RECT 1034.240 510.000 1034.590 510.340 ;
        RECT 1034.240 497.490 1034.380 510.000 ;
        RECT 1034.240 497.350 1034.840 497.490 ;
        RECT 1034.700 327.750 1034.840 497.350 ;
        RECT 1034.640 327.430 1034.900 327.750 ;
        RECT 1518.100 327.430 1518.360 327.750 ;
        RECT 1518.160 16.730 1518.300 327.430 ;
        RECT 1518.160 16.590 1519.220 16.730 ;
        RECT 1519.080 2.400 1519.220 16.590 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 477.550 498.680 477.870 498.740 ;
        RECT 482.610 498.680 482.930 498.740 ;
        RECT 477.550 498.540 482.930 498.680 ;
        RECT 477.550 498.480 477.870 498.540 ;
        RECT 482.610 498.480 482.930 498.540 ;
        RECT 482.610 18.940 482.930 19.000 ;
        RECT 716.290 18.940 716.610 19.000 ;
        RECT 482.610 18.800 716.610 18.940 ;
        RECT 482.610 18.740 482.930 18.800 ;
        RECT 716.290 18.740 716.610 18.800 ;
      LAYER via ;
        RECT 477.580 498.480 477.840 498.740 ;
        RECT 482.640 498.480 482.900 498.740 ;
        RECT 482.640 18.740 482.900 19.000 ;
        RECT 716.320 18.740 716.580 19.000 ;
      LAYER met2 ;
        RECT 477.710 510.340 477.990 514.000 ;
        RECT 477.640 510.000 477.990 510.340 ;
        RECT 477.640 498.770 477.780 510.000 ;
        RECT 477.580 498.450 477.840 498.770 ;
        RECT 482.640 498.450 482.900 498.770 ;
        RECT 482.700 19.030 482.840 498.450 ;
        RECT 482.640 18.710 482.900 19.030 ;
        RECT 716.320 18.710 716.580 19.030 ;
        RECT 716.380 2.400 716.520 18.710 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1048.410 348.740 1048.730 348.800 ;
        RECT 1531.870 348.740 1532.190 348.800 ;
        RECT 1048.410 348.600 1532.190 348.740 ;
        RECT 1048.410 348.540 1048.730 348.600 ;
        RECT 1531.870 348.540 1532.190 348.600 ;
        RECT 1531.870 2.960 1532.190 3.020 ;
        RECT 1536.930 2.960 1537.250 3.020 ;
        RECT 1531.870 2.820 1537.250 2.960 ;
        RECT 1531.870 2.760 1532.190 2.820 ;
        RECT 1536.930 2.760 1537.250 2.820 ;
      LAYER via ;
        RECT 1048.440 348.540 1048.700 348.800 ;
        RECT 1531.900 348.540 1532.160 348.800 ;
        RECT 1531.900 2.760 1532.160 3.020 ;
        RECT 1536.960 2.760 1537.220 3.020 ;
      LAYER met2 ;
        RECT 1046.730 510.410 1047.010 514.000 ;
        RECT 1046.730 510.270 1048.640 510.410 ;
        RECT 1046.730 510.000 1047.010 510.270 ;
        RECT 1048.500 348.830 1048.640 510.270 ;
        RECT 1048.440 348.510 1048.700 348.830 ;
        RECT 1531.900 348.510 1532.160 348.830 ;
        RECT 1531.960 3.050 1532.100 348.510 ;
        RECT 1531.900 2.730 1532.160 3.050 ;
        RECT 1536.960 2.730 1537.220 3.050 ;
        RECT 1537.020 2.400 1537.160 2.730 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1062.210 334.460 1062.530 334.520 ;
        RECT 1552.570 334.460 1552.890 334.520 ;
        RECT 1062.210 334.320 1552.890 334.460 ;
        RECT 1062.210 334.260 1062.530 334.320 ;
        RECT 1552.570 334.260 1552.890 334.320 ;
        RECT 1552.570 2.960 1552.890 3.020 ;
        RECT 1554.870 2.960 1555.190 3.020 ;
        RECT 1552.570 2.820 1555.190 2.960 ;
        RECT 1552.570 2.760 1552.890 2.820 ;
        RECT 1554.870 2.760 1555.190 2.820 ;
      LAYER via ;
        RECT 1062.240 334.260 1062.500 334.520 ;
        RECT 1552.600 334.260 1552.860 334.520 ;
        RECT 1552.600 2.760 1552.860 3.020 ;
        RECT 1554.900 2.760 1555.160 3.020 ;
      LAYER met2 ;
        RECT 1059.150 510.410 1059.430 514.000 ;
        RECT 1059.150 510.270 1062.440 510.410 ;
        RECT 1059.150 510.000 1059.430 510.270 ;
        RECT 1062.300 334.550 1062.440 510.270 ;
        RECT 1062.240 334.230 1062.500 334.550 ;
        RECT 1552.600 334.230 1552.860 334.550 ;
        RECT 1552.660 3.050 1552.800 334.230 ;
        RECT 1552.600 2.730 1552.860 3.050 ;
        RECT 1554.900 2.730 1555.160 3.050 ;
        RECT 1554.960 2.400 1555.100 2.730 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1071.410 496.980 1071.730 497.040 ;
        RECT 1079.690 496.980 1080.010 497.040 ;
        RECT 1071.410 496.840 1080.010 496.980 ;
        RECT 1071.410 496.780 1071.730 496.840 ;
        RECT 1079.690 496.780 1080.010 496.840 ;
        RECT 1079.690 341.600 1080.010 341.660 ;
        RECT 1566.830 341.600 1567.150 341.660 ;
        RECT 1079.690 341.460 1567.150 341.600 ;
        RECT 1079.690 341.400 1080.010 341.460 ;
        RECT 1566.830 341.400 1567.150 341.460 ;
        RECT 1566.830 17.920 1567.150 17.980 ;
        RECT 1572.810 17.920 1573.130 17.980 ;
        RECT 1566.830 17.780 1573.130 17.920 ;
        RECT 1566.830 17.720 1567.150 17.780 ;
        RECT 1572.810 17.720 1573.130 17.780 ;
      LAYER via ;
        RECT 1071.440 496.780 1071.700 497.040 ;
        RECT 1079.720 496.780 1079.980 497.040 ;
        RECT 1079.720 341.400 1079.980 341.660 ;
        RECT 1566.860 341.400 1567.120 341.660 ;
        RECT 1566.860 17.720 1567.120 17.980 ;
        RECT 1572.840 17.720 1573.100 17.980 ;
      LAYER met2 ;
        RECT 1071.570 510.340 1071.850 514.000 ;
        RECT 1071.500 510.000 1071.850 510.340 ;
        RECT 1071.500 497.070 1071.640 510.000 ;
        RECT 1071.440 496.750 1071.700 497.070 ;
        RECT 1079.720 496.750 1079.980 497.070 ;
        RECT 1079.780 341.690 1079.920 496.750 ;
        RECT 1079.720 341.370 1079.980 341.690 ;
        RECT 1566.860 341.370 1567.120 341.690 ;
        RECT 1566.920 18.010 1567.060 341.370 ;
        RECT 1566.860 17.690 1567.120 18.010 ;
        RECT 1572.840 17.690 1573.100 18.010 ;
        RECT 1572.900 2.400 1573.040 17.690 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1083.830 496.980 1084.150 497.040 ;
        RECT 1089.810 496.980 1090.130 497.040 ;
        RECT 1083.830 496.840 1090.130 496.980 ;
        RECT 1083.830 496.780 1084.150 496.840 ;
        RECT 1089.810 496.780 1090.130 496.840 ;
        RECT 1089.810 107.000 1090.130 107.060 ;
        RECT 1587.070 107.000 1587.390 107.060 ;
        RECT 1089.810 106.860 1587.390 107.000 ;
        RECT 1089.810 106.800 1090.130 106.860 ;
        RECT 1587.070 106.800 1587.390 106.860 ;
      LAYER via ;
        RECT 1083.860 496.780 1084.120 497.040 ;
        RECT 1089.840 496.780 1090.100 497.040 ;
        RECT 1089.840 106.800 1090.100 107.060 ;
        RECT 1587.100 106.800 1587.360 107.060 ;
      LAYER met2 ;
        RECT 1083.990 510.340 1084.270 514.000 ;
        RECT 1083.920 510.000 1084.270 510.340 ;
        RECT 1083.920 497.070 1084.060 510.000 ;
        RECT 1083.860 496.750 1084.120 497.070 ;
        RECT 1089.840 496.750 1090.100 497.070 ;
        RECT 1089.900 107.090 1090.040 496.750 ;
        RECT 1089.840 106.770 1090.100 107.090 ;
        RECT 1587.100 106.770 1587.360 107.090 ;
        RECT 1587.160 16.730 1587.300 106.770 ;
        RECT 1587.160 16.590 1590.520 16.730 ;
        RECT 1590.380 2.400 1590.520 16.590 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 355.200 1097.030 355.260 ;
        RECT 1607.770 355.200 1608.090 355.260 ;
        RECT 1096.710 355.060 1608.090 355.200 ;
        RECT 1096.710 355.000 1097.030 355.060 ;
        RECT 1607.770 355.000 1608.090 355.060 ;
      LAYER via ;
        RECT 1096.740 355.000 1097.000 355.260 ;
        RECT 1607.800 355.000 1608.060 355.260 ;
      LAYER met2 ;
        RECT 1095.950 510.410 1096.230 514.000 ;
        RECT 1095.950 510.270 1096.940 510.410 ;
        RECT 1095.950 510.000 1096.230 510.270 ;
        RECT 1096.800 355.290 1096.940 510.270 ;
        RECT 1096.740 354.970 1097.000 355.290 ;
        RECT 1607.800 354.970 1608.060 355.290 ;
        RECT 1607.860 17.410 1608.000 354.970 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1108.210 500.380 1108.530 500.440 ;
        RECT 1155.590 500.380 1155.910 500.440 ;
        RECT 1108.210 500.240 1155.910 500.380 ;
        RECT 1108.210 500.180 1108.530 500.240 ;
        RECT 1155.590 500.180 1155.910 500.240 ;
        RECT 1155.590 286.180 1155.910 286.240 ;
        RECT 1621.570 286.180 1621.890 286.240 ;
        RECT 1155.590 286.040 1621.890 286.180 ;
        RECT 1155.590 285.980 1155.910 286.040 ;
        RECT 1621.570 285.980 1621.890 286.040 ;
      LAYER via ;
        RECT 1108.240 500.180 1108.500 500.440 ;
        RECT 1155.620 500.180 1155.880 500.440 ;
        RECT 1155.620 285.980 1155.880 286.240 ;
        RECT 1621.600 285.980 1621.860 286.240 ;
      LAYER met2 ;
        RECT 1108.370 510.340 1108.650 514.000 ;
        RECT 1108.300 510.000 1108.650 510.340 ;
        RECT 1108.300 500.470 1108.440 510.000 ;
        RECT 1108.240 500.150 1108.500 500.470 ;
        RECT 1155.620 500.150 1155.880 500.470 ;
        RECT 1155.680 286.270 1155.820 500.150 ;
        RECT 1155.620 285.950 1155.880 286.270 ;
        RECT 1621.600 285.950 1621.860 286.270 ;
        RECT 1621.660 16.730 1621.800 285.950 ;
        RECT 1621.660 16.590 1626.400 16.730 ;
        RECT 1626.260 2.400 1626.400 16.590 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1120.630 496.980 1120.950 497.040 ;
        RECT 1124.310 496.980 1124.630 497.040 ;
        RECT 1120.630 496.840 1124.630 496.980 ;
        RECT 1120.630 496.780 1120.950 496.840 ;
        RECT 1124.310 496.780 1124.630 496.840 ;
        RECT 1124.310 362.340 1124.630 362.400 ;
        RECT 1642.270 362.340 1642.590 362.400 ;
        RECT 1124.310 362.200 1642.590 362.340 ;
        RECT 1124.310 362.140 1124.630 362.200 ;
        RECT 1642.270 362.140 1642.590 362.200 ;
      LAYER via ;
        RECT 1120.660 496.780 1120.920 497.040 ;
        RECT 1124.340 496.780 1124.600 497.040 ;
        RECT 1124.340 362.140 1124.600 362.400 ;
        RECT 1642.300 362.140 1642.560 362.400 ;
      LAYER met2 ;
        RECT 1120.790 510.340 1121.070 514.000 ;
        RECT 1120.720 510.000 1121.070 510.340 ;
        RECT 1120.720 497.070 1120.860 510.000 ;
        RECT 1120.660 496.750 1120.920 497.070 ;
        RECT 1124.340 496.750 1124.600 497.070 ;
        RECT 1124.400 362.430 1124.540 496.750 ;
        RECT 1124.340 362.110 1124.600 362.430 ;
        RECT 1642.300 362.110 1642.560 362.430 ;
        RECT 1642.360 17.410 1642.500 362.110 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1133.050 496.980 1133.370 497.040 ;
        RECT 1138.110 496.980 1138.430 497.040 ;
        RECT 1133.050 496.840 1138.430 496.980 ;
        RECT 1133.050 496.780 1133.370 496.840 ;
        RECT 1138.110 496.780 1138.430 496.840 ;
        RECT 1138.110 113.800 1138.430 113.860 ;
        RECT 1656.530 113.800 1656.850 113.860 ;
        RECT 1138.110 113.660 1656.850 113.800 ;
        RECT 1138.110 113.600 1138.430 113.660 ;
        RECT 1656.530 113.600 1656.850 113.660 ;
      LAYER via ;
        RECT 1133.080 496.780 1133.340 497.040 ;
        RECT 1138.140 496.780 1138.400 497.040 ;
        RECT 1138.140 113.600 1138.400 113.860 ;
        RECT 1656.560 113.600 1656.820 113.860 ;
      LAYER met2 ;
        RECT 1133.210 510.340 1133.490 514.000 ;
        RECT 1133.140 510.000 1133.490 510.340 ;
        RECT 1133.140 497.070 1133.280 510.000 ;
        RECT 1133.080 496.750 1133.340 497.070 ;
        RECT 1138.140 496.750 1138.400 497.070 ;
        RECT 1138.200 113.890 1138.340 496.750 ;
        RECT 1138.140 113.570 1138.400 113.890 ;
        RECT 1656.560 113.570 1656.820 113.890 ;
        RECT 1656.620 17.410 1656.760 113.570 ;
        RECT 1656.620 17.270 1662.280 17.410 ;
        RECT 1662.140 2.400 1662.280 17.270 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.470 496.980 1145.790 497.040 ;
        RECT 1151.450 496.980 1151.770 497.040 ;
        RECT 1145.470 496.840 1151.770 496.980 ;
        RECT 1145.470 496.780 1145.790 496.840 ;
        RECT 1151.450 496.780 1151.770 496.840 ;
        RECT 1151.450 279.380 1151.770 279.440 ;
        RECT 1676.770 279.380 1677.090 279.440 ;
        RECT 1151.450 279.240 1677.090 279.380 ;
        RECT 1151.450 279.180 1151.770 279.240 ;
        RECT 1676.770 279.180 1677.090 279.240 ;
      LAYER via ;
        RECT 1145.500 496.780 1145.760 497.040 ;
        RECT 1151.480 496.780 1151.740 497.040 ;
        RECT 1151.480 279.180 1151.740 279.440 ;
        RECT 1676.800 279.180 1677.060 279.440 ;
      LAYER met2 ;
        RECT 1145.630 510.340 1145.910 514.000 ;
        RECT 1145.560 510.000 1145.910 510.340 ;
        RECT 1145.560 497.070 1145.700 510.000 ;
        RECT 1145.500 496.750 1145.760 497.070 ;
        RECT 1151.480 496.750 1151.740 497.070 ;
        RECT 1151.540 279.470 1151.680 496.750 ;
        RECT 1151.480 279.150 1151.740 279.470 ;
        RECT 1676.800 279.150 1677.060 279.470 ;
        RECT 1676.860 17.410 1677.000 279.150 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.810 252.180 1159.130 252.240 ;
        RECT 1697.470 252.180 1697.790 252.240 ;
        RECT 1158.810 252.040 1697.790 252.180 ;
        RECT 1158.810 251.980 1159.130 252.040 ;
        RECT 1697.470 251.980 1697.790 252.040 ;
      LAYER via ;
        RECT 1158.840 251.980 1159.100 252.240 ;
        RECT 1697.500 251.980 1697.760 252.240 ;
      LAYER met2 ;
        RECT 1158.050 510.410 1158.330 514.000 ;
        RECT 1158.050 510.270 1159.040 510.410 ;
        RECT 1158.050 510.000 1158.330 510.270 ;
        RECT 1158.900 252.270 1159.040 510.270 ;
        RECT 1158.840 251.950 1159.100 252.270 ;
        RECT 1697.500 251.950 1697.760 252.270 ;
        RECT 1697.560 2.400 1697.700 251.950 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.970 503.440 490.290 503.500 ;
        RECT 496.410 503.440 496.730 503.500 ;
        RECT 489.970 503.300 496.730 503.440 ;
        RECT 489.970 503.240 490.290 503.300 ;
        RECT 496.410 503.240 496.730 503.300 ;
        RECT 496.410 18.600 496.730 18.660 ;
        RECT 734.230 18.600 734.550 18.660 ;
        RECT 496.410 18.460 734.550 18.600 ;
        RECT 496.410 18.400 496.730 18.460 ;
        RECT 734.230 18.400 734.550 18.460 ;
      LAYER via ;
        RECT 490.000 503.240 490.260 503.500 ;
        RECT 496.440 503.240 496.700 503.500 ;
        RECT 496.440 18.400 496.700 18.660 ;
        RECT 734.260 18.400 734.520 18.660 ;
      LAYER met2 ;
        RECT 490.130 510.340 490.410 514.000 ;
        RECT 490.060 510.000 490.410 510.340 ;
        RECT 490.060 503.530 490.200 510.000 ;
        RECT 490.000 503.210 490.260 503.530 ;
        RECT 496.440 503.210 496.700 503.530 ;
        RECT 496.500 18.690 496.640 503.210 ;
        RECT 496.440 18.370 496.700 18.690 ;
        RECT 734.260 18.370 734.520 18.690 ;
        RECT 734.320 2.400 734.460 18.370 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 120.600 1172.930 120.660 ;
        RECT 1711.270 120.600 1711.590 120.660 ;
        RECT 1172.610 120.460 1711.590 120.600 ;
        RECT 1172.610 120.400 1172.930 120.460 ;
        RECT 1711.270 120.400 1711.590 120.460 ;
      LAYER via ;
        RECT 1172.640 120.400 1172.900 120.660 ;
        RECT 1711.300 120.400 1711.560 120.660 ;
      LAYER met2 ;
        RECT 1170.470 510.410 1170.750 514.000 ;
        RECT 1170.470 510.270 1172.840 510.410 ;
        RECT 1170.470 510.000 1170.750 510.270 ;
        RECT 1172.700 120.690 1172.840 510.270 ;
        RECT 1172.640 120.370 1172.900 120.690 ;
        RECT 1711.300 120.370 1711.560 120.690 ;
        RECT 1711.360 17.410 1711.500 120.370 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 189.620 1186.730 189.680 ;
        RECT 1731.970 189.620 1732.290 189.680 ;
        RECT 1186.410 189.480 1732.290 189.620 ;
        RECT 1186.410 189.420 1186.730 189.480 ;
        RECT 1731.970 189.420 1732.290 189.480 ;
      LAYER via ;
        RECT 1186.440 189.420 1186.700 189.680 ;
        RECT 1732.000 189.420 1732.260 189.680 ;
      LAYER met2 ;
        RECT 1182.890 510.410 1183.170 514.000 ;
        RECT 1182.890 510.270 1186.640 510.410 ;
        RECT 1182.890 510.000 1183.170 510.270 ;
        RECT 1186.500 189.710 1186.640 510.270 ;
        RECT 1186.440 189.390 1186.700 189.710 ;
        RECT 1732.000 189.390 1732.260 189.710 ;
        RECT 1732.060 17.410 1732.200 189.390 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1195.150 498.680 1195.470 498.740 ;
        RECT 1200.210 498.680 1200.530 498.740 ;
        RECT 1195.150 498.540 1200.530 498.680 ;
        RECT 1195.150 498.480 1195.470 498.540 ;
        RECT 1200.210 498.480 1200.530 498.540 ;
        RECT 1200.210 37.980 1200.530 38.040 ;
        RECT 1751.290 37.980 1751.610 38.040 ;
        RECT 1200.210 37.840 1751.610 37.980 ;
        RECT 1200.210 37.780 1200.530 37.840 ;
        RECT 1751.290 37.780 1751.610 37.840 ;
      LAYER via ;
        RECT 1195.180 498.480 1195.440 498.740 ;
        RECT 1200.240 498.480 1200.500 498.740 ;
        RECT 1200.240 37.780 1200.500 38.040 ;
        RECT 1751.320 37.780 1751.580 38.040 ;
      LAYER met2 ;
        RECT 1195.310 510.340 1195.590 514.000 ;
        RECT 1195.240 510.000 1195.590 510.340 ;
        RECT 1195.240 498.770 1195.380 510.000 ;
        RECT 1195.180 498.450 1195.440 498.770 ;
        RECT 1200.240 498.450 1200.500 498.770 ;
        RECT 1200.300 38.070 1200.440 498.450 ;
        RECT 1200.240 37.750 1200.500 38.070 ;
        RECT 1751.320 37.750 1751.580 38.070 ;
        RECT 1751.380 2.400 1751.520 37.750 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.570 497.320 1207.890 497.380 ;
        RECT 1252.190 497.320 1252.510 497.380 ;
        RECT 1207.570 497.180 1252.510 497.320 ;
        RECT 1207.570 497.120 1207.890 497.180 ;
        RECT 1252.190 497.120 1252.510 497.180 ;
        RECT 1252.190 314.060 1252.510 314.120 ;
        RECT 1766.470 314.060 1766.790 314.120 ;
        RECT 1252.190 313.920 1766.790 314.060 ;
        RECT 1252.190 313.860 1252.510 313.920 ;
        RECT 1766.470 313.860 1766.790 313.920 ;
      LAYER via ;
        RECT 1207.600 497.120 1207.860 497.380 ;
        RECT 1252.220 497.120 1252.480 497.380 ;
        RECT 1252.220 313.860 1252.480 314.120 ;
        RECT 1766.500 313.860 1766.760 314.120 ;
      LAYER met2 ;
        RECT 1207.730 510.340 1208.010 514.000 ;
        RECT 1207.660 510.000 1208.010 510.340 ;
        RECT 1207.660 497.410 1207.800 510.000 ;
        RECT 1207.600 497.090 1207.860 497.410 ;
        RECT 1252.220 497.090 1252.480 497.410 ;
        RECT 1252.280 314.150 1252.420 497.090 ;
        RECT 1252.220 313.830 1252.480 314.150 ;
        RECT 1766.500 313.830 1766.760 314.150 ;
        RECT 1766.560 17.410 1766.700 313.830 ;
        RECT 1766.560 17.270 1769.000 17.410 ;
        RECT 1768.860 2.400 1769.000 17.270 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 44.780 1221.230 44.840 ;
        RECT 1786.710 44.780 1787.030 44.840 ;
        RECT 1220.910 44.640 1787.030 44.780 ;
        RECT 1220.910 44.580 1221.230 44.640 ;
        RECT 1786.710 44.580 1787.030 44.640 ;
      LAYER via ;
        RECT 1220.940 44.580 1221.200 44.840 ;
        RECT 1786.740 44.580 1787.000 44.840 ;
      LAYER met2 ;
        RECT 1219.690 510.410 1219.970 514.000 ;
        RECT 1219.690 510.270 1221.140 510.410 ;
        RECT 1219.690 510.000 1219.970 510.270 ;
        RECT 1221.000 44.870 1221.140 510.270 ;
        RECT 1220.940 44.550 1221.200 44.870 ;
        RECT 1786.740 44.550 1787.000 44.870 ;
        RECT 1786.800 2.400 1786.940 44.550 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 258.640 1235.030 258.700 ;
        RECT 1800.970 258.640 1801.290 258.700 ;
        RECT 1234.710 258.500 1801.290 258.640 ;
        RECT 1234.710 258.440 1235.030 258.500 ;
        RECT 1800.970 258.440 1801.290 258.500 ;
      LAYER via ;
        RECT 1234.740 258.440 1235.000 258.700 ;
        RECT 1801.000 258.440 1801.260 258.700 ;
      LAYER met2 ;
        RECT 1232.110 510.410 1232.390 514.000 ;
        RECT 1232.110 510.270 1234.940 510.410 ;
        RECT 1232.110 510.000 1232.390 510.270 ;
        RECT 1234.800 258.730 1234.940 510.270 ;
        RECT 1234.740 258.410 1235.000 258.730 ;
        RECT 1801.000 258.410 1801.260 258.730 ;
        RECT 1801.060 17.410 1801.200 258.410 ;
        RECT 1801.060 17.270 1804.880 17.410 ;
        RECT 1804.740 2.400 1804.880 17.270 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.050 265.440 1248.370 265.500 ;
        RECT 1821.670 265.440 1821.990 265.500 ;
        RECT 1248.050 265.300 1821.990 265.440 ;
        RECT 1248.050 265.240 1248.370 265.300 ;
        RECT 1821.670 265.240 1821.990 265.300 ;
      LAYER via ;
        RECT 1248.080 265.240 1248.340 265.500 ;
        RECT 1821.700 265.240 1821.960 265.500 ;
      LAYER met2 ;
        RECT 1244.530 510.410 1244.810 514.000 ;
        RECT 1244.530 510.270 1248.280 510.410 ;
        RECT 1244.530 510.000 1244.810 510.270 ;
        RECT 1248.140 265.530 1248.280 510.270 ;
        RECT 1248.080 265.210 1248.340 265.530 ;
        RECT 1821.700 265.210 1821.960 265.530 ;
        RECT 1821.760 17.410 1821.900 265.210 ;
        RECT 1821.760 17.270 1822.820 17.410 ;
        RECT 1822.680 2.400 1822.820 17.270 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.790 496.980 1257.110 497.040 ;
        RECT 1262.310 496.980 1262.630 497.040 ;
        RECT 1256.790 496.840 1262.630 496.980 ;
        RECT 1256.790 496.780 1257.110 496.840 ;
        RECT 1262.310 496.780 1262.630 496.840 ;
        RECT 1262.310 176.020 1262.630 176.080 ;
        RECT 1835.470 176.020 1835.790 176.080 ;
        RECT 1262.310 175.880 1835.790 176.020 ;
        RECT 1262.310 175.820 1262.630 175.880 ;
        RECT 1835.470 175.820 1835.790 175.880 ;
      LAYER via ;
        RECT 1256.820 496.780 1257.080 497.040 ;
        RECT 1262.340 496.780 1262.600 497.040 ;
        RECT 1262.340 175.820 1262.600 176.080 ;
        RECT 1835.500 175.820 1835.760 176.080 ;
      LAYER met2 ;
        RECT 1256.950 510.340 1257.230 514.000 ;
        RECT 1256.880 510.000 1257.230 510.340 ;
        RECT 1256.880 497.070 1257.020 510.000 ;
        RECT 1256.820 496.750 1257.080 497.070 ;
        RECT 1262.340 496.750 1262.600 497.070 ;
        RECT 1262.400 176.110 1262.540 496.750 ;
        RECT 1262.340 175.790 1262.600 176.110 ;
        RECT 1835.500 175.790 1835.760 176.110 ;
        RECT 1835.560 17.410 1835.700 175.790 ;
        RECT 1835.560 17.270 1840.300 17.410 ;
        RECT 1840.160 2.400 1840.300 17.270 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 320.860 1269.530 320.920 ;
        RECT 1856.170 320.860 1856.490 320.920 ;
        RECT 1269.210 320.720 1856.490 320.860 ;
        RECT 1269.210 320.660 1269.530 320.720 ;
        RECT 1856.170 320.660 1856.490 320.720 ;
      LAYER via ;
        RECT 1269.240 320.660 1269.500 320.920 ;
        RECT 1856.200 320.660 1856.460 320.920 ;
      LAYER met2 ;
        RECT 1269.370 510.340 1269.650 514.000 ;
        RECT 1269.300 510.000 1269.650 510.340 ;
        RECT 1269.300 320.950 1269.440 510.000 ;
        RECT 1269.240 320.630 1269.500 320.950 ;
        RECT 1856.200 320.630 1856.460 320.950 ;
        RECT 1856.260 17.410 1856.400 320.630 ;
        RECT 1856.260 17.270 1858.240 17.410 ;
        RECT 1858.100 2.400 1858.240 17.270 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.010 348.400 1283.330 348.460 ;
        RECT 1869.970 348.400 1870.290 348.460 ;
        RECT 1283.010 348.260 1870.290 348.400 ;
        RECT 1283.010 348.200 1283.330 348.260 ;
        RECT 1869.970 348.200 1870.290 348.260 ;
        RECT 1869.970 16.900 1870.290 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1869.970 16.760 1876.270 16.900 ;
        RECT 1869.970 16.700 1870.290 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1283.040 348.200 1283.300 348.460 ;
        RECT 1870.000 348.200 1870.260 348.460 ;
        RECT 1870.000 16.700 1870.260 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 1281.790 510.410 1282.070 514.000 ;
        RECT 1281.790 510.270 1283.240 510.410 ;
        RECT 1281.790 510.000 1282.070 510.270 ;
        RECT 1283.100 348.490 1283.240 510.270 ;
        RECT 1283.040 348.170 1283.300 348.490 ;
        RECT 1870.000 348.170 1870.260 348.490 ;
        RECT 1870.060 16.990 1870.200 348.170 ;
        RECT 1870.000 16.670 1870.260 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.310 17.920 503.630 17.980 ;
        RECT 752.170 17.920 752.490 17.980 ;
        RECT 503.310 17.780 752.490 17.920 ;
        RECT 503.310 17.720 503.630 17.780 ;
        RECT 752.170 17.720 752.490 17.780 ;
      LAYER via ;
        RECT 503.340 17.720 503.600 17.980 ;
        RECT 752.200 17.720 752.460 17.980 ;
      LAYER met2 ;
        RECT 502.550 510.410 502.830 514.000 ;
        RECT 502.550 510.270 503.540 510.410 ;
        RECT 502.550 510.000 502.830 510.270 ;
        RECT 503.400 18.010 503.540 510.270 ;
        RECT 503.340 17.690 503.600 18.010 ;
        RECT 752.200 17.690 752.460 18.010 ;
        RECT 752.260 2.400 752.400 17.690 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 58.720 1297.130 58.780 ;
        RECT 1890.670 58.720 1890.990 58.780 ;
        RECT 1296.810 58.580 1890.990 58.720 ;
        RECT 1296.810 58.520 1297.130 58.580 ;
        RECT 1890.670 58.520 1890.990 58.580 ;
      LAYER via ;
        RECT 1296.840 58.520 1297.100 58.780 ;
        RECT 1890.700 58.520 1890.960 58.780 ;
      LAYER met2 ;
        RECT 1294.210 510.410 1294.490 514.000 ;
        RECT 1294.210 510.270 1297.040 510.410 ;
        RECT 1294.210 510.000 1294.490 510.270 ;
        RECT 1296.900 58.810 1297.040 510.270 ;
        RECT 1296.840 58.490 1297.100 58.810 ;
        RECT 1890.700 58.490 1890.960 58.810 ;
        RECT 1890.760 17.410 1890.900 58.490 ;
        RECT 1890.760 17.270 1894.120 17.410 ;
        RECT 1893.980 2.400 1894.120 17.270 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.470 500.380 1306.790 500.440 ;
        RECT 1472.990 500.380 1473.310 500.440 ;
        RECT 1306.470 500.240 1473.310 500.380 ;
        RECT 1306.470 500.180 1306.790 500.240 ;
        RECT 1472.990 500.180 1473.310 500.240 ;
        RECT 1472.990 65.860 1473.310 65.920 ;
        RECT 1911.370 65.860 1911.690 65.920 ;
        RECT 1472.990 65.720 1911.690 65.860 ;
        RECT 1472.990 65.660 1473.310 65.720 ;
        RECT 1911.370 65.660 1911.690 65.720 ;
      LAYER via ;
        RECT 1306.500 500.180 1306.760 500.440 ;
        RECT 1473.020 500.180 1473.280 500.440 ;
        RECT 1473.020 65.660 1473.280 65.920 ;
        RECT 1911.400 65.660 1911.660 65.920 ;
      LAYER met2 ;
        RECT 1306.630 510.340 1306.910 514.000 ;
        RECT 1306.560 510.000 1306.910 510.340 ;
        RECT 1306.560 500.470 1306.700 510.000 ;
        RECT 1306.500 500.150 1306.760 500.470 ;
        RECT 1473.020 500.150 1473.280 500.470 ;
        RECT 1473.080 65.950 1473.220 500.150 ;
        RECT 1473.020 65.630 1473.280 65.950 ;
        RECT 1911.400 65.630 1911.660 65.950 ;
        RECT 1911.460 17.410 1911.600 65.630 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.890 503.440 1319.210 503.500 ;
        RECT 1323.950 503.440 1324.270 503.500 ;
        RECT 1318.890 503.300 1324.270 503.440 ;
        RECT 1318.890 503.240 1319.210 503.300 ;
        RECT 1323.950 503.240 1324.270 503.300 ;
        RECT 1323.950 438.500 1324.270 438.560 ;
        RECT 1925.170 438.500 1925.490 438.560 ;
        RECT 1323.950 438.360 1925.490 438.500 ;
        RECT 1323.950 438.300 1324.270 438.360 ;
        RECT 1925.170 438.300 1925.490 438.360 ;
      LAYER via ;
        RECT 1318.920 503.240 1319.180 503.500 ;
        RECT 1323.980 503.240 1324.240 503.500 ;
        RECT 1323.980 438.300 1324.240 438.560 ;
        RECT 1925.200 438.300 1925.460 438.560 ;
      LAYER met2 ;
        RECT 1319.050 510.340 1319.330 514.000 ;
        RECT 1318.980 510.000 1319.330 510.340 ;
        RECT 1318.980 503.530 1319.120 510.000 ;
        RECT 1318.920 503.210 1319.180 503.530 ;
        RECT 1323.980 503.210 1324.240 503.530 ;
        RECT 1324.040 438.590 1324.180 503.210 ;
        RECT 1323.980 438.270 1324.240 438.590 ;
        RECT 1925.200 438.270 1925.460 438.590 ;
        RECT 1925.260 17.410 1925.400 438.270 ;
        RECT 1925.260 17.270 1929.540 17.410 ;
        RECT 1929.400 2.400 1929.540 17.270 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 52.260 1331.630 52.320 ;
        RECT 1945.870 52.260 1946.190 52.320 ;
        RECT 1331.310 52.120 1946.190 52.260 ;
        RECT 1331.310 52.060 1331.630 52.120 ;
        RECT 1945.870 52.060 1946.190 52.120 ;
      LAYER via ;
        RECT 1331.340 52.060 1331.600 52.320 ;
        RECT 1945.900 52.060 1946.160 52.320 ;
      LAYER met2 ;
        RECT 1331.010 510.340 1331.290 514.000 ;
        RECT 1330.940 510.000 1331.290 510.340 ;
        RECT 1330.940 503.610 1331.080 510.000 ;
        RECT 1330.940 503.470 1331.540 503.610 ;
        RECT 1331.400 52.350 1331.540 503.470 ;
        RECT 1331.340 52.030 1331.600 52.350 ;
        RECT 1945.900 52.030 1946.160 52.350 ;
        RECT 1945.960 17.410 1946.100 52.030 ;
        RECT 1945.960 17.270 1947.480 17.410 ;
        RECT 1947.340 2.400 1947.480 17.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1344.650 328.340 1344.970 328.400 ;
        RECT 1959.670 328.340 1959.990 328.400 ;
        RECT 1344.650 328.200 1959.990 328.340 ;
        RECT 1344.650 328.140 1344.970 328.200 ;
        RECT 1959.670 328.140 1959.990 328.200 ;
      LAYER via ;
        RECT 1344.680 328.140 1344.940 328.400 ;
        RECT 1959.700 328.140 1959.960 328.400 ;
      LAYER met2 ;
        RECT 1343.430 510.410 1343.710 514.000 ;
        RECT 1343.430 510.270 1344.880 510.410 ;
        RECT 1343.430 510.000 1343.710 510.270 ;
        RECT 1344.740 328.430 1344.880 510.270 ;
        RECT 1344.680 328.110 1344.940 328.430 ;
        RECT 1959.700 328.110 1959.960 328.430 ;
        RECT 1959.760 17.410 1959.900 328.110 ;
        RECT 1959.760 17.270 1965.420 17.410 ;
        RECT 1965.280 2.400 1965.420 17.270 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.690 500.040 1356.010 500.100 ;
        RECT 1362.590 500.040 1362.910 500.100 ;
        RECT 1355.690 499.900 1362.910 500.040 ;
        RECT 1355.690 499.840 1356.010 499.900 ;
        RECT 1362.590 499.840 1362.910 499.900 ;
        RECT 1362.590 86.600 1362.910 86.660 ;
        RECT 1980.370 86.600 1980.690 86.660 ;
        RECT 1362.590 86.460 1980.690 86.600 ;
        RECT 1362.590 86.400 1362.910 86.460 ;
        RECT 1980.370 86.400 1980.690 86.460 ;
      LAYER via ;
        RECT 1355.720 499.840 1355.980 500.100 ;
        RECT 1362.620 499.840 1362.880 500.100 ;
        RECT 1362.620 86.400 1362.880 86.660 ;
        RECT 1980.400 86.400 1980.660 86.660 ;
      LAYER met2 ;
        RECT 1355.850 510.340 1356.130 514.000 ;
        RECT 1355.780 510.000 1356.130 510.340 ;
        RECT 1355.780 500.130 1355.920 510.000 ;
        RECT 1355.720 499.810 1355.980 500.130 ;
        RECT 1362.620 499.810 1362.880 500.130 ;
        RECT 1362.680 86.690 1362.820 499.810 ;
        RECT 1362.620 86.370 1362.880 86.690 ;
        RECT 1980.400 86.370 1980.660 86.690 ;
        RECT 1980.460 17.410 1980.600 86.370 ;
        RECT 1980.460 17.270 1983.360 17.410 ;
        RECT 1983.220 2.400 1983.360 17.270 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1368.110 500.040 1368.430 500.100 ;
        RECT 1417.790 500.040 1418.110 500.100 ;
        RECT 1368.110 499.900 1418.110 500.040 ;
        RECT 1368.110 499.840 1368.430 499.900 ;
        RECT 1417.790 499.840 1418.110 499.900 ;
        RECT 1417.790 93.740 1418.110 93.800 ;
        RECT 2001.530 93.740 2001.850 93.800 ;
        RECT 1417.790 93.600 2001.850 93.740 ;
        RECT 1417.790 93.540 1418.110 93.600 ;
        RECT 2001.530 93.540 2001.850 93.600 ;
      LAYER via ;
        RECT 1368.140 499.840 1368.400 500.100 ;
        RECT 1417.820 499.840 1418.080 500.100 ;
        RECT 1417.820 93.540 1418.080 93.800 ;
        RECT 2001.560 93.540 2001.820 93.800 ;
      LAYER met2 ;
        RECT 1368.270 510.340 1368.550 514.000 ;
        RECT 1368.200 510.000 1368.550 510.340 ;
        RECT 1368.200 500.130 1368.340 510.000 ;
        RECT 1368.140 499.810 1368.400 500.130 ;
        RECT 1417.820 499.810 1418.080 500.130 ;
        RECT 1417.880 93.830 1418.020 499.810 ;
        RECT 1417.820 93.510 1418.080 93.830 ;
        RECT 2001.560 93.510 2001.820 93.830 ;
        RECT 2001.620 17.410 2001.760 93.510 ;
        RECT 2001.160 17.270 2001.760 17.410 ;
        RECT 2001.160 2.400 2001.300 17.270 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.530 503.440 1380.850 503.500 ;
        RECT 1386.510 503.440 1386.830 503.500 ;
        RECT 1380.530 503.300 1386.830 503.440 ;
        RECT 1380.530 503.240 1380.850 503.300 ;
        RECT 1386.510 503.240 1386.830 503.300 ;
        RECT 1386.510 403.820 1386.830 403.880 ;
        RECT 2014.870 403.820 2015.190 403.880 ;
        RECT 1386.510 403.680 2015.190 403.820 ;
        RECT 1386.510 403.620 1386.830 403.680 ;
        RECT 2014.870 403.620 2015.190 403.680 ;
      LAYER via ;
        RECT 1380.560 503.240 1380.820 503.500 ;
        RECT 1386.540 503.240 1386.800 503.500 ;
        RECT 1386.540 403.620 1386.800 403.880 ;
        RECT 2014.900 403.620 2015.160 403.880 ;
      LAYER met2 ;
        RECT 1380.690 510.340 1380.970 514.000 ;
        RECT 1380.620 510.000 1380.970 510.340 ;
        RECT 1380.620 503.530 1380.760 510.000 ;
        RECT 1380.560 503.210 1380.820 503.530 ;
        RECT 1386.540 503.210 1386.800 503.530 ;
        RECT 1386.600 403.910 1386.740 503.210 ;
        RECT 1386.540 403.590 1386.800 403.910 ;
        RECT 2014.900 403.590 2015.160 403.910 ;
        RECT 2014.960 17.410 2015.100 403.590 ;
        RECT 2014.960 17.270 2018.780 17.410 ;
        RECT 2018.640 2.400 2018.780 17.270 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1393.025 434.945 1393.195 483.055 ;
      LAYER mcon ;
        RECT 1393.025 482.885 1393.195 483.055 ;
      LAYER met1 ;
        RECT 1392.490 483.720 1392.810 483.780 ;
        RECT 1393.410 483.720 1393.730 483.780 ;
        RECT 1392.490 483.580 1393.730 483.720 ;
        RECT 1392.490 483.520 1392.810 483.580 ;
        RECT 1393.410 483.520 1393.730 483.580 ;
        RECT 1392.965 483.040 1393.255 483.085 ;
        RECT 1393.410 483.040 1393.730 483.100 ;
        RECT 1392.965 482.900 1393.730 483.040 ;
        RECT 1392.965 482.855 1393.255 482.900 ;
        RECT 1393.410 482.840 1393.730 482.900 ;
        RECT 1392.950 435.100 1393.270 435.160 ;
        RECT 1392.755 434.960 1393.270 435.100 ;
        RECT 1392.950 434.900 1393.270 434.960 ;
        RECT 1392.950 400.220 1393.270 400.480 ;
        RECT 1393.040 399.740 1393.180 400.220 ;
        RECT 1393.410 399.740 1393.730 399.800 ;
        RECT 1393.040 399.600 1393.730 399.740 ;
        RECT 1393.410 399.540 1393.730 399.600 ;
        RECT 1392.950 335.140 1393.270 335.200 ;
        RECT 2035.570 335.140 2035.890 335.200 ;
        RECT 1392.950 335.000 2035.890 335.140 ;
        RECT 1392.950 334.940 1393.270 335.000 ;
        RECT 2035.570 334.940 2035.890 335.000 ;
      LAYER via ;
        RECT 1392.520 483.520 1392.780 483.780 ;
        RECT 1393.440 483.520 1393.700 483.780 ;
        RECT 1393.440 482.840 1393.700 483.100 ;
        RECT 1392.980 434.900 1393.240 435.160 ;
        RECT 1392.980 400.220 1393.240 400.480 ;
        RECT 1393.440 399.540 1393.700 399.800 ;
        RECT 1392.980 334.940 1393.240 335.200 ;
        RECT 2035.600 334.940 2035.860 335.200 ;
      LAYER met2 ;
        RECT 1393.110 510.410 1393.390 514.000 ;
        RECT 1392.580 510.270 1393.390 510.410 ;
        RECT 1392.580 483.810 1392.720 510.270 ;
        RECT 1393.110 510.000 1393.390 510.270 ;
        RECT 1392.520 483.490 1392.780 483.810 ;
        RECT 1393.440 483.490 1393.700 483.810 ;
        RECT 1393.500 483.130 1393.640 483.490 ;
        RECT 1393.440 482.810 1393.700 483.130 ;
        RECT 1392.980 434.870 1393.240 435.190 ;
        RECT 1393.040 400.510 1393.180 434.870 ;
        RECT 1392.980 400.190 1393.240 400.510 ;
        RECT 1393.440 399.510 1393.700 399.830 ;
        RECT 1393.500 352.650 1393.640 399.510 ;
        RECT 1393.040 352.510 1393.640 352.650 ;
        RECT 1393.040 335.230 1393.180 352.510 ;
        RECT 1392.980 334.910 1393.240 335.230 ;
        RECT 2035.600 334.910 2035.860 335.230 ;
        RECT 2035.660 17.410 2035.800 334.910 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1407.210 272.920 1407.530 272.980 ;
        RECT 2049.370 272.920 2049.690 272.980 ;
        RECT 1407.210 272.780 2049.690 272.920 ;
        RECT 1407.210 272.720 1407.530 272.780 ;
        RECT 2049.370 272.720 2049.690 272.780 ;
      LAYER via ;
        RECT 1407.240 272.720 1407.500 272.980 ;
        RECT 2049.400 272.720 2049.660 272.980 ;
      LAYER met2 ;
        RECT 1405.530 510.410 1405.810 514.000 ;
        RECT 1405.530 510.270 1407.440 510.410 ;
        RECT 1405.530 510.000 1405.810 510.270 ;
        RECT 1407.300 273.010 1407.440 510.270 ;
        RECT 1407.240 272.690 1407.500 273.010 ;
        RECT 2049.400 272.690 2049.660 273.010 ;
        RECT 2049.460 17.410 2049.600 272.690 ;
        RECT 2049.460 17.270 2054.660 17.410 ;
        RECT 2054.520 2.400 2054.660 17.270 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 18.260 517.430 18.320 ;
        RECT 769.650 18.260 769.970 18.320 ;
        RECT 517.110 18.120 769.970 18.260 ;
        RECT 517.110 18.060 517.430 18.120 ;
        RECT 769.650 18.060 769.970 18.120 ;
      LAYER via ;
        RECT 517.140 18.060 517.400 18.320 ;
        RECT 769.680 18.060 769.940 18.320 ;
      LAYER met2 ;
        RECT 514.970 510.410 515.250 514.000 ;
        RECT 514.970 510.270 517.340 510.410 ;
        RECT 514.970 510.000 515.250 510.270 ;
        RECT 517.200 18.350 517.340 510.270 ;
        RECT 517.140 18.030 517.400 18.350 ;
        RECT 769.680 18.030 769.940 18.350 ;
        RECT 769.740 2.400 769.880 18.030 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 203.560 1421.330 203.620 ;
        RECT 2070.070 203.560 2070.390 203.620 ;
        RECT 1421.010 203.420 2070.390 203.560 ;
        RECT 1421.010 203.360 1421.330 203.420 ;
        RECT 2070.070 203.360 2070.390 203.420 ;
      LAYER via ;
        RECT 1421.040 203.360 1421.300 203.620 ;
        RECT 2070.100 203.360 2070.360 203.620 ;
      LAYER met2 ;
        RECT 1417.950 510.410 1418.230 514.000 ;
        RECT 1417.950 510.270 1421.240 510.410 ;
        RECT 1417.950 510.000 1418.230 510.270 ;
        RECT 1421.100 203.650 1421.240 510.270 ;
        RECT 1421.040 203.330 1421.300 203.650 ;
        RECT 2070.100 203.330 2070.360 203.650 ;
        RECT 2070.160 17.410 2070.300 203.330 ;
        RECT 2070.160 17.270 2072.600 17.410 ;
        RECT 2072.460 2.400 2072.600 17.270 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1430.210 496.980 1430.530 497.040 ;
        RECT 1434.350 496.980 1434.670 497.040 ;
        RECT 1430.210 496.840 1434.670 496.980 ;
        RECT 1430.210 496.780 1430.530 496.840 ;
        RECT 1434.350 496.780 1434.670 496.840 ;
        RECT 1434.350 286.860 1434.670 286.920 ;
        RECT 2084.330 286.860 2084.650 286.920 ;
        RECT 1434.350 286.720 2084.650 286.860 ;
        RECT 1434.350 286.660 1434.670 286.720 ;
        RECT 2084.330 286.660 2084.650 286.720 ;
      LAYER via ;
        RECT 1430.240 496.780 1430.500 497.040 ;
        RECT 1434.380 496.780 1434.640 497.040 ;
        RECT 1434.380 286.660 1434.640 286.920 ;
        RECT 2084.360 286.660 2084.620 286.920 ;
      LAYER met2 ;
        RECT 1430.370 510.340 1430.650 514.000 ;
        RECT 1430.300 510.000 1430.650 510.340 ;
        RECT 1430.300 497.070 1430.440 510.000 ;
        RECT 1430.240 496.750 1430.500 497.070 ;
        RECT 1434.380 496.750 1434.640 497.070 ;
        RECT 1434.440 286.950 1434.580 496.750 ;
        RECT 1434.380 286.630 1434.640 286.950 ;
        RECT 2084.360 286.630 2084.620 286.950 ;
        RECT 2084.420 18.090 2084.560 286.630 ;
        RECT 2084.420 17.950 2090.080 18.090 ;
        RECT 2089.940 2.400 2090.080 17.950 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.170 496.980 1442.490 497.040 ;
        RECT 1448.610 496.980 1448.930 497.040 ;
        RECT 1442.170 496.840 1448.930 496.980 ;
        RECT 1442.170 496.780 1442.490 496.840 ;
        RECT 1448.610 496.780 1448.930 496.840 ;
        RECT 1448.610 424.560 1448.930 424.620 ;
        RECT 2104.570 424.560 2104.890 424.620 ;
        RECT 1448.610 424.420 2104.890 424.560 ;
        RECT 1448.610 424.360 1448.930 424.420 ;
        RECT 2104.570 424.360 2104.890 424.420 ;
      LAYER via ;
        RECT 1442.200 496.780 1442.460 497.040 ;
        RECT 1448.640 496.780 1448.900 497.040 ;
        RECT 1448.640 424.360 1448.900 424.620 ;
        RECT 2104.600 424.360 2104.860 424.620 ;
      LAYER met2 ;
        RECT 1442.330 510.340 1442.610 514.000 ;
        RECT 1442.260 510.000 1442.610 510.340 ;
        RECT 1442.260 497.070 1442.400 510.000 ;
        RECT 1442.200 496.750 1442.460 497.070 ;
        RECT 1448.640 496.750 1448.900 497.070 ;
        RECT 1448.700 424.650 1448.840 496.750 ;
        RECT 1448.640 424.330 1448.900 424.650 ;
        RECT 2104.600 424.330 2104.860 424.650 ;
        RECT 2104.660 17.410 2104.800 424.330 ;
        RECT 2104.660 17.270 2108.020 17.410 ;
        RECT 2107.880 2.400 2108.020 17.270 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.510 79.800 1455.830 79.860 ;
        RECT 2125.730 79.800 2126.050 79.860 ;
        RECT 1455.510 79.660 2126.050 79.800 ;
        RECT 1455.510 79.600 1455.830 79.660 ;
        RECT 2125.730 79.600 2126.050 79.660 ;
      LAYER via ;
        RECT 1455.540 79.600 1455.800 79.860 ;
        RECT 2125.760 79.600 2126.020 79.860 ;
      LAYER met2 ;
        RECT 1454.750 510.410 1455.030 514.000 ;
        RECT 1454.750 510.270 1455.740 510.410 ;
        RECT 1454.750 510.000 1455.030 510.270 ;
        RECT 1455.600 79.890 1455.740 510.270 ;
        RECT 1455.540 79.570 1455.800 79.890 ;
        RECT 2125.760 79.570 2126.020 79.890 ;
        RECT 2125.820 2.400 2125.960 79.570 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1467.010 501.060 1467.330 501.120 ;
        RECT 1548.890 501.060 1549.210 501.120 ;
        RECT 1467.010 500.920 1549.210 501.060 ;
        RECT 1467.010 500.860 1467.330 500.920 ;
        RECT 1548.890 500.860 1549.210 500.920 ;
        RECT 1548.890 432.040 1549.210 432.100 ;
        RECT 2139.070 432.040 2139.390 432.100 ;
        RECT 1548.890 431.900 2139.390 432.040 ;
        RECT 1548.890 431.840 1549.210 431.900 ;
        RECT 2139.070 431.840 2139.390 431.900 ;
      LAYER via ;
        RECT 1467.040 500.860 1467.300 501.120 ;
        RECT 1548.920 500.860 1549.180 501.120 ;
        RECT 1548.920 431.840 1549.180 432.100 ;
        RECT 2139.100 431.840 2139.360 432.100 ;
      LAYER met2 ;
        RECT 1467.170 510.340 1467.450 514.000 ;
        RECT 1467.100 510.000 1467.450 510.340 ;
        RECT 1467.100 501.150 1467.240 510.000 ;
        RECT 1467.040 500.830 1467.300 501.150 ;
        RECT 1548.920 500.830 1549.180 501.150 ;
        RECT 1548.980 432.130 1549.120 500.830 ;
        RECT 1548.920 431.810 1549.180 432.130 ;
        RECT 2139.100 431.810 2139.360 432.130 ;
        RECT 2139.160 17.410 2139.300 431.810 ;
        RECT 2139.160 17.270 2143.900 17.410 ;
        RECT 2143.760 2.400 2143.900 17.270 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1479.430 496.980 1479.750 497.040 ;
        RECT 1483.110 496.980 1483.430 497.040 ;
        RECT 1479.430 496.840 1483.430 496.980 ;
        RECT 1479.430 496.780 1479.750 496.840 ;
        RECT 1483.110 496.780 1483.430 496.840 ;
        RECT 1483.110 279.720 1483.430 279.780 ;
        RECT 2159.770 279.720 2160.090 279.780 ;
        RECT 1483.110 279.580 2160.090 279.720 ;
        RECT 1483.110 279.520 1483.430 279.580 ;
        RECT 2159.770 279.520 2160.090 279.580 ;
      LAYER via ;
        RECT 1479.460 496.780 1479.720 497.040 ;
        RECT 1483.140 496.780 1483.400 497.040 ;
        RECT 1483.140 279.520 1483.400 279.780 ;
        RECT 2159.800 279.520 2160.060 279.780 ;
      LAYER met2 ;
        RECT 1479.590 510.340 1479.870 514.000 ;
        RECT 1479.520 510.000 1479.870 510.340 ;
        RECT 1479.520 497.070 1479.660 510.000 ;
        RECT 1479.460 496.750 1479.720 497.070 ;
        RECT 1483.140 496.750 1483.400 497.070 ;
        RECT 1483.200 279.810 1483.340 496.750 ;
        RECT 1483.140 279.490 1483.400 279.810 ;
        RECT 2159.800 279.490 2160.060 279.810 ;
        RECT 2159.860 17.410 2160.000 279.490 ;
        RECT 2159.860 17.270 2161.840 17.410 ;
        RECT 2161.700 2.400 2161.840 17.270 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1491.850 496.980 1492.170 497.040 ;
        RECT 1496.450 496.980 1496.770 497.040 ;
        RECT 1491.850 496.840 1496.770 496.980 ;
        RECT 1491.850 496.780 1492.170 496.840 ;
        RECT 1496.450 496.780 1496.770 496.840 ;
        RECT 1496.450 445.300 1496.770 445.360 ;
        RECT 2173.570 445.300 2173.890 445.360 ;
        RECT 1496.450 445.160 2173.890 445.300 ;
        RECT 1496.450 445.100 1496.770 445.160 ;
        RECT 2173.570 445.100 2173.890 445.160 ;
      LAYER via ;
        RECT 1491.880 496.780 1492.140 497.040 ;
        RECT 1496.480 496.780 1496.740 497.040 ;
        RECT 1496.480 445.100 1496.740 445.360 ;
        RECT 2173.600 445.100 2173.860 445.360 ;
      LAYER met2 ;
        RECT 1492.010 510.340 1492.290 514.000 ;
        RECT 1491.940 510.000 1492.290 510.340 ;
        RECT 1491.940 497.070 1492.080 510.000 ;
        RECT 1491.880 496.750 1492.140 497.070 ;
        RECT 1496.480 496.750 1496.740 497.070 ;
        RECT 1496.540 445.390 1496.680 496.750 ;
        RECT 1496.480 445.070 1496.740 445.390 ;
        RECT 2173.600 445.070 2173.860 445.390 ;
        RECT 2173.660 17.410 2173.800 445.070 ;
        RECT 2173.660 17.270 2179.320 17.410 ;
        RECT 2179.180 2.400 2179.320 17.270 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1504.270 496.980 1504.590 497.040 ;
        RECT 1510.250 496.980 1510.570 497.040 ;
        RECT 1504.270 496.840 1510.570 496.980 ;
        RECT 1504.270 496.780 1504.590 496.840 ;
        RECT 1510.250 496.780 1510.570 496.840 ;
        RECT 1510.250 341.940 1510.570 342.000 ;
        RECT 2194.270 341.940 2194.590 342.000 ;
        RECT 1510.250 341.800 2194.590 341.940 ;
        RECT 1510.250 341.740 1510.570 341.800 ;
        RECT 2194.270 341.740 2194.590 341.800 ;
      LAYER via ;
        RECT 1504.300 496.780 1504.560 497.040 ;
        RECT 1510.280 496.780 1510.540 497.040 ;
        RECT 1510.280 341.740 1510.540 342.000 ;
        RECT 2194.300 341.740 2194.560 342.000 ;
      LAYER met2 ;
        RECT 1504.430 510.340 1504.710 514.000 ;
        RECT 1504.360 510.000 1504.710 510.340 ;
        RECT 1504.360 497.070 1504.500 510.000 ;
        RECT 1504.300 496.750 1504.560 497.070 ;
        RECT 1510.280 496.750 1510.540 497.070 ;
        RECT 1510.340 342.030 1510.480 496.750 ;
        RECT 1510.280 341.710 1510.540 342.030 ;
        RECT 2194.300 341.710 2194.560 342.030 ;
        RECT 2194.360 17.410 2194.500 341.710 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 355.540 1517.930 355.600 ;
        RECT 2214.970 355.540 2215.290 355.600 ;
        RECT 1517.610 355.400 2215.290 355.540 ;
        RECT 1517.610 355.340 1517.930 355.400 ;
        RECT 2214.970 355.340 2215.290 355.400 ;
      LAYER via ;
        RECT 1517.640 355.340 1517.900 355.600 ;
        RECT 2215.000 355.340 2215.260 355.600 ;
      LAYER met2 ;
        RECT 1516.850 510.410 1517.130 514.000 ;
        RECT 1516.850 510.270 1517.840 510.410 ;
        RECT 1516.850 510.000 1517.130 510.270 ;
        RECT 1517.700 355.630 1517.840 510.270 ;
        RECT 1517.640 355.310 1517.900 355.630 ;
        RECT 2215.000 355.310 2215.260 355.630 ;
        RECT 2215.060 2.400 2215.200 355.310 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.410 20.640 1531.730 20.700 ;
        RECT 2232.910 20.640 2233.230 20.700 ;
        RECT 1531.410 20.500 2233.230 20.640 ;
        RECT 1531.410 20.440 1531.730 20.500 ;
        RECT 2232.910 20.440 2233.230 20.500 ;
      LAYER via ;
        RECT 1531.440 20.440 1531.700 20.700 ;
        RECT 2232.940 20.440 2233.200 20.700 ;
      LAYER met2 ;
        RECT 1529.270 510.410 1529.550 514.000 ;
        RECT 1529.270 510.270 1531.640 510.410 ;
        RECT 1529.270 510.000 1529.550 510.270 ;
        RECT 1531.500 20.730 1531.640 510.270 ;
        RECT 1531.440 20.410 1531.700 20.730 ;
        RECT 2232.940 20.410 2233.200 20.730 ;
        RECT 2233.000 2.400 2233.140 20.410 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 526.770 503.440 527.090 503.500 ;
        RECT 530.910 503.440 531.230 503.500 ;
        RECT 526.770 503.300 531.230 503.440 ;
        RECT 526.770 503.240 527.090 503.300 ;
        RECT 530.910 503.240 531.230 503.300 ;
        RECT 530.910 17.580 531.230 17.640 ;
        RECT 787.590 17.580 787.910 17.640 ;
        RECT 530.910 17.440 787.910 17.580 ;
        RECT 530.910 17.380 531.230 17.440 ;
        RECT 787.590 17.380 787.910 17.440 ;
      LAYER via ;
        RECT 526.800 503.240 527.060 503.500 ;
        RECT 530.940 503.240 531.200 503.500 ;
        RECT 530.940 17.380 531.200 17.640 ;
        RECT 787.620 17.380 787.880 17.640 ;
      LAYER met2 ;
        RECT 526.930 510.340 527.210 514.000 ;
        RECT 526.860 510.000 527.210 510.340 ;
        RECT 526.860 503.530 527.000 510.000 ;
        RECT 526.800 503.210 527.060 503.530 ;
        RECT 530.940 503.210 531.200 503.530 ;
        RECT 531.000 17.670 531.140 503.210 ;
        RECT 530.940 17.350 531.200 17.670 ;
        RECT 787.620 17.350 787.880 17.670 ;
        RECT 787.680 2.400 787.820 17.350 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 20.300 1545.530 20.360 ;
        RECT 2250.850 20.300 2251.170 20.360 ;
        RECT 1545.210 20.160 2251.170 20.300 ;
        RECT 1545.210 20.100 1545.530 20.160 ;
        RECT 2250.850 20.100 2251.170 20.160 ;
      LAYER via ;
        RECT 1545.240 20.100 1545.500 20.360 ;
        RECT 2250.880 20.100 2251.140 20.360 ;
      LAYER met2 ;
        RECT 1541.690 510.410 1541.970 514.000 ;
        RECT 1541.690 510.270 1545.440 510.410 ;
        RECT 1541.690 510.000 1541.970 510.270 ;
        RECT 1545.300 20.390 1545.440 510.270 ;
        RECT 1545.240 20.070 1545.500 20.390 ;
        RECT 2250.880 20.070 2251.140 20.390 ;
        RECT 2250.940 2.400 2251.080 20.070 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1553.490 496.980 1553.810 497.040 ;
        RECT 1559.010 496.980 1559.330 497.040 ;
        RECT 1553.490 496.840 1559.330 496.980 ;
        RECT 1553.490 496.780 1553.810 496.840 ;
        RECT 1559.010 496.780 1559.330 496.840 ;
        RECT 1559.010 19.960 1559.330 20.020 ;
        RECT 2268.330 19.960 2268.650 20.020 ;
        RECT 1559.010 19.820 2268.650 19.960 ;
        RECT 1559.010 19.760 1559.330 19.820 ;
        RECT 2268.330 19.760 2268.650 19.820 ;
      LAYER via ;
        RECT 1553.520 496.780 1553.780 497.040 ;
        RECT 1559.040 496.780 1559.300 497.040 ;
        RECT 1559.040 19.760 1559.300 20.020 ;
        RECT 2268.360 19.760 2268.620 20.020 ;
      LAYER met2 ;
        RECT 1553.650 510.340 1553.930 514.000 ;
        RECT 1553.580 510.000 1553.930 510.340 ;
        RECT 1553.580 497.070 1553.720 510.000 ;
        RECT 1553.520 496.750 1553.780 497.070 ;
        RECT 1559.040 496.750 1559.300 497.070 ;
        RECT 1559.100 20.050 1559.240 496.750 ;
        RECT 1559.040 19.730 1559.300 20.050 ;
        RECT 2268.360 19.730 2268.620 20.050 ;
        RECT 2268.420 2.400 2268.560 19.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 19.280 1566.230 19.340 ;
        RECT 2286.270 19.280 2286.590 19.340 ;
        RECT 1565.910 19.140 2286.590 19.280 ;
        RECT 1565.910 19.080 1566.230 19.140 ;
        RECT 2286.270 19.080 2286.590 19.140 ;
      LAYER via ;
        RECT 1565.940 19.080 1566.200 19.340 ;
        RECT 2286.300 19.080 2286.560 19.340 ;
      LAYER met2 ;
        RECT 1566.070 510.340 1566.350 514.000 ;
        RECT 1566.000 510.000 1566.350 510.340 ;
        RECT 1566.000 19.370 1566.140 510.000 ;
        RECT 1565.940 19.050 1566.200 19.370 ;
        RECT 2286.300 19.050 2286.560 19.370 ;
        RECT 2286.360 2.400 2286.500 19.050 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 19.620 1580.030 19.680 ;
        RECT 2304.210 19.620 2304.530 19.680 ;
        RECT 1579.710 19.480 2304.530 19.620 ;
        RECT 1579.710 19.420 1580.030 19.480 ;
        RECT 2304.210 19.420 2304.530 19.480 ;
      LAYER via ;
        RECT 1579.740 19.420 1580.000 19.680 ;
        RECT 2304.240 19.420 2304.500 19.680 ;
      LAYER met2 ;
        RECT 1578.490 510.410 1578.770 514.000 ;
        RECT 1578.490 510.270 1579.940 510.410 ;
        RECT 1578.490 510.000 1578.770 510.270 ;
        RECT 1579.800 19.710 1579.940 510.270 ;
        RECT 1579.740 19.390 1580.000 19.710 ;
        RECT 2304.240 19.390 2304.500 19.710 ;
        RECT 2304.300 2.400 2304.440 19.390 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 18.940 1593.830 19.000 ;
        RECT 2322.150 18.940 2322.470 19.000 ;
        RECT 1593.510 18.800 2322.470 18.940 ;
        RECT 1593.510 18.740 1593.830 18.800 ;
        RECT 2322.150 18.740 2322.470 18.800 ;
      LAYER via ;
        RECT 1593.540 18.740 1593.800 19.000 ;
        RECT 2322.180 18.740 2322.440 19.000 ;
      LAYER met2 ;
        RECT 1590.910 510.410 1591.190 514.000 ;
        RECT 1590.910 510.270 1593.740 510.410 ;
        RECT 1590.910 510.000 1591.190 510.270 ;
        RECT 1593.600 19.030 1593.740 510.270 ;
        RECT 1593.540 18.710 1593.800 19.030 ;
        RECT 2322.180 18.710 2322.440 19.030 ;
        RECT 2322.240 2.400 2322.380 18.710 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1603.170 496.980 1603.490 497.040 ;
        RECT 1607.310 496.980 1607.630 497.040 ;
        RECT 1603.170 496.840 1607.630 496.980 ;
        RECT 1603.170 496.780 1603.490 496.840 ;
        RECT 1607.310 496.780 1607.630 496.840 ;
        RECT 1607.310 18.600 1607.630 18.660 ;
        RECT 2339.170 18.600 2339.490 18.660 ;
        RECT 1607.310 18.460 2339.490 18.600 ;
        RECT 1607.310 18.400 1607.630 18.460 ;
        RECT 2339.170 18.400 2339.490 18.460 ;
      LAYER via ;
        RECT 1603.200 496.780 1603.460 497.040 ;
        RECT 1607.340 496.780 1607.600 497.040 ;
        RECT 1607.340 18.400 1607.600 18.660 ;
        RECT 2339.200 18.400 2339.460 18.660 ;
      LAYER met2 ;
        RECT 1603.330 510.340 1603.610 514.000 ;
        RECT 1603.260 510.000 1603.610 510.340 ;
        RECT 1603.260 497.070 1603.400 510.000 ;
        RECT 1603.200 496.750 1603.460 497.070 ;
        RECT 1607.340 496.750 1607.600 497.070 ;
        RECT 1607.400 18.690 1607.540 496.750 ;
        RECT 1607.340 18.370 1607.600 18.690 ;
        RECT 2339.200 18.370 2339.460 18.690 ;
        RECT 2339.260 16.050 2339.400 18.370 ;
        RECT 2339.260 15.910 2339.860 16.050 ;
        RECT 2339.720 2.400 2339.860 15.910 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.590 496.980 1615.910 497.040 ;
        RECT 1621.110 496.980 1621.430 497.040 ;
        RECT 1615.590 496.840 1621.430 496.980 ;
        RECT 1615.590 496.780 1615.910 496.840 ;
        RECT 1621.110 496.780 1621.430 496.840 ;
        RECT 1621.110 18.260 1621.430 18.320 ;
        RECT 2357.570 18.260 2357.890 18.320 ;
        RECT 1621.110 18.120 2357.890 18.260 ;
        RECT 1621.110 18.060 1621.430 18.120 ;
        RECT 2357.570 18.060 2357.890 18.120 ;
      LAYER via ;
        RECT 1615.620 496.780 1615.880 497.040 ;
        RECT 1621.140 496.780 1621.400 497.040 ;
        RECT 1621.140 18.060 1621.400 18.320 ;
        RECT 2357.600 18.060 2357.860 18.320 ;
      LAYER met2 ;
        RECT 1615.750 510.340 1616.030 514.000 ;
        RECT 1615.680 510.000 1616.030 510.340 ;
        RECT 1615.680 497.070 1615.820 510.000 ;
        RECT 1615.620 496.750 1615.880 497.070 ;
        RECT 1621.140 496.750 1621.400 497.070 ;
        RECT 1621.200 18.350 1621.340 496.750 ;
        RECT 1621.140 18.030 1621.400 18.350 ;
        RECT 2357.600 18.030 2357.860 18.350 ;
        RECT 2357.660 2.400 2357.800 18.030 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 17.920 1628.330 17.980 ;
        RECT 2375.510 17.920 2375.830 17.980 ;
        RECT 1628.010 17.780 2375.830 17.920 ;
        RECT 1628.010 17.720 1628.330 17.780 ;
        RECT 2375.510 17.720 2375.830 17.780 ;
      LAYER via ;
        RECT 1628.040 17.720 1628.300 17.980 ;
        RECT 2375.540 17.720 2375.800 17.980 ;
      LAYER met2 ;
        RECT 1628.170 510.340 1628.450 514.000 ;
        RECT 1628.100 510.000 1628.450 510.340 ;
        RECT 1628.100 18.010 1628.240 510.000 ;
        RECT 1628.040 17.690 1628.300 18.010 ;
        RECT 2375.540 17.690 2375.800 18.010 ;
        RECT 2375.600 2.400 2375.740 17.690 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.810 17.580 1642.130 17.640 ;
        RECT 2393.450 17.580 2393.770 17.640 ;
        RECT 1641.810 17.440 2393.770 17.580 ;
        RECT 1641.810 17.380 1642.130 17.440 ;
        RECT 2393.450 17.380 2393.770 17.440 ;
      LAYER via ;
        RECT 1641.840 17.380 1642.100 17.640 ;
        RECT 2393.480 17.380 2393.740 17.640 ;
      LAYER met2 ;
        RECT 1640.590 510.410 1640.870 514.000 ;
        RECT 1640.590 510.270 1642.040 510.410 ;
        RECT 1640.590 510.000 1640.870 510.270 ;
        RECT 1641.900 17.670 1642.040 510.270 ;
        RECT 1641.840 17.350 1642.100 17.670 ;
        RECT 2393.480 17.350 2393.740 17.670 ;
        RECT 2393.540 2.400 2393.680 17.350 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.610 17.240 1655.930 17.300 ;
        RECT 2411.390 17.240 2411.710 17.300 ;
        RECT 1655.610 17.100 2411.710 17.240 ;
        RECT 1655.610 17.040 1655.930 17.100 ;
        RECT 2411.390 17.040 2411.710 17.100 ;
      LAYER via ;
        RECT 1655.640 17.040 1655.900 17.300 ;
        RECT 2411.420 17.040 2411.680 17.300 ;
      LAYER met2 ;
        RECT 1653.010 510.410 1653.290 514.000 ;
        RECT 1653.010 510.270 1655.840 510.410 ;
        RECT 1653.010 510.000 1653.290 510.270 ;
        RECT 1655.700 17.330 1655.840 510.270 ;
        RECT 1655.640 17.010 1655.900 17.330 ;
        RECT 2411.420 17.010 2411.680 17.330 ;
        RECT 2411.480 2.400 2411.620 17.010 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 539.190 503.440 539.510 503.500 ;
        RECT 544.710 503.440 545.030 503.500 ;
        RECT 539.190 503.300 545.030 503.440 ;
        RECT 539.190 503.240 539.510 503.300 ;
        RECT 544.710 503.240 545.030 503.300 ;
        RECT 544.710 17.240 545.030 17.300 ;
        RECT 805.530 17.240 805.850 17.300 ;
        RECT 544.710 17.100 805.850 17.240 ;
        RECT 544.710 17.040 545.030 17.100 ;
        RECT 805.530 17.040 805.850 17.100 ;
      LAYER via ;
        RECT 539.220 503.240 539.480 503.500 ;
        RECT 544.740 503.240 545.000 503.500 ;
        RECT 544.740 17.040 545.000 17.300 ;
        RECT 805.560 17.040 805.820 17.300 ;
      LAYER met2 ;
        RECT 539.350 510.340 539.630 514.000 ;
        RECT 539.280 510.000 539.630 510.340 ;
        RECT 539.280 503.530 539.420 510.000 ;
        RECT 539.220 503.210 539.480 503.530 ;
        RECT 544.740 503.210 545.000 503.530 ;
        RECT 544.800 17.330 544.940 503.210 ;
        RECT 544.740 17.010 545.000 17.330 ;
        RECT 805.560 17.010 805.820 17.330 ;
        RECT 805.620 2.400 805.760 17.010 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 407.170 17.580 407.490 17.640 ;
        RECT 2.830 17.440 407.490 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 407.170 17.380 407.490 17.440 ;
      LAYER via ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 407.200 17.380 407.460 17.640 ;
      LAYER met2 ;
        RECT 411.930 510.410 412.210 514.000 ;
        RECT 407.260 510.270 412.210 510.410 ;
        RECT 407.260 17.670 407.400 510.270 ;
        RECT 411.930 510.000 412.210 510.270 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 407.200 17.350 407.460 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.240 8.670 17.300 ;
        RECT 414.530 17.240 414.850 17.300 ;
        RECT 8.350 17.100 414.850 17.240 ;
        RECT 8.350 17.040 8.670 17.100 ;
        RECT 414.530 17.040 414.850 17.100 ;
      LAYER via ;
        RECT 8.380 17.040 8.640 17.300 ;
        RECT 414.560 17.040 414.820 17.300 ;
      LAYER met2 ;
        RECT 415.610 510.410 415.890 514.000 ;
        RECT 414.620 510.270 415.890 510.410 ;
        RECT 414.620 17.330 414.760 510.270 ;
        RECT 415.610 510.000 415.890 510.270 ;
        RECT 8.380 17.010 8.640 17.330 ;
        RECT 414.560 17.010 414.820 17.330 ;
        RECT 8.440 2.400 8.580 17.010 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.580 -14.220 -16.580 3533.900 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.420 7.020 3529.100 ;
        RECT 22.020 -19.020 25.020 3538.700 ;
        RECT 184.020 -9.420 187.020 3529.100 ;
        RECT 202.020 -19.020 205.020 3538.700 ;
        RECT 364.020 -9.420 367.020 3529.100 ;
        RECT 382.020 -19.020 385.020 3538.700 ;
        RECT 544.020 2112.185 547.020 3529.100 ;
        RECT 562.020 2112.185 565.020 3538.700 ;
        RECT 724.020 2112.185 727.020 3529.100 ;
        RECT 742.020 2112.185 745.020 3538.700 ;
        RECT 904.020 2112.185 907.020 3529.100 ;
        RECT 922.020 2112.185 925.020 3538.700 ;
        RECT 1084.020 2112.185 1087.020 3529.100 ;
        RECT 1102.020 2112.185 1105.020 3538.700 ;
        RECT 1264.020 2112.185 1267.020 3529.100 ;
        RECT 1282.020 2112.185 1285.020 3538.700 ;
        RECT 1444.020 2112.185 1447.020 3529.100 ;
        RECT 1462.020 2112.185 1465.020 3538.700 ;
        RECT 1624.020 2112.185 1627.020 3529.100 ;
        RECT 1642.020 2112.185 1645.020 3538.700 ;
        RECT 1804.020 2112.185 1807.020 3529.100 ;
        RECT 1822.020 2112.185 1825.020 3538.700 ;
        RECT 1984.020 2112.185 1987.020 3529.100 ;
        RECT 431.040 520.640 432.640 2101.440 ;
        RECT 544.020 -9.420 547.020 510.000 ;
        RECT 562.020 -19.020 565.020 510.000 ;
        RECT 724.020 -9.420 727.020 510.000 ;
        RECT 742.020 -19.020 745.020 510.000 ;
        RECT 904.020 -9.420 907.020 510.000 ;
        RECT 922.020 -19.020 925.020 510.000 ;
        RECT 1084.020 -9.420 1087.020 510.000 ;
        RECT 1102.020 -19.020 1105.020 510.000 ;
        RECT 1264.020 -9.420 1267.020 510.000 ;
        RECT 1282.020 -19.020 1285.020 510.000 ;
        RECT 1444.020 -9.420 1447.020 510.000 ;
        RECT 1462.020 -19.020 1465.020 510.000 ;
        RECT 1624.020 -9.420 1627.020 510.000 ;
        RECT 1642.020 -19.020 1645.020 510.000 ;
        RECT 1804.020 -9.420 1807.020 510.000 ;
        RECT 1822.020 -19.020 1825.020 510.000 ;
        RECT 1984.020 -9.420 1987.020 510.000 ;
        RECT 2002.020 -19.020 2005.020 3538.700 ;
        RECT 2164.020 -9.420 2167.020 3529.100 ;
        RECT 2182.020 -19.020 2185.020 3538.700 ;
        RECT 2344.020 -9.420 2347.020 3529.100 ;
        RECT 2362.020 -19.020 2365.020 3538.700 ;
        RECT 2524.020 -9.420 2527.020 3529.100 ;
        RECT 2542.020 -19.020 2545.020 3538.700 ;
        RECT 2704.020 -9.420 2707.020 3529.100 ;
        RECT 2722.020 -19.020 2725.020 3538.700 ;
        RECT 2884.020 -9.420 2887.020 3529.100 ;
        RECT 2902.020 -19.020 2905.020 3538.700 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.200 -14.220 2939.200 3533.900 ;
      LAYER via4 ;
        RECT -18.670 3532.610 -17.490 3533.790 ;
        RECT -18.670 3531.010 -17.490 3532.190 ;
        RECT 22.930 3532.610 24.110 3533.790 ;
        RECT 22.930 3531.010 24.110 3532.190 ;
        RECT -18.670 3449.090 -17.490 3450.270 ;
        RECT -18.670 3447.490 -17.490 3448.670 ;
        RECT -18.670 3269.090 -17.490 3270.270 ;
        RECT -18.670 3267.490 -17.490 3268.670 ;
        RECT -18.670 3089.090 -17.490 3090.270 ;
        RECT -18.670 3087.490 -17.490 3088.670 ;
        RECT -18.670 2909.090 -17.490 2910.270 ;
        RECT -18.670 2907.490 -17.490 2908.670 ;
        RECT -18.670 2729.090 -17.490 2730.270 ;
        RECT -18.670 2727.490 -17.490 2728.670 ;
        RECT -18.670 2549.090 -17.490 2550.270 ;
        RECT -18.670 2547.490 -17.490 2548.670 ;
        RECT -18.670 2369.090 -17.490 2370.270 ;
        RECT -18.670 2367.490 -17.490 2368.670 ;
        RECT -18.670 2189.090 -17.490 2190.270 ;
        RECT -18.670 2187.490 -17.490 2188.670 ;
        RECT -18.670 2009.090 -17.490 2010.270 ;
        RECT -18.670 2007.490 -17.490 2008.670 ;
        RECT -18.670 1829.090 -17.490 1830.270 ;
        RECT -18.670 1827.490 -17.490 1828.670 ;
        RECT -18.670 1649.090 -17.490 1650.270 ;
        RECT -18.670 1647.490 -17.490 1648.670 ;
        RECT -18.670 1469.090 -17.490 1470.270 ;
        RECT -18.670 1467.490 -17.490 1468.670 ;
        RECT -18.670 1289.090 -17.490 1290.270 ;
        RECT -18.670 1287.490 -17.490 1288.670 ;
        RECT -18.670 1109.090 -17.490 1110.270 ;
        RECT -18.670 1107.490 -17.490 1108.670 ;
        RECT -18.670 929.090 -17.490 930.270 ;
        RECT -18.670 927.490 -17.490 928.670 ;
        RECT -18.670 749.090 -17.490 750.270 ;
        RECT -18.670 747.490 -17.490 748.670 ;
        RECT -18.670 569.090 -17.490 570.270 ;
        RECT -18.670 567.490 -17.490 568.670 ;
        RECT -18.670 389.090 -17.490 390.270 ;
        RECT -18.670 387.490 -17.490 388.670 ;
        RECT -18.670 209.090 -17.490 210.270 ;
        RECT -18.670 207.490 -17.490 208.670 ;
        RECT -18.670 29.090 -17.490 30.270 ;
        RECT -18.670 27.490 -17.490 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 202.930 3532.610 204.110 3533.790 ;
        RECT 202.930 3531.010 204.110 3532.190 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.670 -12.510 -17.490 -11.330 ;
        RECT -18.670 -14.110 -17.490 -12.930 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 382.930 3532.610 384.110 3533.790 ;
        RECT 382.930 3531.010 384.110 3532.190 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 22.930 -12.510 24.110 -11.330 ;
        RECT 22.930 -14.110 24.110 -12.930 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 562.930 3532.610 564.110 3533.790 ;
        RECT 562.930 3531.010 564.110 3532.190 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 742.930 3532.610 744.110 3533.790 ;
        RECT 742.930 3531.010 744.110 3532.190 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 922.930 3532.610 924.110 3533.790 ;
        RECT 922.930 3531.010 924.110 3532.190 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 1102.930 3532.610 1104.110 3533.790 ;
        RECT 1102.930 3531.010 1104.110 3532.190 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1282.930 3532.610 1284.110 3533.790 ;
        RECT 1282.930 3531.010 1284.110 3532.190 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1462.930 3532.610 1464.110 3533.790 ;
        RECT 1462.930 3531.010 1464.110 3532.190 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1642.930 3532.610 1644.110 3533.790 ;
        RECT 1642.930 3531.010 1644.110 3532.190 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1822.930 3532.610 1824.110 3533.790 ;
        RECT 1822.930 3531.010 1824.110 3532.190 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 2002.930 3532.610 2004.110 3533.790 ;
        RECT 2002.930 3531.010 2004.110 3532.190 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 2182.930 3532.610 2184.110 3533.790 ;
        RECT 2182.930 3531.010 2184.110 3532.190 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 431.250 2009.090 432.430 2010.270 ;
        RECT 431.250 2007.490 432.430 2008.670 ;
        RECT 431.250 1991.090 432.430 1992.270 ;
        RECT 431.250 1989.490 432.430 1990.670 ;
        RECT 431.250 1829.090 432.430 1830.270 ;
        RECT 431.250 1827.490 432.430 1828.670 ;
        RECT 431.250 1811.090 432.430 1812.270 ;
        RECT 431.250 1809.490 432.430 1810.670 ;
        RECT 431.250 1649.090 432.430 1650.270 ;
        RECT 431.250 1647.490 432.430 1648.670 ;
        RECT 431.250 1631.090 432.430 1632.270 ;
        RECT 431.250 1629.490 432.430 1630.670 ;
        RECT 431.250 1469.090 432.430 1470.270 ;
        RECT 431.250 1467.490 432.430 1468.670 ;
        RECT 431.250 1451.090 432.430 1452.270 ;
        RECT 431.250 1449.490 432.430 1450.670 ;
        RECT 431.250 1289.090 432.430 1290.270 ;
        RECT 431.250 1287.490 432.430 1288.670 ;
        RECT 431.250 1271.090 432.430 1272.270 ;
        RECT 431.250 1269.490 432.430 1270.670 ;
        RECT 431.250 1109.090 432.430 1110.270 ;
        RECT 431.250 1107.490 432.430 1108.670 ;
        RECT 431.250 1091.090 432.430 1092.270 ;
        RECT 431.250 1089.490 432.430 1090.670 ;
        RECT 431.250 929.090 432.430 930.270 ;
        RECT 431.250 927.490 432.430 928.670 ;
        RECT 431.250 911.090 432.430 912.270 ;
        RECT 431.250 909.490 432.430 910.670 ;
        RECT 431.250 749.090 432.430 750.270 ;
        RECT 431.250 747.490 432.430 748.670 ;
        RECT 431.250 731.090 432.430 732.270 ;
        RECT 431.250 729.490 432.430 730.670 ;
        RECT 431.250 569.090 432.430 570.270 ;
        RECT 431.250 567.490 432.430 568.670 ;
        RECT 431.250 551.090 432.430 552.270 ;
        RECT 431.250 549.490 432.430 550.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 202.930 -12.510 204.110 -11.330 ;
        RECT 202.930 -14.110 204.110 -12.930 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 382.930 -12.510 384.110 -11.330 ;
        RECT 382.930 -14.110 384.110 -12.930 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 562.930 -12.510 564.110 -11.330 ;
        RECT 562.930 -14.110 564.110 -12.930 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 742.930 -12.510 744.110 -11.330 ;
        RECT 742.930 -14.110 744.110 -12.930 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 922.930 -12.510 924.110 -11.330 ;
        RECT 922.930 -14.110 924.110 -12.930 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1102.930 -12.510 1104.110 -11.330 ;
        RECT 1102.930 -14.110 1104.110 -12.930 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1282.930 -12.510 1284.110 -11.330 ;
        RECT 1282.930 -14.110 1284.110 -12.930 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1462.930 -12.510 1464.110 -11.330 ;
        RECT 1462.930 -14.110 1464.110 -12.930 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1642.930 -12.510 1644.110 -11.330 ;
        RECT 1642.930 -14.110 1644.110 -12.930 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 1822.930 -12.510 1824.110 -11.330 ;
        RECT 1822.930 -14.110 1824.110 -12.930 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2362.930 3532.610 2364.110 3533.790 ;
        RECT 2362.930 3531.010 2364.110 3532.190 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2002.930 -12.510 2004.110 -11.330 ;
        RECT 2002.930 -14.110 2004.110 -12.930 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2542.930 3532.610 2544.110 3533.790 ;
        RECT 2542.930 3531.010 2544.110 3532.190 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2182.930 -12.510 2184.110 -11.330 ;
        RECT 2182.930 -14.110 2184.110 -12.930 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2722.930 3532.610 2724.110 3533.790 ;
        RECT 2722.930 3531.010 2724.110 3532.190 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2362.930 -12.510 2364.110 -11.330 ;
        RECT 2362.930 -14.110 2364.110 -12.930 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2902.930 3532.610 2904.110 3533.790 ;
        RECT 2902.930 3531.010 2904.110 3532.190 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2542.930 -12.510 2544.110 -11.330 ;
        RECT 2542.930 -14.110 2544.110 -12.930 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2937.110 3532.610 2938.290 3533.790 ;
        RECT 2937.110 3531.010 2938.290 3532.190 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2722.930 -12.510 2724.110 -11.330 ;
        RECT 2722.930 -14.110 2724.110 -12.930 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2937.110 3449.090 2938.290 3450.270 ;
        RECT 2937.110 3447.490 2938.290 3448.670 ;
        RECT 2937.110 3269.090 2938.290 3270.270 ;
        RECT 2937.110 3267.490 2938.290 3268.670 ;
        RECT 2937.110 3089.090 2938.290 3090.270 ;
        RECT 2937.110 3087.490 2938.290 3088.670 ;
        RECT 2937.110 2909.090 2938.290 2910.270 ;
        RECT 2937.110 2907.490 2938.290 2908.670 ;
        RECT 2937.110 2729.090 2938.290 2730.270 ;
        RECT 2937.110 2727.490 2938.290 2728.670 ;
        RECT 2937.110 2549.090 2938.290 2550.270 ;
        RECT 2937.110 2547.490 2938.290 2548.670 ;
        RECT 2937.110 2369.090 2938.290 2370.270 ;
        RECT 2937.110 2367.490 2938.290 2368.670 ;
        RECT 2937.110 2189.090 2938.290 2190.270 ;
        RECT 2937.110 2187.490 2938.290 2188.670 ;
        RECT 2937.110 2009.090 2938.290 2010.270 ;
        RECT 2937.110 2007.490 2938.290 2008.670 ;
        RECT 2937.110 1829.090 2938.290 1830.270 ;
        RECT 2937.110 1827.490 2938.290 1828.670 ;
        RECT 2937.110 1649.090 2938.290 1650.270 ;
        RECT 2937.110 1647.490 2938.290 1648.670 ;
        RECT 2937.110 1469.090 2938.290 1470.270 ;
        RECT 2937.110 1467.490 2938.290 1468.670 ;
        RECT 2937.110 1289.090 2938.290 1290.270 ;
        RECT 2937.110 1287.490 2938.290 1288.670 ;
        RECT 2937.110 1109.090 2938.290 1110.270 ;
        RECT 2937.110 1107.490 2938.290 1108.670 ;
        RECT 2937.110 929.090 2938.290 930.270 ;
        RECT 2937.110 927.490 2938.290 928.670 ;
        RECT 2937.110 749.090 2938.290 750.270 ;
        RECT 2937.110 747.490 2938.290 748.670 ;
        RECT 2937.110 569.090 2938.290 570.270 ;
        RECT 2937.110 567.490 2938.290 568.670 ;
        RECT 2937.110 389.090 2938.290 390.270 ;
        RECT 2937.110 387.490 2938.290 388.670 ;
        RECT 2937.110 209.090 2938.290 210.270 ;
        RECT 2937.110 207.490 2938.290 208.670 ;
        RECT 2937.110 29.090 2938.290 30.270 ;
        RECT 2937.110 27.490 2938.290 28.670 ;
        RECT 2902.930 -12.510 2904.110 -11.330 ;
        RECT 2902.930 -14.110 2904.110 -12.930 ;
        RECT 2937.110 -12.510 2938.290 -11.330 ;
        RECT 2937.110 -14.110 2938.290 -12.930 ;
      LAYER met5 ;
        RECT -19.580 3533.900 -16.580 3533.910 ;
        RECT 22.020 3533.900 25.020 3533.910 ;
        RECT 202.020 3533.900 205.020 3533.910 ;
        RECT 382.020 3533.900 385.020 3533.910 ;
        RECT 562.020 3533.900 565.020 3533.910 ;
        RECT 742.020 3533.900 745.020 3533.910 ;
        RECT 922.020 3533.900 925.020 3533.910 ;
        RECT 1102.020 3533.900 1105.020 3533.910 ;
        RECT 1282.020 3533.900 1285.020 3533.910 ;
        RECT 1462.020 3533.900 1465.020 3533.910 ;
        RECT 1642.020 3533.900 1645.020 3533.910 ;
        RECT 1822.020 3533.900 1825.020 3533.910 ;
        RECT 2002.020 3533.900 2005.020 3533.910 ;
        RECT 2182.020 3533.900 2185.020 3533.910 ;
        RECT 2362.020 3533.900 2365.020 3533.910 ;
        RECT 2542.020 3533.900 2545.020 3533.910 ;
        RECT 2722.020 3533.900 2725.020 3533.910 ;
        RECT 2902.020 3533.900 2905.020 3533.910 ;
        RECT 2936.200 3533.900 2939.200 3533.910 ;
        RECT -19.580 3530.900 2939.200 3533.900 ;
        RECT -19.580 3530.890 -16.580 3530.900 ;
        RECT 22.020 3530.890 25.020 3530.900 ;
        RECT 202.020 3530.890 205.020 3530.900 ;
        RECT 382.020 3530.890 385.020 3530.900 ;
        RECT 562.020 3530.890 565.020 3530.900 ;
        RECT 742.020 3530.890 745.020 3530.900 ;
        RECT 922.020 3530.890 925.020 3530.900 ;
        RECT 1102.020 3530.890 1105.020 3530.900 ;
        RECT 1282.020 3530.890 1285.020 3530.900 ;
        RECT 1462.020 3530.890 1465.020 3530.900 ;
        RECT 1642.020 3530.890 1645.020 3530.900 ;
        RECT 1822.020 3530.890 1825.020 3530.900 ;
        RECT 2002.020 3530.890 2005.020 3530.900 ;
        RECT 2182.020 3530.890 2185.020 3530.900 ;
        RECT 2362.020 3530.890 2365.020 3530.900 ;
        RECT 2542.020 3530.890 2545.020 3530.900 ;
        RECT 2722.020 3530.890 2725.020 3530.900 ;
        RECT 2902.020 3530.890 2905.020 3530.900 ;
        RECT 2936.200 3530.890 2939.200 3530.900 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -19.580 3450.380 -16.580 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.200 3450.380 2939.200 3450.390 ;
        RECT -24.380 3447.380 2944.000 3450.380 ;
        RECT -19.580 3447.370 -16.580 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.200 3447.370 2939.200 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.780 3429.380 2934.400 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -19.580 3270.380 -16.580 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.200 3270.380 2939.200 3270.390 ;
        RECT -24.380 3267.380 2944.000 3270.380 ;
        RECT -19.580 3267.370 -16.580 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.200 3267.370 2939.200 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.780 3249.380 2934.400 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -19.580 3090.380 -16.580 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.200 3090.380 2939.200 3090.390 ;
        RECT -24.380 3087.380 2944.000 3090.380 ;
        RECT -19.580 3087.370 -16.580 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.200 3087.370 2939.200 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.780 3069.380 2934.400 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -19.580 2910.380 -16.580 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.200 2910.380 2939.200 2910.390 ;
        RECT -24.380 2907.380 2944.000 2910.380 ;
        RECT -19.580 2907.370 -16.580 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.200 2907.370 2939.200 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.780 2889.380 2934.400 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -19.580 2730.380 -16.580 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.200 2730.380 2939.200 2730.390 ;
        RECT -24.380 2727.380 2944.000 2730.380 ;
        RECT -19.580 2727.370 -16.580 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.200 2727.370 2939.200 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.780 2709.380 2934.400 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -19.580 2550.380 -16.580 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.200 2550.380 2939.200 2550.390 ;
        RECT -24.380 2547.380 2944.000 2550.380 ;
        RECT -19.580 2547.370 -16.580 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.200 2547.370 2939.200 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.780 2529.380 2934.400 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -19.580 2370.380 -16.580 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.200 2370.380 2939.200 2370.390 ;
        RECT -24.380 2367.380 2944.000 2370.380 ;
        RECT -19.580 2367.370 -16.580 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.200 2367.370 2939.200 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.780 2349.380 2934.400 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -19.580 2190.380 -16.580 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.200 2190.380 2939.200 2190.390 ;
        RECT -24.380 2187.380 2944.000 2190.380 ;
        RECT -19.580 2187.370 -16.580 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.200 2187.370 2939.200 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.780 2169.380 2934.400 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -19.580 2010.380 -16.580 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 431.040 2010.380 432.640 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.200 2010.380 2939.200 2010.390 ;
        RECT -24.380 2007.380 2944.000 2010.380 ;
        RECT -19.580 2007.370 -16.580 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 431.040 2007.370 432.640 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.200 2007.370 2939.200 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 431.040 1992.380 432.640 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.780 1989.380 2934.400 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 431.040 1989.370 432.640 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -19.580 1830.380 -16.580 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 431.040 1830.380 432.640 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.200 1830.380 2939.200 1830.390 ;
        RECT -24.380 1827.380 2944.000 1830.380 ;
        RECT -19.580 1827.370 -16.580 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 431.040 1827.370 432.640 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.200 1827.370 2939.200 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 431.040 1812.380 432.640 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.780 1809.380 2934.400 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 431.040 1809.370 432.640 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -19.580 1650.380 -16.580 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 431.040 1650.380 432.640 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.200 1650.380 2939.200 1650.390 ;
        RECT -24.380 1647.380 2944.000 1650.380 ;
        RECT -19.580 1647.370 -16.580 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 431.040 1647.370 432.640 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.200 1647.370 2939.200 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 431.040 1632.380 432.640 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.780 1629.380 2934.400 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 431.040 1629.370 432.640 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -19.580 1470.380 -16.580 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 431.040 1470.380 432.640 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.200 1470.380 2939.200 1470.390 ;
        RECT -24.380 1467.380 2944.000 1470.380 ;
        RECT -19.580 1467.370 -16.580 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 431.040 1467.370 432.640 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.200 1467.370 2939.200 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 431.040 1452.380 432.640 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.780 1449.380 2934.400 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 431.040 1449.370 432.640 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -19.580 1290.380 -16.580 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 431.040 1290.380 432.640 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.200 1290.380 2939.200 1290.390 ;
        RECT -24.380 1287.380 2944.000 1290.380 ;
        RECT -19.580 1287.370 -16.580 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 431.040 1287.370 432.640 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.200 1287.370 2939.200 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 431.040 1272.380 432.640 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.780 1269.380 2934.400 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 431.040 1269.370 432.640 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -19.580 1110.380 -16.580 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 431.040 1110.380 432.640 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.200 1110.380 2939.200 1110.390 ;
        RECT -24.380 1107.380 2944.000 1110.380 ;
        RECT -19.580 1107.370 -16.580 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 431.040 1107.370 432.640 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.200 1107.370 2939.200 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 431.040 1092.380 432.640 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.780 1089.380 2934.400 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 431.040 1089.370 432.640 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -19.580 930.380 -16.580 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 431.040 930.380 432.640 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.200 930.380 2939.200 930.390 ;
        RECT -24.380 927.380 2944.000 930.380 ;
        RECT -19.580 927.370 -16.580 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 431.040 927.370 432.640 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.200 927.370 2939.200 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 431.040 912.380 432.640 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.780 909.380 2934.400 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 431.040 909.370 432.640 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -19.580 750.380 -16.580 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 431.040 750.380 432.640 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.200 750.380 2939.200 750.390 ;
        RECT -24.380 747.380 2944.000 750.380 ;
        RECT -19.580 747.370 -16.580 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 431.040 747.370 432.640 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.200 747.370 2939.200 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 431.040 732.380 432.640 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.780 729.380 2934.400 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 431.040 729.370 432.640 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -19.580 570.380 -16.580 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 431.040 570.380 432.640 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.200 570.380 2939.200 570.390 ;
        RECT -24.380 567.380 2944.000 570.380 ;
        RECT -19.580 567.370 -16.580 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 431.040 567.370 432.640 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.200 567.370 2939.200 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 431.040 552.380 432.640 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.780 549.380 2934.400 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 431.040 549.370 432.640 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -19.580 390.380 -16.580 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.200 390.380 2939.200 390.390 ;
        RECT -24.380 387.380 2944.000 390.380 ;
        RECT -19.580 387.370 -16.580 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.200 387.370 2939.200 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.780 369.380 2934.400 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -19.580 210.380 -16.580 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.200 210.380 2939.200 210.390 ;
        RECT -24.380 207.380 2944.000 210.380 ;
        RECT -19.580 207.370 -16.580 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.200 207.370 2939.200 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.780 189.380 2934.400 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -19.580 30.380 -16.580 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.200 30.380 2939.200 30.390 ;
        RECT -24.380 27.380 2944.000 30.380 ;
        RECT -19.580 27.370 -16.580 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.200 27.370 2939.200 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.780 9.380 2934.400 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.580 -11.220 -16.580 -11.210 ;
        RECT 22.020 -11.220 25.020 -11.210 ;
        RECT 202.020 -11.220 205.020 -11.210 ;
        RECT 382.020 -11.220 385.020 -11.210 ;
        RECT 562.020 -11.220 565.020 -11.210 ;
        RECT 742.020 -11.220 745.020 -11.210 ;
        RECT 922.020 -11.220 925.020 -11.210 ;
        RECT 1102.020 -11.220 1105.020 -11.210 ;
        RECT 1282.020 -11.220 1285.020 -11.210 ;
        RECT 1462.020 -11.220 1465.020 -11.210 ;
        RECT 1642.020 -11.220 1645.020 -11.210 ;
        RECT 1822.020 -11.220 1825.020 -11.210 ;
        RECT 2002.020 -11.220 2005.020 -11.210 ;
        RECT 2182.020 -11.220 2185.020 -11.210 ;
        RECT 2362.020 -11.220 2365.020 -11.210 ;
        RECT 2542.020 -11.220 2545.020 -11.210 ;
        RECT 2722.020 -11.220 2725.020 -11.210 ;
        RECT 2902.020 -11.220 2905.020 -11.210 ;
        RECT 2936.200 -11.220 2939.200 -11.210 ;
        RECT -19.580 -14.220 2939.200 -11.220 ;
        RECT -19.580 -14.230 -16.580 -14.220 ;
        RECT 22.020 -14.230 25.020 -14.220 ;
        RECT 202.020 -14.230 205.020 -14.220 ;
        RECT 382.020 -14.230 385.020 -14.220 ;
        RECT 562.020 -14.230 565.020 -14.220 ;
        RECT 742.020 -14.230 745.020 -14.220 ;
        RECT 922.020 -14.230 925.020 -14.220 ;
        RECT 1102.020 -14.230 1105.020 -14.220 ;
        RECT 1282.020 -14.230 1285.020 -14.220 ;
        RECT 1462.020 -14.230 1465.020 -14.220 ;
        RECT 1642.020 -14.230 1645.020 -14.220 ;
        RECT 1822.020 -14.230 1825.020 -14.220 ;
        RECT 2002.020 -14.230 2005.020 -14.220 ;
        RECT 2182.020 -14.230 2185.020 -14.220 ;
        RECT 2362.020 -14.230 2365.020 -14.220 ;
        RECT 2542.020 -14.230 2545.020 -14.220 ;
        RECT 2722.020 -14.230 2725.020 -14.220 ;
        RECT 2902.020 -14.230 2905.020 -14.220 ;
        RECT 2936.200 -14.230 2939.200 -14.220 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.380 -19.020 -21.380 3538.700 ;
        RECT -14.780 -9.420 -11.780 3529.100 ;
        RECT 94.020 -9.420 97.020 3529.100 ;
        RECT 112.020 -19.020 115.020 3538.700 ;
        RECT 274.020 -9.420 277.020 3529.100 ;
        RECT 292.020 -19.020 295.020 3538.700 ;
        RECT 454.020 2112.185 457.020 3529.100 ;
        RECT 472.020 2112.185 475.020 3538.700 ;
        RECT 634.020 2112.185 637.020 3529.100 ;
        RECT 652.020 2112.185 655.020 3538.700 ;
        RECT 814.020 2112.185 817.020 3529.100 ;
        RECT 832.020 2112.185 835.020 3538.700 ;
        RECT 994.020 2112.185 997.020 3529.100 ;
        RECT 1012.020 2112.185 1015.020 3538.700 ;
        RECT 1174.020 2112.185 1177.020 3529.100 ;
        RECT 1192.020 2112.185 1195.020 3538.700 ;
        RECT 1354.020 2112.185 1357.020 3529.100 ;
        RECT 1372.020 2112.185 1375.020 3538.700 ;
        RECT 1534.020 2112.185 1537.020 3529.100 ;
        RECT 1552.020 2112.185 1555.020 3538.700 ;
        RECT 1714.020 2112.185 1717.020 3529.100 ;
        RECT 1732.020 2112.185 1735.020 3538.700 ;
        RECT 1894.020 2112.185 1897.020 3529.100 ;
        RECT 1912.020 2112.185 1915.020 3538.700 ;
        RECT 507.840 520.640 509.440 2101.440 ;
        RECT 454.020 -9.420 457.020 510.000 ;
        RECT 472.020 -19.020 475.020 510.000 ;
        RECT 634.020 -9.420 637.020 510.000 ;
        RECT 652.020 -19.020 655.020 510.000 ;
        RECT 814.020 -9.420 817.020 510.000 ;
        RECT 832.020 -19.020 835.020 510.000 ;
        RECT 994.020 -9.420 997.020 510.000 ;
        RECT 1012.020 -19.020 1015.020 510.000 ;
        RECT 1174.020 -9.420 1177.020 510.000 ;
        RECT 1192.020 -19.020 1195.020 510.000 ;
        RECT 1354.020 -9.420 1357.020 510.000 ;
        RECT 1372.020 -19.020 1375.020 510.000 ;
        RECT 1534.020 -9.420 1537.020 510.000 ;
        RECT 1552.020 -19.020 1555.020 510.000 ;
        RECT 1714.020 -9.420 1717.020 510.000 ;
        RECT 1732.020 -19.020 1735.020 510.000 ;
        RECT 1894.020 -9.420 1897.020 510.000 ;
        RECT 1912.020 -19.020 1915.020 510.000 ;
        RECT 2074.020 -9.420 2077.020 3529.100 ;
        RECT 2092.020 -19.020 2095.020 3538.700 ;
        RECT 2254.020 -9.420 2257.020 3529.100 ;
        RECT 2272.020 -19.020 2275.020 3538.700 ;
        RECT 2434.020 -9.420 2437.020 3529.100 ;
        RECT 2452.020 -19.020 2455.020 3538.700 ;
        RECT 2614.020 -9.420 2617.020 3529.100 ;
        RECT 2632.020 -19.020 2635.020 3538.700 ;
        RECT 2794.020 -9.420 2797.020 3529.100 ;
        RECT 2812.020 -19.020 2815.020 3538.700 ;
        RECT 2931.400 -9.420 2934.400 3529.100 ;
        RECT 2941.000 -19.020 2944.000 3538.700 ;
      LAYER via4 ;
        RECT -23.470 3537.410 -22.290 3538.590 ;
        RECT -23.470 3535.810 -22.290 3536.990 ;
        RECT 112.930 3537.410 114.110 3538.590 ;
        RECT 112.930 3535.810 114.110 3536.990 ;
        RECT -23.470 3359.090 -22.290 3360.270 ;
        RECT -23.470 3357.490 -22.290 3358.670 ;
        RECT -23.470 3179.090 -22.290 3180.270 ;
        RECT -23.470 3177.490 -22.290 3178.670 ;
        RECT -23.470 2999.090 -22.290 3000.270 ;
        RECT -23.470 2997.490 -22.290 2998.670 ;
        RECT -23.470 2819.090 -22.290 2820.270 ;
        RECT -23.470 2817.490 -22.290 2818.670 ;
        RECT -23.470 2639.090 -22.290 2640.270 ;
        RECT -23.470 2637.490 -22.290 2638.670 ;
        RECT -23.470 2459.090 -22.290 2460.270 ;
        RECT -23.470 2457.490 -22.290 2458.670 ;
        RECT -23.470 2279.090 -22.290 2280.270 ;
        RECT -23.470 2277.490 -22.290 2278.670 ;
        RECT -23.470 2099.090 -22.290 2100.270 ;
        RECT -23.470 2097.490 -22.290 2098.670 ;
        RECT -23.470 1919.090 -22.290 1920.270 ;
        RECT -23.470 1917.490 -22.290 1918.670 ;
        RECT -23.470 1739.090 -22.290 1740.270 ;
        RECT -23.470 1737.490 -22.290 1738.670 ;
        RECT -23.470 1559.090 -22.290 1560.270 ;
        RECT -23.470 1557.490 -22.290 1558.670 ;
        RECT -23.470 1379.090 -22.290 1380.270 ;
        RECT -23.470 1377.490 -22.290 1378.670 ;
        RECT -23.470 1199.090 -22.290 1200.270 ;
        RECT -23.470 1197.490 -22.290 1198.670 ;
        RECT -23.470 1019.090 -22.290 1020.270 ;
        RECT -23.470 1017.490 -22.290 1018.670 ;
        RECT -23.470 839.090 -22.290 840.270 ;
        RECT -23.470 837.490 -22.290 838.670 ;
        RECT -23.470 659.090 -22.290 660.270 ;
        RECT -23.470 657.490 -22.290 658.670 ;
        RECT -23.470 479.090 -22.290 480.270 ;
        RECT -23.470 477.490 -22.290 478.670 ;
        RECT -23.470 299.090 -22.290 300.270 ;
        RECT -23.470 297.490 -22.290 298.670 ;
        RECT -23.470 119.090 -22.290 120.270 ;
        RECT -23.470 117.490 -22.290 118.670 ;
        RECT -13.870 3527.810 -12.690 3528.990 ;
        RECT -13.870 3526.210 -12.690 3527.390 ;
        RECT -13.870 3341.090 -12.690 3342.270 ;
        RECT -13.870 3339.490 -12.690 3340.670 ;
        RECT -13.870 3161.090 -12.690 3162.270 ;
        RECT -13.870 3159.490 -12.690 3160.670 ;
        RECT -13.870 2981.090 -12.690 2982.270 ;
        RECT -13.870 2979.490 -12.690 2980.670 ;
        RECT -13.870 2801.090 -12.690 2802.270 ;
        RECT -13.870 2799.490 -12.690 2800.670 ;
        RECT -13.870 2621.090 -12.690 2622.270 ;
        RECT -13.870 2619.490 -12.690 2620.670 ;
        RECT -13.870 2441.090 -12.690 2442.270 ;
        RECT -13.870 2439.490 -12.690 2440.670 ;
        RECT -13.870 2261.090 -12.690 2262.270 ;
        RECT -13.870 2259.490 -12.690 2260.670 ;
        RECT -13.870 2081.090 -12.690 2082.270 ;
        RECT -13.870 2079.490 -12.690 2080.670 ;
        RECT -13.870 1901.090 -12.690 1902.270 ;
        RECT -13.870 1899.490 -12.690 1900.670 ;
        RECT -13.870 1721.090 -12.690 1722.270 ;
        RECT -13.870 1719.490 -12.690 1720.670 ;
        RECT -13.870 1541.090 -12.690 1542.270 ;
        RECT -13.870 1539.490 -12.690 1540.670 ;
        RECT -13.870 1361.090 -12.690 1362.270 ;
        RECT -13.870 1359.490 -12.690 1360.670 ;
        RECT -13.870 1181.090 -12.690 1182.270 ;
        RECT -13.870 1179.490 -12.690 1180.670 ;
        RECT -13.870 1001.090 -12.690 1002.270 ;
        RECT -13.870 999.490 -12.690 1000.670 ;
        RECT -13.870 821.090 -12.690 822.270 ;
        RECT -13.870 819.490 -12.690 820.670 ;
        RECT -13.870 641.090 -12.690 642.270 ;
        RECT -13.870 639.490 -12.690 640.670 ;
        RECT -13.870 461.090 -12.690 462.270 ;
        RECT -13.870 459.490 -12.690 460.670 ;
        RECT -13.870 281.090 -12.690 282.270 ;
        RECT -13.870 279.490 -12.690 280.670 ;
        RECT -13.870 101.090 -12.690 102.270 ;
        RECT -13.870 99.490 -12.690 100.670 ;
        RECT -13.870 -7.710 -12.690 -6.530 ;
        RECT -13.870 -9.310 -12.690 -8.130 ;
        RECT 94.930 3527.810 96.110 3528.990 ;
        RECT 94.930 3526.210 96.110 3527.390 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.710 96.110 -6.530 ;
        RECT 94.930 -9.310 96.110 -8.130 ;
        RECT 292.930 3537.410 294.110 3538.590 ;
        RECT 292.930 3535.810 294.110 3536.990 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.470 -17.310 -22.290 -16.130 ;
        RECT -23.470 -18.910 -22.290 -17.730 ;
        RECT 274.930 3527.810 276.110 3528.990 ;
        RECT 274.930 3526.210 276.110 3527.390 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.710 276.110 -6.530 ;
        RECT 274.930 -9.310 276.110 -8.130 ;
        RECT 472.930 3537.410 474.110 3538.590 ;
        RECT 472.930 3535.810 474.110 3536.990 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 454.930 3527.810 456.110 3528.990 ;
        RECT 454.930 3526.210 456.110 3527.390 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 652.930 3537.410 654.110 3538.590 ;
        RECT 652.930 3535.810 654.110 3536.990 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 634.930 3527.810 636.110 3528.990 ;
        RECT 634.930 3526.210 636.110 3527.390 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 832.930 3537.410 834.110 3538.590 ;
        RECT 832.930 3535.810 834.110 3536.990 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 814.930 3527.810 816.110 3528.990 ;
        RECT 814.930 3526.210 816.110 3527.390 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 1012.930 3537.410 1014.110 3538.590 ;
        RECT 1012.930 3535.810 1014.110 3536.990 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 994.930 3527.810 996.110 3528.990 ;
        RECT 994.930 3526.210 996.110 3527.390 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 1192.930 3537.410 1194.110 3538.590 ;
        RECT 1192.930 3535.810 1194.110 3536.990 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1174.930 3527.810 1176.110 3528.990 ;
        RECT 1174.930 3526.210 1176.110 3527.390 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1372.930 3537.410 1374.110 3538.590 ;
        RECT 1372.930 3535.810 1374.110 3536.990 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1354.930 3527.810 1356.110 3528.990 ;
        RECT 1354.930 3526.210 1356.110 3527.390 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1552.930 3537.410 1554.110 3538.590 ;
        RECT 1552.930 3535.810 1554.110 3536.990 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1534.930 3527.810 1536.110 3528.990 ;
        RECT 1534.930 3526.210 1536.110 3527.390 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1732.930 3537.410 1734.110 3538.590 ;
        RECT 1732.930 3535.810 1734.110 3536.990 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1714.930 3527.810 1716.110 3528.990 ;
        RECT 1714.930 3526.210 1716.110 3527.390 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1912.930 3537.410 1914.110 3538.590 ;
        RECT 1912.930 3535.810 1914.110 3536.990 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1894.930 3527.810 1896.110 3528.990 ;
        RECT 1894.930 3526.210 1896.110 3527.390 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 2092.930 3537.410 2094.110 3538.590 ;
        RECT 2092.930 3535.810 2094.110 3536.990 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 2074.930 3527.810 2076.110 3528.990 ;
        RECT 2074.930 3526.210 2076.110 3527.390 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 508.050 2099.090 509.230 2100.270 ;
        RECT 508.050 2097.490 509.230 2098.670 ;
        RECT 508.050 2081.090 509.230 2082.270 ;
        RECT 508.050 2079.490 509.230 2080.670 ;
        RECT 508.050 1919.090 509.230 1920.270 ;
        RECT 508.050 1917.490 509.230 1918.670 ;
        RECT 508.050 1901.090 509.230 1902.270 ;
        RECT 508.050 1899.490 509.230 1900.670 ;
        RECT 508.050 1739.090 509.230 1740.270 ;
        RECT 508.050 1737.490 509.230 1738.670 ;
        RECT 508.050 1721.090 509.230 1722.270 ;
        RECT 508.050 1719.490 509.230 1720.670 ;
        RECT 508.050 1559.090 509.230 1560.270 ;
        RECT 508.050 1557.490 509.230 1558.670 ;
        RECT 508.050 1541.090 509.230 1542.270 ;
        RECT 508.050 1539.490 509.230 1540.670 ;
        RECT 508.050 1379.090 509.230 1380.270 ;
        RECT 508.050 1377.490 509.230 1378.670 ;
        RECT 508.050 1361.090 509.230 1362.270 ;
        RECT 508.050 1359.490 509.230 1360.670 ;
        RECT 508.050 1199.090 509.230 1200.270 ;
        RECT 508.050 1197.490 509.230 1198.670 ;
        RECT 508.050 1181.090 509.230 1182.270 ;
        RECT 508.050 1179.490 509.230 1180.670 ;
        RECT 508.050 1019.090 509.230 1020.270 ;
        RECT 508.050 1017.490 509.230 1018.670 ;
        RECT 508.050 1001.090 509.230 1002.270 ;
        RECT 508.050 999.490 509.230 1000.670 ;
        RECT 508.050 839.090 509.230 840.270 ;
        RECT 508.050 837.490 509.230 838.670 ;
        RECT 508.050 821.090 509.230 822.270 ;
        RECT 508.050 819.490 509.230 820.670 ;
        RECT 508.050 659.090 509.230 660.270 ;
        RECT 508.050 657.490 509.230 658.670 ;
        RECT 508.050 641.090 509.230 642.270 ;
        RECT 508.050 639.490 509.230 640.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 112.930 -17.310 114.110 -16.130 ;
        RECT 112.930 -18.910 114.110 -17.730 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.710 456.110 -6.530 ;
        RECT 454.930 -9.310 456.110 -8.130 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 292.930 -17.310 294.110 -16.130 ;
        RECT 292.930 -18.910 294.110 -17.730 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.710 636.110 -6.530 ;
        RECT 634.930 -9.310 636.110 -8.130 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 472.930 -17.310 474.110 -16.130 ;
        RECT 472.930 -18.910 474.110 -17.730 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.710 816.110 -6.530 ;
        RECT 814.930 -9.310 816.110 -8.130 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 652.930 -17.310 654.110 -16.130 ;
        RECT 652.930 -18.910 654.110 -17.730 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.710 996.110 -6.530 ;
        RECT 994.930 -9.310 996.110 -8.130 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 832.930 -17.310 834.110 -16.130 ;
        RECT 832.930 -18.910 834.110 -17.730 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.710 1176.110 -6.530 ;
        RECT 1174.930 -9.310 1176.110 -8.130 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1012.930 -17.310 1014.110 -16.130 ;
        RECT 1012.930 -18.910 1014.110 -17.730 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.710 1356.110 -6.530 ;
        RECT 1354.930 -9.310 1356.110 -8.130 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1192.930 -17.310 1194.110 -16.130 ;
        RECT 1192.930 -18.910 1194.110 -17.730 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.710 1536.110 -6.530 ;
        RECT 1534.930 -9.310 1536.110 -8.130 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1372.930 -17.310 1374.110 -16.130 ;
        RECT 1372.930 -18.910 1374.110 -17.730 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.710 1716.110 -6.530 ;
        RECT 1714.930 -9.310 1716.110 -8.130 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1552.930 -17.310 1554.110 -16.130 ;
        RECT 1552.930 -18.910 1554.110 -17.730 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.710 1896.110 -6.530 ;
        RECT 1894.930 -9.310 1896.110 -8.130 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1732.930 -17.310 1734.110 -16.130 ;
        RECT 1732.930 -18.910 1734.110 -17.730 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.710 2076.110 -6.530 ;
        RECT 2074.930 -9.310 2076.110 -8.130 ;
        RECT 2272.930 3537.410 2274.110 3538.590 ;
        RECT 2272.930 3535.810 2274.110 3536.990 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 1912.930 -17.310 1914.110 -16.130 ;
        RECT 1912.930 -18.910 1914.110 -17.730 ;
        RECT 2254.930 3527.810 2256.110 3528.990 ;
        RECT 2254.930 3526.210 2256.110 3527.390 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.710 2256.110 -6.530 ;
        RECT 2254.930 -9.310 2256.110 -8.130 ;
        RECT 2452.930 3537.410 2454.110 3538.590 ;
        RECT 2452.930 3535.810 2454.110 3536.990 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2092.930 -17.310 2094.110 -16.130 ;
        RECT 2092.930 -18.910 2094.110 -17.730 ;
        RECT 2434.930 3527.810 2436.110 3528.990 ;
        RECT 2434.930 3526.210 2436.110 3527.390 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.710 2436.110 -6.530 ;
        RECT 2434.930 -9.310 2436.110 -8.130 ;
        RECT 2632.930 3537.410 2634.110 3538.590 ;
        RECT 2632.930 3535.810 2634.110 3536.990 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2272.930 -17.310 2274.110 -16.130 ;
        RECT 2272.930 -18.910 2274.110 -17.730 ;
        RECT 2614.930 3527.810 2616.110 3528.990 ;
        RECT 2614.930 3526.210 2616.110 3527.390 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.710 2616.110 -6.530 ;
        RECT 2614.930 -9.310 2616.110 -8.130 ;
        RECT 2812.930 3537.410 2814.110 3538.590 ;
        RECT 2812.930 3535.810 2814.110 3536.990 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2452.930 -17.310 2454.110 -16.130 ;
        RECT 2452.930 -18.910 2454.110 -17.730 ;
        RECT 2794.930 3527.810 2796.110 3528.990 ;
        RECT 2794.930 3526.210 2796.110 3527.390 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.710 2796.110 -6.530 ;
        RECT 2794.930 -9.310 2796.110 -8.130 ;
        RECT 2941.910 3537.410 2943.090 3538.590 ;
        RECT 2941.910 3535.810 2943.090 3536.990 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2632.930 -17.310 2634.110 -16.130 ;
        RECT 2632.930 -18.910 2634.110 -17.730 ;
        RECT 2932.310 3527.810 2933.490 3528.990 ;
        RECT 2932.310 3526.210 2933.490 3527.390 ;
        RECT 2932.310 3341.090 2933.490 3342.270 ;
        RECT 2932.310 3339.490 2933.490 3340.670 ;
        RECT 2932.310 3161.090 2933.490 3162.270 ;
        RECT 2932.310 3159.490 2933.490 3160.670 ;
        RECT 2932.310 2981.090 2933.490 2982.270 ;
        RECT 2932.310 2979.490 2933.490 2980.670 ;
        RECT 2932.310 2801.090 2933.490 2802.270 ;
        RECT 2932.310 2799.490 2933.490 2800.670 ;
        RECT 2932.310 2621.090 2933.490 2622.270 ;
        RECT 2932.310 2619.490 2933.490 2620.670 ;
        RECT 2932.310 2441.090 2933.490 2442.270 ;
        RECT 2932.310 2439.490 2933.490 2440.670 ;
        RECT 2932.310 2261.090 2933.490 2262.270 ;
        RECT 2932.310 2259.490 2933.490 2260.670 ;
        RECT 2932.310 2081.090 2933.490 2082.270 ;
        RECT 2932.310 2079.490 2933.490 2080.670 ;
        RECT 2932.310 1901.090 2933.490 1902.270 ;
        RECT 2932.310 1899.490 2933.490 1900.670 ;
        RECT 2932.310 1721.090 2933.490 1722.270 ;
        RECT 2932.310 1719.490 2933.490 1720.670 ;
        RECT 2932.310 1541.090 2933.490 1542.270 ;
        RECT 2932.310 1539.490 2933.490 1540.670 ;
        RECT 2932.310 1361.090 2933.490 1362.270 ;
        RECT 2932.310 1359.490 2933.490 1360.670 ;
        RECT 2932.310 1181.090 2933.490 1182.270 ;
        RECT 2932.310 1179.490 2933.490 1180.670 ;
        RECT 2932.310 1001.090 2933.490 1002.270 ;
        RECT 2932.310 999.490 2933.490 1000.670 ;
        RECT 2932.310 821.090 2933.490 822.270 ;
        RECT 2932.310 819.490 2933.490 820.670 ;
        RECT 2932.310 641.090 2933.490 642.270 ;
        RECT 2932.310 639.490 2933.490 640.670 ;
        RECT 2932.310 461.090 2933.490 462.270 ;
        RECT 2932.310 459.490 2933.490 460.670 ;
        RECT 2932.310 281.090 2933.490 282.270 ;
        RECT 2932.310 279.490 2933.490 280.670 ;
        RECT 2932.310 101.090 2933.490 102.270 ;
        RECT 2932.310 99.490 2933.490 100.670 ;
        RECT 2932.310 -7.710 2933.490 -6.530 ;
        RECT 2932.310 -9.310 2933.490 -8.130 ;
        RECT 2941.910 3359.090 2943.090 3360.270 ;
        RECT 2941.910 3357.490 2943.090 3358.670 ;
        RECT 2941.910 3179.090 2943.090 3180.270 ;
        RECT 2941.910 3177.490 2943.090 3178.670 ;
        RECT 2941.910 2999.090 2943.090 3000.270 ;
        RECT 2941.910 2997.490 2943.090 2998.670 ;
        RECT 2941.910 2819.090 2943.090 2820.270 ;
        RECT 2941.910 2817.490 2943.090 2818.670 ;
        RECT 2941.910 2639.090 2943.090 2640.270 ;
        RECT 2941.910 2637.490 2943.090 2638.670 ;
        RECT 2941.910 2459.090 2943.090 2460.270 ;
        RECT 2941.910 2457.490 2943.090 2458.670 ;
        RECT 2941.910 2279.090 2943.090 2280.270 ;
        RECT 2941.910 2277.490 2943.090 2278.670 ;
        RECT 2941.910 2099.090 2943.090 2100.270 ;
        RECT 2941.910 2097.490 2943.090 2098.670 ;
        RECT 2941.910 1919.090 2943.090 1920.270 ;
        RECT 2941.910 1917.490 2943.090 1918.670 ;
        RECT 2941.910 1739.090 2943.090 1740.270 ;
        RECT 2941.910 1737.490 2943.090 1738.670 ;
        RECT 2941.910 1559.090 2943.090 1560.270 ;
        RECT 2941.910 1557.490 2943.090 1558.670 ;
        RECT 2941.910 1379.090 2943.090 1380.270 ;
        RECT 2941.910 1377.490 2943.090 1378.670 ;
        RECT 2941.910 1199.090 2943.090 1200.270 ;
        RECT 2941.910 1197.490 2943.090 1198.670 ;
        RECT 2941.910 1019.090 2943.090 1020.270 ;
        RECT 2941.910 1017.490 2943.090 1018.670 ;
        RECT 2941.910 839.090 2943.090 840.270 ;
        RECT 2941.910 837.490 2943.090 838.670 ;
        RECT 2941.910 659.090 2943.090 660.270 ;
        RECT 2941.910 657.490 2943.090 658.670 ;
        RECT 2941.910 479.090 2943.090 480.270 ;
        RECT 2941.910 477.490 2943.090 478.670 ;
        RECT 2941.910 299.090 2943.090 300.270 ;
        RECT 2941.910 297.490 2943.090 298.670 ;
        RECT 2941.910 119.090 2943.090 120.270 ;
        RECT 2941.910 117.490 2943.090 118.670 ;
        RECT 2812.930 -17.310 2814.110 -16.130 ;
        RECT 2812.930 -18.910 2814.110 -17.730 ;
        RECT 2941.910 -17.310 2943.090 -16.130 ;
        RECT 2941.910 -18.910 2943.090 -17.730 ;
      LAYER met5 ;
        RECT -24.380 3538.700 -21.380 3538.710 ;
        RECT 112.020 3538.700 115.020 3538.710 ;
        RECT 292.020 3538.700 295.020 3538.710 ;
        RECT 472.020 3538.700 475.020 3538.710 ;
        RECT 652.020 3538.700 655.020 3538.710 ;
        RECT 832.020 3538.700 835.020 3538.710 ;
        RECT 1012.020 3538.700 1015.020 3538.710 ;
        RECT 1192.020 3538.700 1195.020 3538.710 ;
        RECT 1372.020 3538.700 1375.020 3538.710 ;
        RECT 1552.020 3538.700 1555.020 3538.710 ;
        RECT 1732.020 3538.700 1735.020 3538.710 ;
        RECT 1912.020 3538.700 1915.020 3538.710 ;
        RECT 2092.020 3538.700 2095.020 3538.710 ;
        RECT 2272.020 3538.700 2275.020 3538.710 ;
        RECT 2452.020 3538.700 2455.020 3538.710 ;
        RECT 2632.020 3538.700 2635.020 3538.710 ;
        RECT 2812.020 3538.700 2815.020 3538.710 ;
        RECT 2941.000 3538.700 2944.000 3538.710 ;
        RECT -24.380 3535.700 2944.000 3538.700 ;
        RECT -24.380 3535.690 -21.380 3535.700 ;
        RECT 112.020 3535.690 115.020 3535.700 ;
        RECT 292.020 3535.690 295.020 3535.700 ;
        RECT 472.020 3535.690 475.020 3535.700 ;
        RECT 652.020 3535.690 655.020 3535.700 ;
        RECT 832.020 3535.690 835.020 3535.700 ;
        RECT 1012.020 3535.690 1015.020 3535.700 ;
        RECT 1192.020 3535.690 1195.020 3535.700 ;
        RECT 1372.020 3535.690 1375.020 3535.700 ;
        RECT 1552.020 3535.690 1555.020 3535.700 ;
        RECT 1732.020 3535.690 1735.020 3535.700 ;
        RECT 1912.020 3535.690 1915.020 3535.700 ;
        RECT 2092.020 3535.690 2095.020 3535.700 ;
        RECT 2272.020 3535.690 2275.020 3535.700 ;
        RECT 2452.020 3535.690 2455.020 3535.700 ;
        RECT 2632.020 3535.690 2635.020 3535.700 ;
        RECT 2812.020 3535.690 2815.020 3535.700 ;
        RECT 2941.000 3535.690 2944.000 3535.700 ;
        RECT -14.780 3529.100 -11.780 3529.110 ;
        RECT 94.020 3529.100 97.020 3529.110 ;
        RECT 274.020 3529.100 277.020 3529.110 ;
        RECT 454.020 3529.100 457.020 3529.110 ;
        RECT 634.020 3529.100 637.020 3529.110 ;
        RECT 814.020 3529.100 817.020 3529.110 ;
        RECT 994.020 3529.100 997.020 3529.110 ;
        RECT 1174.020 3529.100 1177.020 3529.110 ;
        RECT 1354.020 3529.100 1357.020 3529.110 ;
        RECT 1534.020 3529.100 1537.020 3529.110 ;
        RECT 1714.020 3529.100 1717.020 3529.110 ;
        RECT 1894.020 3529.100 1897.020 3529.110 ;
        RECT 2074.020 3529.100 2077.020 3529.110 ;
        RECT 2254.020 3529.100 2257.020 3529.110 ;
        RECT 2434.020 3529.100 2437.020 3529.110 ;
        RECT 2614.020 3529.100 2617.020 3529.110 ;
        RECT 2794.020 3529.100 2797.020 3529.110 ;
        RECT 2931.400 3529.100 2934.400 3529.110 ;
        RECT -14.780 3526.100 2934.400 3529.100 ;
        RECT -14.780 3526.090 -11.780 3526.100 ;
        RECT 94.020 3526.090 97.020 3526.100 ;
        RECT 274.020 3526.090 277.020 3526.100 ;
        RECT 454.020 3526.090 457.020 3526.100 ;
        RECT 634.020 3526.090 637.020 3526.100 ;
        RECT 814.020 3526.090 817.020 3526.100 ;
        RECT 994.020 3526.090 997.020 3526.100 ;
        RECT 1174.020 3526.090 1177.020 3526.100 ;
        RECT 1354.020 3526.090 1357.020 3526.100 ;
        RECT 1534.020 3526.090 1537.020 3526.100 ;
        RECT 1714.020 3526.090 1717.020 3526.100 ;
        RECT 1894.020 3526.090 1897.020 3526.100 ;
        RECT 2074.020 3526.090 2077.020 3526.100 ;
        RECT 2254.020 3526.090 2257.020 3526.100 ;
        RECT 2434.020 3526.090 2437.020 3526.100 ;
        RECT 2614.020 3526.090 2617.020 3526.100 ;
        RECT 2794.020 3526.090 2797.020 3526.100 ;
        RECT 2931.400 3526.090 2934.400 3526.100 ;
        RECT -24.380 3360.380 -21.380 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2941.000 3360.380 2944.000 3360.390 ;
        RECT -24.380 3357.380 2944.000 3360.380 ;
        RECT -24.380 3357.370 -21.380 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2941.000 3357.370 2944.000 3357.380 ;
        RECT -14.780 3342.380 -11.780 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.400 3342.380 2934.400 3342.390 ;
        RECT -14.780 3339.380 2934.400 3342.380 ;
        RECT -14.780 3339.370 -11.780 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.400 3339.370 2934.400 3339.380 ;
        RECT -24.380 3180.380 -21.380 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2941.000 3180.380 2944.000 3180.390 ;
        RECT -24.380 3177.380 2944.000 3180.380 ;
        RECT -24.380 3177.370 -21.380 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2941.000 3177.370 2944.000 3177.380 ;
        RECT -14.780 3162.380 -11.780 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.400 3162.380 2934.400 3162.390 ;
        RECT -14.780 3159.380 2934.400 3162.380 ;
        RECT -14.780 3159.370 -11.780 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.400 3159.370 2934.400 3159.380 ;
        RECT -24.380 3000.380 -21.380 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2941.000 3000.380 2944.000 3000.390 ;
        RECT -24.380 2997.380 2944.000 3000.380 ;
        RECT -24.380 2997.370 -21.380 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2941.000 2997.370 2944.000 2997.380 ;
        RECT -14.780 2982.380 -11.780 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.400 2982.380 2934.400 2982.390 ;
        RECT -14.780 2979.380 2934.400 2982.380 ;
        RECT -14.780 2979.370 -11.780 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.400 2979.370 2934.400 2979.380 ;
        RECT -24.380 2820.380 -21.380 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2941.000 2820.380 2944.000 2820.390 ;
        RECT -24.380 2817.380 2944.000 2820.380 ;
        RECT -24.380 2817.370 -21.380 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2941.000 2817.370 2944.000 2817.380 ;
        RECT -14.780 2802.380 -11.780 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.400 2802.380 2934.400 2802.390 ;
        RECT -14.780 2799.380 2934.400 2802.380 ;
        RECT -14.780 2799.370 -11.780 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.400 2799.370 2934.400 2799.380 ;
        RECT -24.380 2640.380 -21.380 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2941.000 2640.380 2944.000 2640.390 ;
        RECT -24.380 2637.380 2944.000 2640.380 ;
        RECT -24.380 2637.370 -21.380 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2941.000 2637.370 2944.000 2637.380 ;
        RECT -14.780 2622.380 -11.780 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.400 2622.380 2934.400 2622.390 ;
        RECT -14.780 2619.380 2934.400 2622.380 ;
        RECT -14.780 2619.370 -11.780 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.400 2619.370 2934.400 2619.380 ;
        RECT -24.380 2460.380 -21.380 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2941.000 2460.380 2944.000 2460.390 ;
        RECT -24.380 2457.380 2944.000 2460.380 ;
        RECT -24.380 2457.370 -21.380 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2941.000 2457.370 2944.000 2457.380 ;
        RECT -14.780 2442.380 -11.780 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.400 2442.380 2934.400 2442.390 ;
        RECT -14.780 2439.380 2934.400 2442.380 ;
        RECT -14.780 2439.370 -11.780 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.400 2439.370 2934.400 2439.380 ;
        RECT -24.380 2280.380 -21.380 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2941.000 2280.380 2944.000 2280.390 ;
        RECT -24.380 2277.380 2944.000 2280.380 ;
        RECT -24.380 2277.370 -21.380 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2941.000 2277.370 2944.000 2277.380 ;
        RECT -14.780 2262.380 -11.780 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.400 2262.380 2934.400 2262.390 ;
        RECT -14.780 2259.380 2934.400 2262.380 ;
        RECT -14.780 2259.370 -11.780 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.400 2259.370 2934.400 2259.380 ;
        RECT -24.380 2100.380 -21.380 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 507.840 2100.380 509.440 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2941.000 2100.380 2944.000 2100.390 ;
        RECT -24.380 2097.380 2944.000 2100.380 ;
        RECT -24.380 2097.370 -21.380 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 507.840 2097.370 509.440 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2941.000 2097.370 2944.000 2097.380 ;
        RECT -14.780 2082.380 -11.780 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 507.840 2082.380 509.440 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.400 2082.380 2934.400 2082.390 ;
        RECT -14.780 2079.380 2934.400 2082.380 ;
        RECT -14.780 2079.370 -11.780 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 507.840 2079.370 509.440 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.400 2079.370 2934.400 2079.380 ;
        RECT -24.380 1920.380 -21.380 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 507.840 1920.380 509.440 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2941.000 1920.380 2944.000 1920.390 ;
        RECT -24.380 1917.380 2944.000 1920.380 ;
        RECT -24.380 1917.370 -21.380 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 507.840 1917.370 509.440 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2941.000 1917.370 2944.000 1917.380 ;
        RECT -14.780 1902.380 -11.780 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 507.840 1902.380 509.440 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.400 1902.380 2934.400 1902.390 ;
        RECT -14.780 1899.380 2934.400 1902.380 ;
        RECT -14.780 1899.370 -11.780 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 507.840 1899.370 509.440 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.400 1899.370 2934.400 1899.380 ;
        RECT -24.380 1740.380 -21.380 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 507.840 1740.380 509.440 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2941.000 1740.380 2944.000 1740.390 ;
        RECT -24.380 1737.380 2944.000 1740.380 ;
        RECT -24.380 1737.370 -21.380 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 507.840 1737.370 509.440 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2941.000 1737.370 2944.000 1737.380 ;
        RECT -14.780 1722.380 -11.780 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 507.840 1722.380 509.440 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.400 1722.380 2934.400 1722.390 ;
        RECT -14.780 1719.380 2934.400 1722.380 ;
        RECT -14.780 1719.370 -11.780 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 507.840 1719.370 509.440 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.400 1719.370 2934.400 1719.380 ;
        RECT -24.380 1560.380 -21.380 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 507.840 1560.380 509.440 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2941.000 1560.380 2944.000 1560.390 ;
        RECT -24.380 1557.380 2944.000 1560.380 ;
        RECT -24.380 1557.370 -21.380 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 507.840 1557.370 509.440 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2941.000 1557.370 2944.000 1557.380 ;
        RECT -14.780 1542.380 -11.780 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 507.840 1542.380 509.440 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.400 1542.380 2934.400 1542.390 ;
        RECT -14.780 1539.380 2934.400 1542.380 ;
        RECT -14.780 1539.370 -11.780 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 507.840 1539.370 509.440 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.400 1539.370 2934.400 1539.380 ;
        RECT -24.380 1380.380 -21.380 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 507.840 1380.380 509.440 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2941.000 1380.380 2944.000 1380.390 ;
        RECT -24.380 1377.380 2944.000 1380.380 ;
        RECT -24.380 1377.370 -21.380 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 507.840 1377.370 509.440 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2941.000 1377.370 2944.000 1377.380 ;
        RECT -14.780 1362.380 -11.780 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 507.840 1362.380 509.440 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.400 1362.380 2934.400 1362.390 ;
        RECT -14.780 1359.380 2934.400 1362.380 ;
        RECT -14.780 1359.370 -11.780 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 507.840 1359.370 509.440 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.400 1359.370 2934.400 1359.380 ;
        RECT -24.380 1200.380 -21.380 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 507.840 1200.380 509.440 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2941.000 1200.380 2944.000 1200.390 ;
        RECT -24.380 1197.380 2944.000 1200.380 ;
        RECT -24.380 1197.370 -21.380 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 507.840 1197.370 509.440 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2941.000 1197.370 2944.000 1197.380 ;
        RECT -14.780 1182.380 -11.780 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 507.840 1182.380 509.440 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.400 1182.380 2934.400 1182.390 ;
        RECT -14.780 1179.380 2934.400 1182.380 ;
        RECT -14.780 1179.370 -11.780 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 507.840 1179.370 509.440 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.400 1179.370 2934.400 1179.380 ;
        RECT -24.380 1020.380 -21.380 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 507.840 1020.380 509.440 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2941.000 1020.380 2944.000 1020.390 ;
        RECT -24.380 1017.380 2944.000 1020.380 ;
        RECT -24.380 1017.370 -21.380 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 507.840 1017.370 509.440 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2941.000 1017.370 2944.000 1017.380 ;
        RECT -14.780 1002.380 -11.780 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 507.840 1002.380 509.440 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.400 1002.380 2934.400 1002.390 ;
        RECT -14.780 999.380 2934.400 1002.380 ;
        RECT -14.780 999.370 -11.780 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 507.840 999.370 509.440 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.400 999.370 2934.400 999.380 ;
        RECT -24.380 840.380 -21.380 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 507.840 840.380 509.440 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2941.000 840.380 2944.000 840.390 ;
        RECT -24.380 837.380 2944.000 840.380 ;
        RECT -24.380 837.370 -21.380 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 507.840 837.370 509.440 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2941.000 837.370 2944.000 837.380 ;
        RECT -14.780 822.380 -11.780 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 507.840 822.380 509.440 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.400 822.380 2934.400 822.390 ;
        RECT -14.780 819.380 2934.400 822.380 ;
        RECT -14.780 819.370 -11.780 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 507.840 819.370 509.440 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.400 819.370 2934.400 819.380 ;
        RECT -24.380 660.380 -21.380 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 507.840 660.380 509.440 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2941.000 660.380 2944.000 660.390 ;
        RECT -24.380 657.380 2944.000 660.380 ;
        RECT -24.380 657.370 -21.380 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 507.840 657.370 509.440 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2941.000 657.370 2944.000 657.380 ;
        RECT -14.780 642.380 -11.780 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 507.840 642.380 509.440 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.400 642.380 2934.400 642.390 ;
        RECT -14.780 639.380 2934.400 642.380 ;
        RECT -14.780 639.370 -11.780 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 507.840 639.370 509.440 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.400 639.370 2934.400 639.380 ;
        RECT -24.380 480.380 -21.380 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2941.000 480.380 2944.000 480.390 ;
        RECT -24.380 477.380 2944.000 480.380 ;
        RECT -24.380 477.370 -21.380 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2941.000 477.370 2944.000 477.380 ;
        RECT -14.780 462.380 -11.780 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.400 462.380 2934.400 462.390 ;
        RECT -14.780 459.380 2934.400 462.380 ;
        RECT -14.780 459.370 -11.780 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.400 459.370 2934.400 459.380 ;
        RECT -24.380 300.380 -21.380 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2941.000 300.380 2944.000 300.390 ;
        RECT -24.380 297.380 2944.000 300.380 ;
        RECT -24.380 297.370 -21.380 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2941.000 297.370 2944.000 297.380 ;
        RECT -14.780 282.380 -11.780 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.400 282.380 2934.400 282.390 ;
        RECT -14.780 279.380 2934.400 282.380 ;
        RECT -14.780 279.370 -11.780 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.400 279.370 2934.400 279.380 ;
        RECT -24.380 120.380 -21.380 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2941.000 120.380 2944.000 120.390 ;
        RECT -24.380 117.380 2944.000 120.380 ;
        RECT -24.380 117.370 -21.380 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2941.000 117.370 2944.000 117.380 ;
        RECT -14.780 102.380 -11.780 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.400 102.380 2934.400 102.390 ;
        RECT -14.780 99.380 2934.400 102.380 ;
        RECT -14.780 99.370 -11.780 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.400 99.370 2934.400 99.380 ;
        RECT -14.780 -6.420 -11.780 -6.410 ;
        RECT 94.020 -6.420 97.020 -6.410 ;
        RECT 274.020 -6.420 277.020 -6.410 ;
        RECT 454.020 -6.420 457.020 -6.410 ;
        RECT 634.020 -6.420 637.020 -6.410 ;
        RECT 814.020 -6.420 817.020 -6.410 ;
        RECT 994.020 -6.420 997.020 -6.410 ;
        RECT 1174.020 -6.420 1177.020 -6.410 ;
        RECT 1354.020 -6.420 1357.020 -6.410 ;
        RECT 1534.020 -6.420 1537.020 -6.410 ;
        RECT 1714.020 -6.420 1717.020 -6.410 ;
        RECT 1894.020 -6.420 1897.020 -6.410 ;
        RECT 2074.020 -6.420 2077.020 -6.410 ;
        RECT 2254.020 -6.420 2257.020 -6.410 ;
        RECT 2434.020 -6.420 2437.020 -6.410 ;
        RECT 2614.020 -6.420 2617.020 -6.410 ;
        RECT 2794.020 -6.420 2797.020 -6.410 ;
        RECT 2931.400 -6.420 2934.400 -6.410 ;
        RECT -14.780 -9.420 2934.400 -6.420 ;
        RECT -14.780 -9.430 -11.780 -9.420 ;
        RECT 94.020 -9.430 97.020 -9.420 ;
        RECT 274.020 -9.430 277.020 -9.420 ;
        RECT 454.020 -9.430 457.020 -9.420 ;
        RECT 634.020 -9.430 637.020 -9.420 ;
        RECT 814.020 -9.430 817.020 -9.420 ;
        RECT 994.020 -9.430 997.020 -9.420 ;
        RECT 1174.020 -9.430 1177.020 -9.420 ;
        RECT 1354.020 -9.430 1357.020 -9.420 ;
        RECT 1534.020 -9.430 1537.020 -9.420 ;
        RECT 1714.020 -9.430 1717.020 -9.420 ;
        RECT 1894.020 -9.430 1897.020 -9.420 ;
        RECT 2074.020 -9.430 2077.020 -9.420 ;
        RECT 2254.020 -9.430 2257.020 -9.420 ;
        RECT 2434.020 -9.430 2437.020 -9.420 ;
        RECT 2614.020 -9.430 2617.020 -9.420 ;
        RECT 2794.020 -9.430 2797.020 -9.420 ;
        RECT 2931.400 -9.430 2934.400 -9.420 ;
        RECT -24.380 -16.020 -21.380 -16.010 ;
        RECT 112.020 -16.020 115.020 -16.010 ;
        RECT 292.020 -16.020 295.020 -16.010 ;
        RECT 472.020 -16.020 475.020 -16.010 ;
        RECT 652.020 -16.020 655.020 -16.010 ;
        RECT 832.020 -16.020 835.020 -16.010 ;
        RECT 1012.020 -16.020 1015.020 -16.010 ;
        RECT 1192.020 -16.020 1195.020 -16.010 ;
        RECT 1372.020 -16.020 1375.020 -16.010 ;
        RECT 1552.020 -16.020 1555.020 -16.010 ;
        RECT 1732.020 -16.020 1735.020 -16.010 ;
        RECT 1912.020 -16.020 1915.020 -16.010 ;
        RECT 2092.020 -16.020 2095.020 -16.010 ;
        RECT 2272.020 -16.020 2275.020 -16.010 ;
        RECT 2452.020 -16.020 2455.020 -16.010 ;
        RECT 2632.020 -16.020 2635.020 -16.010 ;
        RECT 2812.020 -16.020 2815.020 -16.010 ;
        RECT 2941.000 -16.020 2944.000 -16.010 ;
        RECT -24.380 -19.020 2944.000 -16.020 ;
        RECT -24.380 -19.030 -21.380 -19.020 ;
        RECT 112.020 -19.030 115.020 -19.020 ;
        RECT 292.020 -19.030 295.020 -19.020 ;
        RECT 472.020 -19.030 475.020 -19.020 ;
        RECT 652.020 -19.030 655.020 -19.020 ;
        RECT 832.020 -19.030 835.020 -19.020 ;
        RECT 1012.020 -19.030 1015.020 -19.020 ;
        RECT 1192.020 -19.030 1195.020 -19.020 ;
        RECT 1372.020 -19.030 1375.020 -19.020 ;
        RECT 1552.020 -19.030 1555.020 -19.020 ;
        RECT 1732.020 -19.030 1735.020 -19.020 ;
        RECT 1912.020 -19.030 1915.020 -19.020 ;
        RECT 2092.020 -19.030 2095.020 -19.020 ;
        RECT 2272.020 -19.030 2275.020 -19.020 ;
        RECT 2452.020 -19.030 2455.020 -19.020 ;
        RECT 2632.020 -19.030 2635.020 -19.020 ;
        RECT 2812.020 -19.030 2815.020 -19.020 ;
        RECT 2941.000 -19.030 2944.000 -19.020 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 415.520 520.795 1995.620 2101.285 ;
      LAYER met1 ;
        RECT 411.910 519.560 1995.620 2101.440 ;
      LAYER met2 ;
        RECT 411.940 2107.905 439.250 2108.185 ;
        RECT 440.090 2107.905 498.130 2108.185 ;
        RECT 498.970 2107.905 557.010 2108.185 ;
        RECT 557.850 2107.905 615.890 2108.185 ;
        RECT 616.730 2107.905 674.770 2108.185 ;
        RECT 675.610 2107.905 733.650 2108.185 ;
        RECT 734.490 2107.905 792.530 2108.185 ;
        RECT 793.370 2107.905 851.870 2108.185 ;
        RECT 852.710 2107.905 910.750 2108.185 ;
        RECT 911.590 2107.905 969.630 2108.185 ;
        RECT 970.470 2107.905 1028.510 2108.185 ;
        RECT 1029.350 2107.905 1087.390 2108.185 ;
        RECT 1088.230 2107.905 1146.270 2108.185 ;
        RECT 1147.110 2107.905 1205.150 2108.185 ;
        RECT 1205.990 2107.905 1264.490 2108.185 ;
        RECT 1265.330 2107.905 1323.370 2108.185 ;
        RECT 1324.210 2107.905 1382.250 2108.185 ;
        RECT 1383.090 2107.905 1441.130 2108.185 ;
        RECT 1441.970 2107.905 1500.010 2108.185 ;
        RECT 1500.850 2107.905 1558.890 2108.185 ;
        RECT 1559.730 2107.905 1617.770 2108.185 ;
        RECT 1618.610 2107.905 1677.110 2108.185 ;
        RECT 1677.950 2107.905 1735.990 2108.185 ;
        RECT 1736.830 2107.905 1794.870 2108.185 ;
        RECT 1795.710 2107.905 1853.750 2108.185 ;
        RECT 1854.590 2107.905 1912.630 2108.185 ;
        RECT 1913.470 2107.905 1971.510 2108.185 ;
        RECT 1972.350 2107.905 1995.520 2108.185 ;
        RECT 411.940 514.280 1995.520 2107.905 ;
        RECT 412.490 514.000 415.330 514.280 ;
        RECT 416.170 514.000 419.470 514.280 ;
        RECT 420.310 514.000 423.610 514.280 ;
        RECT 424.450 514.000 427.750 514.280 ;
        RECT 428.590 514.000 431.890 514.280 ;
        RECT 432.730 514.000 436.030 514.280 ;
        RECT 436.870 514.000 440.170 514.280 ;
        RECT 441.010 514.000 444.310 514.280 ;
        RECT 445.150 514.000 448.450 514.280 ;
        RECT 449.290 514.000 452.590 514.280 ;
        RECT 453.430 514.000 456.730 514.280 ;
        RECT 457.570 514.000 460.870 514.280 ;
        RECT 461.710 514.000 465.010 514.280 ;
        RECT 465.850 514.000 469.150 514.280 ;
        RECT 469.990 514.000 473.290 514.280 ;
        RECT 474.130 514.000 477.430 514.280 ;
        RECT 478.270 514.000 481.570 514.280 ;
        RECT 482.410 514.000 485.710 514.280 ;
        RECT 486.550 514.000 489.850 514.280 ;
        RECT 490.690 514.000 493.990 514.280 ;
        RECT 494.830 514.000 498.130 514.280 ;
        RECT 498.970 514.000 502.270 514.280 ;
        RECT 503.110 514.000 506.410 514.280 ;
        RECT 507.250 514.000 510.550 514.280 ;
        RECT 511.390 514.000 514.690 514.280 ;
        RECT 515.530 514.000 518.830 514.280 ;
        RECT 519.670 514.000 522.970 514.280 ;
        RECT 523.810 514.000 526.650 514.280 ;
        RECT 527.490 514.000 530.790 514.280 ;
        RECT 531.630 514.000 534.930 514.280 ;
        RECT 535.770 514.000 539.070 514.280 ;
        RECT 539.910 514.000 543.210 514.280 ;
        RECT 544.050 514.000 547.350 514.280 ;
        RECT 548.190 514.000 551.490 514.280 ;
        RECT 552.330 514.000 555.630 514.280 ;
        RECT 556.470 514.000 559.770 514.280 ;
        RECT 560.610 514.000 563.910 514.280 ;
        RECT 564.750 514.000 568.050 514.280 ;
        RECT 568.890 514.000 572.190 514.280 ;
        RECT 573.030 514.000 576.330 514.280 ;
        RECT 577.170 514.000 580.470 514.280 ;
        RECT 581.310 514.000 584.610 514.280 ;
        RECT 585.450 514.000 588.750 514.280 ;
        RECT 589.590 514.000 592.890 514.280 ;
        RECT 593.730 514.000 597.030 514.280 ;
        RECT 597.870 514.000 601.170 514.280 ;
        RECT 602.010 514.000 605.310 514.280 ;
        RECT 606.150 514.000 609.450 514.280 ;
        RECT 610.290 514.000 613.590 514.280 ;
        RECT 614.430 514.000 617.730 514.280 ;
        RECT 618.570 514.000 621.870 514.280 ;
        RECT 622.710 514.000 626.010 514.280 ;
        RECT 626.850 514.000 630.150 514.280 ;
        RECT 630.990 514.000 634.290 514.280 ;
        RECT 635.130 514.000 638.430 514.280 ;
        RECT 639.270 514.000 642.110 514.280 ;
        RECT 642.950 514.000 646.250 514.280 ;
        RECT 647.090 514.000 650.390 514.280 ;
        RECT 651.230 514.000 654.530 514.280 ;
        RECT 655.370 514.000 658.670 514.280 ;
        RECT 659.510 514.000 662.810 514.280 ;
        RECT 663.650 514.000 666.950 514.280 ;
        RECT 667.790 514.000 671.090 514.280 ;
        RECT 671.930 514.000 675.230 514.280 ;
        RECT 676.070 514.000 679.370 514.280 ;
        RECT 680.210 514.000 683.510 514.280 ;
        RECT 684.350 514.000 687.650 514.280 ;
        RECT 688.490 514.000 691.790 514.280 ;
        RECT 692.630 514.000 695.930 514.280 ;
        RECT 696.770 514.000 700.070 514.280 ;
        RECT 700.910 514.000 704.210 514.280 ;
        RECT 705.050 514.000 708.350 514.280 ;
        RECT 709.190 514.000 712.490 514.280 ;
        RECT 713.330 514.000 716.630 514.280 ;
        RECT 717.470 514.000 720.770 514.280 ;
        RECT 721.610 514.000 724.910 514.280 ;
        RECT 725.750 514.000 729.050 514.280 ;
        RECT 729.890 514.000 733.190 514.280 ;
        RECT 734.030 514.000 737.330 514.280 ;
        RECT 738.170 514.000 741.470 514.280 ;
        RECT 742.310 514.000 745.610 514.280 ;
        RECT 746.450 514.000 749.750 514.280 ;
        RECT 750.590 514.000 753.430 514.280 ;
        RECT 754.270 514.000 757.570 514.280 ;
        RECT 758.410 514.000 761.710 514.280 ;
        RECT 762.550 514.000 765.850 514.280 ;
        RECT 766.690 514.000 769.990 514.280 ;
        RECT 770.830 514.000 774.130 514.280 ;
        RECT 774.970 514.000 778.270 514.280 ;
        RECT 779.110 514.000 782.410 514.280 ;
        RECT 783.250 514.000 786.550 514.280 ;
        RECT 787.390 514.000 790.690 514.280 ;
        RECT 791.530 514.000 794.830 514.280 ;
        RECT 795.670 514.000 798.970 514.280 ;
        RECT 799.810 514.000 803.110 514.280 ;
        RECT 803.950 514.000 807.250 514.280 ;
        RECT 808.090 514.000 811.390 514.280 ;
        RECT 812.230 514.000 815.530 514.280 ;
        RECT 816.370 514.000 819.670 514.280 ;
        RECT 820.510 514.000 823.810 514.280 ;
        RECT 824.650 514.000 827.950 514.280 ;
        RECT 828.790 514.000 832.090 514.280 ;
        RECT 832.930 514.000 836.230 514.280 ;
        RECT 837.070 514.000 840.370 514.280 ;
        RECT 841.210 514.000 844.510 514.280 ;
        RECT 845.350 514.000 848.650 514.280 ;
        RECT 849.490 514.000 852.790 514.280 ;
        RECT 853.630 514.000 856.930 514.280 ;
        RECT 857.770 514.000 861.070 514.280 ;
        RECT 861.910 514.000 865.210 514.280 ;
        RECT 866.050 514.000 868.890 514.280 ;
        RECT 869.730 514.000 873.030 514.280 ;
        RECT 873.870 514.000 877.170 514.280 ;
        RECT 878.010 514.000 881.310 514.280 ;
        RECT 882.150 514.000 885.450 514.280 ;
        RECT 886.290 514.000 889.590 514.280 ;
        RECT 890.430 514.000 893.730 514.280 ;
        RECT 894.570 514.000 897.870 514.280 ;
        RECT 898.710 514.000 902.010 514.280 ;
        RECT 902.850 514.000 906.150 514.280 ;
        RECT 906.990 514.000 910.290 514.280 ;
        RECT 911.130 514.000 914.430 514.280 ;
        RECT 915.270 514.000 918.570 514.280 ;
        RECT 919.410 514.000 922.710 514.280 ;
        RECT 923.550 514.000 926.850 514.280 ;
        RECT 927.690 514.000 930.990 514.280 ;
        RECT 931.830 514.000 935.130 514.280 ;
        RECT 935.970 514.000 939.270 514.280 ;
        RECT 940.110 514.000 943.410 514.280 ;
        RECT 944.250 514.000 947.550 514.280 ;
        RECT 948.390 514.000 951.690 514.280 ;
        RECT 952.530 514.000 955.830 514.280 ;
        RECT 956.670 514.000 959.970 514.280 ;
        RECT 960.810 514.000 964.110 514.280 ;
        RECT 964.950 514.000 968.250 514.280 ;
        RECT 969.090 514.000 972.390 514.280 ;
        RECT 973.230 514.000 976.530 514.280 ;
        RECT 977.370 514.000 980.210 514.280 ;
        RECT 981.050 514.000 984.350 514.280 ;
        RECT 985.190 514.000 988.490 514.280 ;
        RECT 989.330 514.000 992.630 514.280 ;
        RECT 993.470 514.000 996.770 514.280 ;
        RECT 997.610 514.000 1000.910 514.280 ;
        RECT 1001.750 514.000 1005.050 514.280 ;
        RECT 1005.890 514.000 1009.190 514.280 ;
        RECT 1010.030 514.000 1013.330 514.280 ;
        RECT 1014.170 514.000 1017.470 514.280 ;
        RECT 1018.310 514.000 1021.610 514.280 ;
        RECT 1022.450 514.000 1025.750 514.280 ;
        RECT 1026.590 514.000 1029.890 514.280 ;
        RECT 1030.730 514.000 1034.030 514.280 ;
        RECT 1034.870 514.000 1038.170 514.280 ;
        RECT 1039.010 514.000 1042.310 514.280 ;
        RECT 1043.150 514.000 1046.450 514.280 ;
        RECT 1047.290 514.000 1050.590 514.280 ;
        RECT 1051.430 514.000 1054.730 514.280 ;
        RECT 1055.570 514.000 1058.870 514.280 ;
        RECT 1059.710 514.000 1063.010 514.280 ;
        RECT 1063.850 514.000 1067.150 514.280 ;
        RECT 1067.990 514.000 1071.290 514.280 ;
        RECT 1072.130 514.000 1075.430 514.280 ;
        RECT 1076.270 514.000 1079.570 514.280 ;
        RECT 1080.410 514.000 1083.710 514.280 ;
        RECT 1084.550 514.000 1087.850 514.280 ;
        RECT 1088.690 514.000 1091.990 514.280 ;
        RECT 1092.830 514.000 1095.670 514.280 ;
        RECT 1096.510 514.000 1099.810 514.280 ;
        RECT 1100.650 514.000 1103.950 514.280 ;
        RECT 1104.790 514.000 1108.090 514.280 ;
        RECT 1108.930 514.000 1112.230 514.280 ;
        RECT 1113.070 514.000 1116.370 514.280 ;
        RECT 1117.210 514.000 1120.510 514.280 ;
        RECT 1121.350 514.000 1124.650 514.280 ;
        RECT 1125.490 514.000 1128.790 514.280 ;
        RECT 1129.630 514.000 1132.930 514.280 ;
        RECT 1133.770 514.000 1137.070 514.280 ;
        RECT 1137.910 514.000 1141.210 514.280 ;
        RECT 1142.050 514.000 1145.350 514.280 ;
        RECT 1146.190 514.000 1149.490 514.280 ;
        RECT 1150.330 514.000 1153.630 514.280 ;
        RECT 1154.470 514.000 1157.770 514.280 ;
        RECT 1158.610 514.000 1161.910 514.280 ;
        RECT 1162.750 514.000 1166.050 514.280 ;
        RECT 1166.890 514.000 1170.190 514.280 ;
        RECT 1171.030 514.000 1174.330 514.280 ;
        RECT 1175.170 514.000 1178.470 514.280 ;
        RECT 1179.310 514.000 1182.610 514.280 ;
        RECT 1183.450 514.000 1186.750 514.280 ;
        RECT 1187.590 514.000 1190.890 514.280 ;
        RECT 1191.730 514.000 1195.030 514.280 ;
        RECT 1195.870 514.000 1199.170 514.280 ;
        RECT 1200.010 514.000 1203.310 514.280 ;
        RECT 1204.150 514.000 1207.450 514.280 ;
        RECT 1208.290 514.000 1211.130 514.280 ;
        RECT 1211.970 514.000 1215.270 514.280 ;
        RECT 1216.110 514.000 1219.410 514.280 ;
        RECT 1220.250 514.000 1223.550 514.280 ;
        RECT 1224.390 514.000 1227.690 514.280 ;
        RECT 1228.530 514.000 1231.830 514.280 ;
        RECT 1232.670 514.000 1235.970 514.280 ;
        RECT 1236.810 514.000 1240.110 514.280 ;
        RECT 1240.950 514.000 1244.250 514.280 ;
        RECT 1245.090 514.000 1248.390 514.280 ;
        RECT 1249.230 514.000 1252.530 514.280 ;
        RECT 1253.370 514.000 1256.670 514.280 ;
        RECT 1257.510 514.000 1260.810 514.280 ;
        RECT 1261.650 514.000 1264.950 514.280 ;
        RECT 1265.790 514.000 1269.090 514.280 ;
        RECT 1269.930 514.000 1273.230 514.280 ;
        RECT 1274.070 514.000 1277.370 514.280 ;
        RECT 1278.210 514.000 1281.510 514.280 ;
        RECT 1282.350 514.000 1285.650 514.280 ;
        RECT 1286.490 514.000 1289.790 514.280 ;
        RECT 1290.630 514.000 1293.930 514.280 ;
        RECT 1294.770 514.000 1298.070 514.280 ;
        RECT 1298.910 514.000 1302.210 514.280 ;
        RECT 1303.050 514.000 1306.350 514.280 ;
        RECT 1307.190 514.000 1310.490 514.280 ;
        RECT 1311.330 514.000 1314.630 514.280 ;
        RECT 1315.470 514.000 1318.770 514.280 ;
        RECT 1319.610 514.000 1322.450 514.280 ;
        RECT 1323.290 514.000 1326.590 514.280 ;
        RECT 1327.430 514.000 1330.730 514.280 ;
        RECT 1331.570 514.000 1334.870 514.280 ;
        RECT 1335.710 514.000 1339.010 514.280 ;
        RECT 1339.850 514.000 1343.150 514.280 ;
        RECT 1343.990 514.000 1347.290 514.280 ;
        RECT 1348.130 514.000 1351.430 514.280 ;
        RECT 1352.270 514.000 1355.570 514.280 ;
        RECT 1356.410 514.000 1359.710 514.280 ;
        RECT 1360.550 514.000 1363.850 514.280 ;
        RECT 1364.690 514.000 1367.990 514.280 ;
        RECT 1368.830 514.000 1372.130 514.280 ;
        RECT 1372.970 514.000 1376.270 514.280 ;
        RECT 1377.110 514.000 1380.410 514.280 ;
        RECT 1381.250 514.000 1384.550 514.280 ;
        RECT 1385.390 514.000 1388.690 514.280 ;
        RECT 1389.530 514.000 1392.830 514.280 ;
        RECT 1393.670 514.000 1396.970 514.280 ;
        RECT 1397.810 514.000 1401.110 514.280 ;
        RECT 1401.950 514.000 1405.250 514.280 ;
        RECT 1406.090 514.000 1409.390 514.280 ;
        RECT 1410.230 514.000 1413.530 514.280 ;
        RECT 1414.370 514.000 1417.670 514.280 ;
        RECT 1418.510 514.000 1421.810 514.280 ;
        RECT 1422.650 514.000 1425.950 514.280 ;
        RECT 1426.790 514.000 1430.090 514.280 ;
        RECT 1430.930 514.000 1434.230 514.280 ;
        RECT 1435.070 514.000 1437.910 514.280 ;
        RECT 1438.750 514.000 1442.050 514.280 ;
        RECT 1442.890 514.000 1446.190 514.280 ;
        RECT 1447.030 514.000 1450.330 514.280 ;
        RECT 1451.170 514.000 1454.470 514.280 ;
        RECT 1455.310 514.000 1458.610 514.280 ;
        RECT 1459.450 514.000 1462.750 514.280 ;
        RECT 1463.590 514.000 1466.890 514.280 ;
        RECT 1467.730 514.000 1471.030 514.280 ;
        RECT 1471.870 514.000 1475.170 514.280 ;
        RECT 1476.010 514.000 1479.310 514.280 ;
        RECT 1480.150 514.000 1483.450 514.280 ;
        RECT 1484.290 514.000 1487.590 514.280 ;
        RECT 1488.430 514.000 1491.730 514.280 ;
        RECT 1492.570 514.000 1495.870 514.280 ;
        RECT 1496.710 514.000 1500.010 514.280 ;
        RECT 1500.850 514.000 1504.150 514.280 ;
        RECT 1504.990 514.000 1508.290 514.280 ;
        RECT 1509.130 514.000 1512.430 514.280 ;
        RECT 1513.270 514.000 1516.570 514.280 ;
        RECT 1517.410 514.000 1520.710 514.280 ;
        RECT 1521.550 514.000 1524.850 514.280 ;
        RECT 1525.690 514.000 1528.990 514.280 ;
        RECT 1529.830 514.000 1533.130 514.280 ;
        RECT 1533.970 514.000 1537.270 514.280 ;
        RECT 1538.110 514.000 1541.410 514.280 ;
        RECT 1542.250 514.000 1545.550 514.280 ;
        RECT 1546.390 514.000 1549.230 514.280 ;
        RECT 1550.070 514.000 1553.370 514.280 ;
        RECT 1554.210 514.000 1557.510 514.280 ;
        RECT 1558.350 514.000 1561.650 514.280 ;
        RECT 1562.490 514.000 1565.790 514.280 ;
        RECT 1566.630 514.000 1569.930 514.280 ;
        RECT 1570.770 514.000 1574.070 514.280 ;
        RECT 1574.910 514.000 1578.210 514.280 ;
        RECT 1579.050 514.000 1582.350 514.280 ;
        RECT 1583.190 514.000 1586.490 514.280 ;
        RECT 1587.330 514.000 1590.630 514.280 ;
        RECT 1591.470 514.000 1594.770 514.280 ;
        RECT 1595.610 514.000 1598.910 514.280 ;
        RECT 1599.750 514.000 1603.050 514.280 ;
        RECT 1603.890 514.000 1607.190 514.280 ;
        RECT 1608.030 514.000 1611.330 514.280 ;
        RECT 1612.170 514.000 1615.470 514.280 ;
        RECT 1616.310 514.000 1619.610 514.280 ;
        RECT 1620.450 514.000 1623.750 514.280 ;
        RECT 1624.590 514.000 1627.890 514.280 ;
        RECT 1628.730 514.000 1632.030 514.280 ;
        RECT 1632.870 514.000 1636.170 514.280 ;
        RECT 1637.010 514.000 1640.310 514.280 ;
        RECT 1641.150 514.000 1644.450 514.280 ;
        RECT 1645.290 514.000 1648.590 514.280 ;
        RECT 1649.430 514.000 1652.730 514.280 ;
        RECT 1653.570 514.000 1656.870 514.280 ;
        RECT 1657.710 514.000 1661.010 514.280 ;
        RECT 1661.850 514.000 1664.690 514.280 ;
        RECT 1665.530 514.000 1668.830 514.280 ;
        RECT 1669.670 514.000 1672.970 514.280 ;
        RECT 1673.810 514.000 1677.110 514.280 ;
        RECT 1677.950 514.000 1681.250 514.280 ;
        RECT 1682.090 514.000 1685.390 514.280 ;
        RECT 1686.230 514.000 1689.530 514.280 ;
        RECT 1690.370 514.000 1693.670 514.280 ;
        RECT 1694.510 514.000 1697.810 514.280 ;
        RECT 1698.650 514.000 1701.950 514.280 ;
        RECT 1702.790 514.000 1706.090 514.280 ;
        RECT 1706.930 514.000 1710.230 514.280 ;
        RECT 1711.070 514.000 1714.370 514.280 ;
        RECT 1715.210 514.000 1718.510 514.280 ;
        RECT 1719.350 514.000 1722.650 514.280 ;
        RECT 1723.490 514.000 1726.790 514.280 ;
        RECT 1727.630 514.000 1730.930 514.280 ;
        RECT 1731.770 514.000 1735.070 514.280 ;
        RECT 1735.910 514.000 1739.210 514.280 ;
        RECT 1740.050 514.000 1743.350 514.280 ;
        RECT 1744.190 514.000 1747.490 514.280 ;
        RECT 1748.330 514.000 1751.630 514.280 ;
        RECT 1752.470 514.000 1755.770 514.280 ;
        RECT 1756.610 514.000 1759.910 514.280 ;
        RECT 1760.750 514.000 1764.050 514.280 ;
        RECT 1764.890 514.000 1768.190 514.280 ;
        RECT 1769.030 514.000 1772.330 514.280 ;
        RECT 1773.170 514.000 1776.010 514.280 ;
        RECT 1776.850 514.000 1780.150 514.280 ;
        RECT 1780.990 514.000 1784.290 514.280 ;
        RECT 1785.130 514.000 1788.430 514.280 ;
        RECT 1789.270 514.000 1792.570 514.280 ;
        RECT 1793.410 514.000 1796.710 514.280 ;
        RECT 1797.550 514.000 1800.850 514.280 ;
        RECT 1801.690 514.000 1804.990 514.280 ;
        RECT 1805.830 514.000 1809.130 514.280 ;
        RECT 1809.970 514.000 1813.270 514.280 ;
        RECT 1814.110 514.000 1817.410 514.280 ;
        RECT 1818.250 514.000 1821.550 514.280 ;
        RECT 1822.390 514.000 1825.690 514.280 ;
        RECT 1826.530 514.000 1829.830 514.280 ;
        RECT 1830.670 514.000 1833.970 514.280 ;
        RECT 1834.810 514.000 1838.110 514.280 ;
        RECT 1838.950 514.000 1842.250 514.280 ;
        RECT 1843.090 514.000 1846.390 514.280 ;
        RECT 1847.230 514.000 1850.530 514.280 ;
        RECT 1851.370 514.000 1854.670 514.280 ;
        RECT 1855.510 514.000 1858.810 514.280 ;
        RECT 1859.650 514.000 1862.950 514.280 ;
        RECT 1863.790 514.000 1867.090 514.280 ;
        RECT 1867.930 514.000 1871.230 514.280 ;
        RECT 1872.070 514.000 1875.370 514.280 ;
        RECT 1876.210 514.000 1879.510 514.280 ;
        RECT 1880.350 514.000 1883.650 514.280 ;
        RECT 1884.490 514.000 1887.790 514.280 ;
        RECT 1888.630 514.000 1891.470 514.280 ;
        RECT 1892.310 514.000 1895.610 514.280 ;
        RECT 1896.450 514.000 1899.750 514.280 ;
        RECT 1900.590 514.000 1903.890 514.280 ;
        RECT 1904.730 514.000 1908.030 514.280 ;
        RECT 1908.870 514.000 1912.170 514.280 ;
        RECT 1913.010 514.000 1916.310 514.280 ;
        RECT 1917.150 514.000 1920.450 514.280 ;
        RECT 1921.290 514.000 1924.590 514.280 ;
        RECT 1925.430 514.000 1928.730 514.280 ;
        RECT 1929.570 514.000 1932.870 514.280 ;
        RECT 1933.710 514.000 1937.010 514.280 ;
        RECT 1937.850 514.000 1941.150 514.280 ;
        RECT 1941.990 514.000 1945.290 514.280 ;
        RECT 1946.130 514.000 1949.430 514.280 ;
        RECT 1950.270 514.000 1953.570 514.280 ;
        RECT 1954.410 514.000 1957.710 514.280 ;
        RECT 1958.550 514.000 1961.850 514.280 ;
        RECT 1962.690 514.000 1965.990 514.280 ;
        RECT 1966.830 514.000 1970.130 514.280 ;
        RECT 1970.970 514.000 1974.270 514.280 ;
        RECT 1975.110 514.000 1978.410 514.280 ;
        RECT 1979.250 514.000 1982.550 514.280 ;
        RECT 1983.390 514.000 1986.690 514.280 ;
        RECT 1987.530 514.000 1990.830 514.280 ;
        RECT 1991.670 514.000 1994.970 514.280 ;
      LAYER met3 ;
        RECT 413.990 2094.760 1997.610 2101.365 ;
        RECT 413.990 2093.400 1997.065 2094.760 ;
        RECT 414.400 2093.360 1997.065 2093.400 ;
        RECT 414.400 2092.000 1997.610 2093.360 ;
        RECT 413.990 2059.400 1997.610 2092.000 ;
        RECT 413.990 2058.000 1997.065 2059.400 ;
        RECT 413.990 2055.320 1997.610 2058.000 ;
        RECT 414.400 2053.920 1997.610 2055.320 ;
        RECT 413.990 2023.360 1997.610 2053.920 ;
        RECT 413.990 2021.960 1997.065 2023.360 ;
        RECT 413.990 2017.240 1997.610 2021.960 ;
        RECT 414.400 2015.840 1997.610 2017.240 ;
        RECT 413.990 1988.000 1997.610 2015.840 ;
        RECT 413.990 1986.600 1997.065 1988.000 ;
        RECT 413.990 1979.160 1997.610 1986.600 ;
        RECT 414.400 1977.760 1997.610 1979.160 ;
        RECT 413.990 1952.640 1997.610 1977.760 ;
        RECT 413.990 1951.240 1997.065 1952.640 ;
        RECT 413.990 1941.080 1997.610 1951.240 ;
        RECT 414.400 1939.680 1997.610 1941.080 ;
        RECT 413.990 1916.600 1997.610 1939.680 ;
        RECT 413.990 1915.200 1997.065 1916.600 ;
        RECT 413.990 1903.000 1997.610 1915.200 ;
        RECT 414.400 1901.600 1997.610 1903.000 ;
        RECT 413.990 1881.240 1997.610 1901.600 ;
        RECT 413.990 1879.840 1997.065 1881.240 ;
        RECT 413.990 1864.920 1997.610 1879.840 ;
        RECT 414.400 1863.520 1997.610 1864.920 ;
        RECT 413.990 1845.880 1997.610 1863.520 ;
        RECT 413.990 1844.480 1997.065 1845.880 ;
        RECT 413.990 1826.840 1997.610 1844.480 ;
        RECT 414.400 1825.440 1997.610 1826.840 ;
        RECT 413.990 1809.840 1997.610 1825.440 ;
        RECT 413.990 1808.440 1997.065 1809.840 ;
        RECT 413.990 1788.760 1997.610 1808.440 ;
        RECT 414.400 1787.360 1997.610 1788.760 ;
        RECT 413.990 1774.480 1997.610 1787.360 ;
        RECT 413.990 1773.080 1997.065 1774.480 ;
        RECT 413.990 1750.680 1997.610 1773.080 ;
        RECT 414.400 1749.280 1997.610 1750.680 ;
        RECT 413.990 1739.120 1997.610 1749.280 ;
        RECT 413.990 1737.720 1997.065 1739.120 ;
        RECT 413.990 1711.920 1997.610 1737.720 ;
        RECT 414.400 1710.520 1997.610 1711.920 ;
        RECT 413.990 1703.080 1997.610 1710.520 ;
        RECT 413.990 1701.680 1997.065 1703.080 ;
        RECT 413.990 1673.840 1997.610 1701.680 ;
        RECT 414.400 1672.440 1997.610 1673.840 ;
        RECT 413.990 1667.720 1997.610 1672.440 ;
        RECT 413.990 1666.320 1997.065 1667.720 ;
        RECT 413.990 1635.760 1997.610 1666.320 ;
        RECT 414.400 1634.360 1997.610 1635.760 ;
        RECT 413.990 1632.360 1997.610 1634.360 ;
        RECT 413.990 1630.960 1997.065 1632.360 ;
        RECT 413.990 1597.680 1997.610 1630.960 ;
        RECT 414.400 1596.320 1997.610 1597.680 ;
        RECT 414.400 1596.280 1997.065 1596.320 ;
        RECT 413.990 1594.920 1997.065 1596.280 ;
        RECT 413.990 1560.960 1997.610 1594.920 ;
        RECT 413.990 1559.600 1997.065 1560.960 ;
        RECT 414.400 1559.560 1997.065 1559.600 ;
        RECT 414.400 1558.200 1997.610 1559.560 ;
        RECT 413.990 1524.920 1997.610 1558.200 ;
        RECT 413.990 1523.520 1997.065 1524.920 ;
        RECT 413.990 1521.520 1997.610 1523.520 ;
        RECT 414.400 1520.120 1997.610 1521.520 ;
        RECT 413.990 1489.560 1997.610 1520.120 ;
        RECT 413.990 1488.160 1997.065 1489.560 ;
        RECT 413.990 1483.440 1997.610 1488.160 ;
        RECT 414.400 1482.040 1997.610 1483.440 ;
        RECT 413.990 1454.200 1997.610 1482.040 ;
        RECT 413.990 1452.800 1997.065 1454.200 ;
        RECT 413.990 1445.360 1997.610 1452.800 ;
        RECT 414.400 1443.960 1997.610 1445.360 ;
        RECT 413.990 1418.160 1997.610 1443.960 ;
        RECT 413.990 1416.760 1997.065 1418.160 ;
        RECT 413.990 1407.280 1997.610 1416.760 ;
        RECT 414.400 1405.880 1997.610 1407.280 ;
        RECT 413.990 1382.800 1997.610 1405.880 ;
        RECT 413.990 1381.400 1997.065 1382.800 ;
        RECT 413.990 1369.200 1997.610 1381.400 ;
        RECT 414.400 1367.800 1997.610 1369.200 ;
        RECT 413.990 1347.440 1997.610 1367.800 ;
        RECT 413.990 1346.040 1997.065 1347.440 ;
        RECT 413.990 1331.120 1997.610 1346.040 ;
        RECT 414.400 1329.720 1997.610 1331.120 ;
        RECT 413.990 1311.400 1997.610 1329.720 ;
        RECT 413.990 1310.000 1997.065 1311.400 ;
        RECT 413.990 1292.360 1997.610 1310.000 ;
        RECT 414.400 1290.960 1997.610 1292.360 ;
        RECT 413.990 1276.040 1997.610 1290.960 ;
        RECT 413.990 1274.640 1997.065 1276.040 ;
        RECT 413.990 1254.280 1997.610 1274.640 ;
        RECT 414.400 1252.880 1997.610 1254.280 ;
        RECT 413.990 1240.680 1997.610 1252.880 ;
        RECT 413.990 1239.280 1997.065 1240.680 ;
        RECT 413.990 1216.200 1997.610 1239.280 ;
        RECT 414.400 1214.800 1997.610 1216.200 ;
        RECT 413.990 1204.640 1997.610 1214.800 ;
        RECT 413.990 1203.240 1997.065 1204.640 ;
        RECT 413.990 1178.120 1997.610 1203.240 ;
        RECT 414.400 1176.720 1997.610 1178.120 ;
        RECT 413.990 1169.280 1997.610 1176.720 ;
        RECT 413.990 1167.880 1997.065 1169.280 ;
        RECT 413.990 1140.040 1997.610 1167.880 ;
        RECT 414.400 1138.640 1997.610 1140.040 ;
        RECT 413.990 1133.920 1997.610 1138.640 ;
        RECT 413.990 1132.520 1997.065 1133.920 ;
        RECT 413.990 1101.960 1997.610 1132.520 ;
        RECT 414.400 1100.560 1997.610 1101.960 ;
        RECT 413.990 1097.880 1997.610 1100.560 ;
        RECT 413.990 1096.480 1997.065 1097.880 ;
        RECT 413.990 1063.880 1997.610 1096.480 ;
        RECT 414.400 1062.520 1997.610 1063.880 ;
        RECT 414.400 1062.480 1997.065 1062.520 ;
        RECT 413.990 1061.120 1997.065 1062.480 ;
        RECT 413.990 1026.480 1997.610 1061.120 ;
        RECT 413.990 1025.800 1997.065 1026.480 ;
        RECT 414.400 1025.080 1997.065 1025.800 ;
        RECT 414.400 1024.400 1997.610 1025.080 ;
        RECT 413.990 991.120 1997.610 1024.400 ;
        RECT 413.990 989.720 1997.065 991.120 ;
        RECT 413.990 987.720 1997.610 989.720 ;
        RECT 414.400 986.320 1997.610 987.720 ;
        RECT 413.990 955.760 1997.610 986.320 ;
        RECT 413.990 954.360 1997.065 955.760 ;
        RECT 413.990 949.640 1997.610 954.360 ;
        RECT 414.400 948.240 1997.610 949.640 ;
        RECT 413.990 919.720 1997.610 948.240 ;
        RECT 413.990 918.320 1997.065 919.720 ;
        RECT 413.990 910.880 1997.610 918.320 ;
        RECT 414.400 909.480 1997.610 910.880 ;
        RECT 413.990 884.360 1997.610 909.480 ;
        RECT 413.990 882.960 1997.065 884.360 ;
        RECT 413.990 872.800 1997.610 882.960 ;
        RECT 414.400 871.400 1997.610 872.800 ;
        RECT 413.990 849.000 1997.610 871.400 ;
        RECT 413.990 847.600 1997.065 849.000 ;
        RECT 413.990 834.720 1997.610 847.600 ;
        RECT 414.400 833.320 1997.610 834.720 ;
        RECT 413.990 812.960 1997.610 833.320 ;
        RECT 413.990 811.560 1997.065 812.960 ;
        RECT 413.990 796.640 1997.610 811.560 ;
        RECT 414.400 795.240 1997.610 796.640 ;
        RECT 413.990 777.600 1997.610 795.240 ;
        RECT 413.990 776.200 1997.065 777.600 ;
        RECT 413.990 758.560 1997.610 776.200 ;
        RECT 414.400 757.160 1997.610 758.560 ;
        RECT 413.990 742.240 1997.610 757.160 ;
        RECT 413.990 740.840 1997.065 742.240 ;
        RECT 413.990 720.480 1997.610 740.840 ;
        RECT 414.400 719.080 1997.610 720.480 ;
        RECT 413.990 706.200 1997.610 719.080 ;
        RECT 413.990 704.800 1997.065 706.200 ;
        RECT 413.990 682.400 1997.610 704.800 ;
        RECT 414.400 681.000 1997.610 682.400 ;
        RECT 413.990 670.840 1997.610 681.000 ;
        RECT 413.990 669.440 1997.065 670.840 ;
        RECT 413.990 644.320 1997.610 669.440 ;
        RECT 414.400 642.920 1997.610 644.320 ;
        RECT 413.990 635.480 1997.610 642.920 ;
        RECT 413.990 634.080 1997.065 635.480 ;
        RECT 413.990 606.240 1997.610 634.080 ;
        RECT 414.400 604.840 1997.610 606.240 ;
        RECT 413.990 599.440 1997.610 604.840 ;
        RECT 413.990 598.040 1997.065 599.440 ;
        RECT 413.990 568.160 1997.610 598.040 ;
        RECT 414.400 566.760 1997.610 568.160 ;
        RECT 413.990 564.080 1997.610 566.760 ;
        RECT 413.990 562.680 1997.065 564.080 ;
        RECT 413.990 530.080 1997.610 562.680 ;
        RECT 414.400 528.720 1997.610 530.080 ;
        RECT 414.400 528.680 1997.065 528.720 ;
        RECT 413.990 527.320 1997.065 528.680 ;
        RECT 413.990 514.255 1997.610 527.320 ;
      LAYER met4 ;
        RECT 428.695 520.640 430.640 2101.440 ;
        RECT 433.040 520.640 507.440 2101.440 ;
        RECT 509.840 520.640 1968.640 2101.440 ;
  END
END user_project_wrapper
END LIBRARY

