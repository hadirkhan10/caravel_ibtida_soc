magic
tech sky130A
magscale 1 2
timestamp 1608140683
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 412649 683247 412683 692733
rect 218989 666587 219023 676141
rect 413017 666587 413051 683077
rect 429577 666587 429611 683077
rect 494069 666587 494103 676141
rect 542737 666587 542771 683077
rect 559297 666587 559331 683077
rect 72985 647275 73019 656829
rect 219265 647275 219299 656829
rect 73077 616879 73111 626501
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 412833 601715 412867 608549
rect 429393 601715 429427 608549
rect 542553 601715 542587 608549
rect 559113 601715 559147 608549
rect 72893 589339 72927 598893
rect 219173 589339 219207 598893
rect 413017 589339 413051 598893
rect 429577 589339 429611 598893
rect 542737 589339 542771 598893
rect 559297 589339 559331 598893
rect 8033 579751 8067 589237
rect 137753 579751 137787 589237
rect 154313 579751 154347 589237
rect 284033 579751 284067 589237
rect 347789 579683 347823 589237
rect 364349 579683 364383 589237
rect 477509 579683 477543 589237
rect 72617 569959 72651 579581
rect 137569 569959 137603 579581
rect 218897 569959 218931 579581
rect 347881 563091 347915 569857
rect 364441 563091 364475 569857
rect 477601 563091 477635 569857
rect 494161 563091 494195 569857
rect 72709 550647 72743 560201
rect 137661 550647 137695 560201
rect 218989 550647 219023 560201
rect 412741 550647 412775 560201
rect 429301 550647 429335 560201
rect 542461 550647 542495 560201
rect 559021 550647 559055 560201
rect 8033 543779 8067 550545
rect 154313 543779 154347 550545
rect 284033 543779 284067 550545
rect 72801 521679 72835 524433
rect 137753 521679 137787 524433
rect 219081 521679 219115 524433
rect 135361 147611 135395 154513
rect 135545 131495 135579 143497
rect 143825 128299 143859 143497
rect 135637 106199 135671 122757
rect 135637 89675 135671 104805
rect 135729 77299 135763 85493
rect 143641 77299 143675 86921
rect 135453 57919 135487 60809
rect 143733 48331 143767 57885
rect 135545 11747 135579 27557
rect 201417 3383 201451 3485
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 412649 692733 412683 692767
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 412649 683213 412683 683247
rect 284033 676209 284067 676243
rect 413017 683077 413051 683111
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 413017 666553 413051 666587
rect 429577 683077 429611 683111
rect 542737 683077 542771 683111
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 542737 666553 542771 666587
rect 559297 683077 559331 683111
rect 559297 666553 559331 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 73077 626501 73111 626535
rect 73077 616845 73111 616879
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 412833 608549 412867 608583
rect 412833 601681 412867 601715
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 542553 608549 542587 608583
rect 542553 601681 542587 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 219265 601545 219299 601579
rect 72893 598893 72927 598927
rect 72893 589305 72927 589339
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 413017 598893 413051 598927
rect 413017 589305 413051 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 542737 598893 542771 598927
rect 542737 589305 542771 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 8033 589237 8067 589271
rect 8033 579717 8067 579751
rect 137753 589237 137787 589271
rect 137753 579717 137787 579751
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 284033 589237 284067 589271
rect 284033 579717 284067 579751
rect 347789 589237 347823 589271
rect 347789 579649 347823 579683
rect 364349 589237 364383 589271
rect 364349 579649 364383 579683
rect 477509 589237 477543 589271
rect 477509 579649 477543 579683
rect 72617 579581 72651 579615
rect 72617 569925 72651 569959
rect 137569 579581 137603 579615
rect 137569 569925 137603 569959
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 347881 569857 347915 569891
rect 347881 563057 347915 563091
rect 364441 569857 364475 569891
rect 364441 563057 364475 563091
rect 477601 569857 477635 569891
rect 477601 563057 477635 563091
rect 494161 569857 494195 569891
rect 494161 563057 494195 563091
rect 72709 560201 72743 560235
rect 72709 550613 72743 550647
rect 137661 560201 137695 560235
rect 137661 550613 137695 550647
rect 218989 560201 219023 560235
rect 218989 550613 219023 550647
rect 412741 560201 412775 560235
rect 412741 550613 412775 550647
rect 429301 560201 429335 560235
rect 429301 550613 429335 550647
rect 542461 560201 542495 560235
rect 542461 550613 542495 550647
rect 559021 560201 559055 560235
rect 559021 550613 559055 550647
rect 8033 550545 8067 550579
rect 8033 543745 8067 543779
rect 154313 550545 154347 550579
rect 154313 543745 154347 543779
rect 284033 550545 284067 550579
rect 284033 543745 284067 543779
rect 72801 524433 72835 524467
rect 72801 521645 72835 521679
rect 137753 524433 137787 524467
rect 137753 521645 137787 521679
rect 219081 524433 219115 524467
rect 219081 521645 219115 521679
rect 135361 154513 135395 154547
rect 135361 147577 135395 147611
rect 135545 143497 135579 143531
rect 135545 131461 135579 131495
rect 143825 143497 143859 143531
rect 143825 128265 143859 128299
rect 135637 122757 135671 122791
rect 135637 106165 135671 106199
rect 135637 104805 135671 104839
rect 135637 89641 135671 89675
rect 143641 86921 143675 86955
rect 135729 85493 135763 85527
rect 135729 77265 135763 77299
rect 143641 77265 143675 77299
rect 135453 60809 135487 60843
rect 135453 57885 135487 57919
rect 143733 57885 143767 57919
rect 143733 48297 143767 48331
rect 135545 27557 135579 27591
rect 135545 11713 135579 11747
rect 201417 3485 201451 3519
rect 201417 3349 201451 3383
<< metal1 >>
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 331214 697552 331220 697604
rect 331272 697592 331278 697604
rect 332502 697592 332508 697604
rect 331272 697564 332508 697592
rect 331272 697552 331278 697564
rect 332502 697552 332508 697564
rect 332560 697552 332566 697604
rect 476758 696940 476764 696992
rect 476816 696980 476822 696992
rect 580166 696980 580172 696992
rect 476816 696952 580172 696980
rect 476816 696940 476822 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 347774 692792 347780 692844
rect 347832 692832 347838 692844
rect 348878 692832 348884 692844
rect 347832 692804 348884 692832
rect 347832 692792 347838 692804
rect 348878 692792 348884 692804
rect 348936 692792 348942 692844
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 542538 692724 542544 692776
rect 542596 692764 542602 692776
rect 542722 692764 542728 692776
rect 542596 692736 542728 692764
rect 542596 692724 542602 692736
rect 542722 692724 542728 692736
rect 542780 692724 542786 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 494238 685856 494244 685908
rect 494296 685896 494302 685908
rect 494882 685896 494888 685908
rect 494296 685868 494888 685896
rect 494296 685856 494302 685868
rect 494882 685856 494888 685868
rect 494940 685856 494946 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 429194 684428 429200 684480
rect 429252 684468 429258 684480
rect 429838 684468 429844 684480
rect 429252 684440 429844 684468
rect 429252 684428 429258 684440
rect 429838 684428 429844 684440
rect 429896 684428 429902 684480
rect 558914 684428 558920 684480
rect 558972 684468 558978 684480
rect 559650 684468 559656 684480
rect 558972 684440 559656 684468
rect 558972 684428 558978 684440
rect 559650 684428 559656 684440
rect 559708 684428 559714 684480
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 429194 683068 429200 683120
rect 429252 683108 429258 683120
rect 429565 683111 429623 683117
rect 429565 683108 429577 683111
rect 429252 683080 429577 683108
rect 429252 683068 429258 683080
rect 429565 683077 429577 683080
rect 429611 683077 429623 683111
rect 429565 683071 429623 683077
rect 542354 683068 542360 683120
rect 542412 683108 542418 683120
rect 542725 683111 542783 683117
rect 542725 683108 542737 683111
rect 542412 683080 542737 683108
rect 542412 683068 542418 683080
rect 542725 683077 542737 683080
rect 542771 683077 542783 683111
rect 542725 683071 542783 683077
rect 558914 683068 558920 683120
rect 558972 683108 558978 683120
rect 559285 683111 559343 683117
rect 559285 683108 559297 683111
rect 558972 683080 559297 683108
rect 558972 683068 558978 683080
rect 559285 683077 559297 683080
rect 559331 683077 559343 683111
rect 559285 683071 559343 683077
rect 3326 681708 3332 681760
rect 3384 681748 3390 681760
rect 6178 681748 6184 681760
rect 3384 681720 6184 681748
rect 3384 681708 3390 681720
rect 6178 681708 6184 681720
rect 6236 681708 6242 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 347774 673480 347780 673532
rect 347832 673520 347838 673532
rect 347958 673520 347964 673532
rect 347832 673492 347964 673520
rect 347832 673480 347838 673492
rect 347958 673480 347964 673492
rect 348016 673480 348022 673532
rect 364334 673480 364340 673532
rect 364392 673520 364398 673532
rect 364518 673520 364524 673532
rect 364392 673492 364524 673520
rect 364392 673480 364398 673492
rect 364518 673480 364524 673492
rect 364576 673480 364582 673532
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 483658 673480 483664 673532
rect 483716 673520 483722 673532
rect 580166 673520 580172 673532
rect 483716 673492 580172 673520
rect 483716 673480 483722 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 284018 654100 284024 654152
rect 284076 654140 284082 654152
rect 284202 654140 284208 654152
rect 284076 654112 284208 654140
rect 284076 654100 284082 654112
rect 284202 654100 284208 654112
rect 284260 654100 284266 654152
rect 347774 654100 347780 654152
rect 347832 654140 347838 654152
rect 347958 654140 347964 654152
rect 347832 654112 347964 654140
rect 347832 654100 347838 654112
rect 347958 654100 347964 654112
rect 348016 654100 348022 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 9030 652780 9036 652792
rect 3108 652752 9036 652780
rect 3108 652740 3114 652752
rect 9030 652740 9036 652752
rect 9088 652740 9094 652792
rect 475378 650020 475384 650072
rect 475436 650060 475442 650072
rect 580166 650060 580172 650072
rect 475436 650032 580172 650060
rect 475436 650020 475442 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 72786 637508 72792 637560
rect 72844 637548 72850 637560
rect 72878 637548 72884 637560
rect 72844 637520 72884 637548
rect 72844 637508 72850 637520
rect 72878 637508 72884 637520
rect 72936 637508 72942 637560
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 284018 634788 284024 634840
rect 284076 634828 284082 634840
rect 284202 634828 284208 634840
rect 284076 634800 284208 634828
rect 284076 634788 284082 634800
rect 284202 634788 284208 634800
rect 284260 634788 284266 634840
rect 347774 634788 347780 634840
rect 347832 634828 347838 634840
rect 347958 634828 347964 634840
rect 347832 634800 347964 634828
rect 347832 634788 347838 634800
rect 347958 634788 347964 634800
rect 348016 634788 348022 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 479518 626560 479524 626612
rect 479576 626600 479582 626612
rect 580166 626600 580172 626612
rect 479576 626572 580172 626600
rect 479576 626560 479582 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 73062 626532 73068 626544
rect 73023 626504 73068 626532
rect 73062 626492 73068 626504
rect 73120 626492 73126 626544
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 9030 624384 9036 624436
rect 9088 624424 9094 624436
rect 128998 624424 129004 624436
rect 9088 624396 129004 624424
rect 9088 624384 9094 624396
rect 128998 624384 129004 624396
rect 129056 624384 129062 624436
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 8938 623812 8944 623824
rect 3292 623784 8944 623812
rect 3292 623772 3298 623784
rect 8938 623772 8944 623784
rect 8996 623772 9002 623824
rect 73062 616876 73068 616888
rect 73023 616848 73068 616876
rect 73062 616836 73068 616848
rect 73120 616836 73126 616888
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 284018 615476 284024 615528
rect 284076 615516 284082 615528
rect 284202 615516 284208 615528
rect 284076 615488 284208 615516
rect 284076 615476 284082 615488
rect 284202 615476 284208 615488
rect 284260 615476 284266 615528
rect 347774 615476 347780 615528
rect 347832 615516 347838 615528
rect 347958 615516 347964 615528
rect 347832 615488 347964 615516
rect 347832 615476 347838 615488
rect 347958 615476 347964 615488
rect 348016 615476 348022 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 477494 615476 477500 615528
rect 477552 615516 477558 615528
rect 477678 615516 477684 615528
rect 477552 615488 477684 615516
rect 477552 615476 477558 615488
rect 477678 615476 477684 615488
rect 477736 615476 477742 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 73062 611436 73068 611448
rect 72896 611408 73068 611436
rect 72896 611312 72924 611408
rect 73062 611396 73068 611408
rect 73120 611396 73126 611448
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 72878 611260 72884 611312
rect 72936 611260 72942 611312
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 412818 608580 412824 608592
rect 412779 608552 412824 608580
rect 219253 608543 219311 608549
rect 412818 608540 412824 608552
rect 412876 608540 412882 608592
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 542538 608580 542544 608592
rect 542499 608552 542544 608580
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 471238 603100 471244 603152
rect 471296 603140 471302 603152
rect 580166 603140 580172 603152
rect 471296 603112 580172 603140
rect 471296 603100 471302 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 412821 601715 412879 601721
rect 412821 601681 412833 601715
rect 412867 601712 412879 601715
rect 413002 601712 413008 601724
rect 412867 601684 413008 601712
rect 412867 601681 412879 601684
rect 412821 601675 412879 601681
rect 413002 601672 413008 601684
rect 413060 601672 413066 601724
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 542541 601715 542599 601721
rect 542541 601681 542553 601715
rect 542587 601712 542599 601715
rect 542722 601712 542728 601724
rect 542587 601684 542728 601712
rect 542587 601681 542599 601684
rect 542541 601675 542599 601681
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 72970 601536 72976 601588
rect 73028 601576 73034 601588
rect 73154 601576 73160 601588
rect 73028 601548 73160 601576
rect 73028 601536 73034 601548
rect 73154 601536 73160 601548
rect 73212 601536 73218 601588
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 72881 598927 72939 598933
rect 72881 598893 72893 598927
rect 72927 598924 72939 598927
rect 72970 598924 72976 598936
rect 72927 598896 72976 598924
rect 72927 598893 72939 598896
rect 72881 598887 72939 598893
rect 72970 598884 72976 598896
rect 73028 598884 73034 598936
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 413002 598924 413008 598936
rect 412963 598896 413008 598924
rect 413002 598884 413008 598896
rect 413060 598884 413066 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 542722 598924 542728 598936
rect 542683 598896 542728 598924
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 137738 596164 137744 596216
rect 137796 596204 137802 596216
rect 137922 596204 137928 596216
rect 137796 596176 137928 596204
rect 137796 596164 137802 596176
rect 137922 596164 137928 596176
rect 137980 596164 137986 596216
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 284018 596164 284024 596216
rect 284076 596204 284082 596216
rect 284202 596204 284208 596216
rect 284076 596176 284208 596204
rect 284076 596164 284082 596176
rect 284202 596164 284208 596176
rect 284260 596164 284266 596216
rect 347774 596164 347780 596216
rect 347832 596204 347838 596216
rect 347958 596204 347964 596216
rect 347832 596176 347964 596204
rect 347832 596164 347838 596176
rect 347958 596164 347964 596176
rect 348016 596164 348022 596216
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 477494 596164 477500 596216
rect 477552 596204 477558 596216
rect 477678 596204 477684 596216
rect 477552 596176 477684 596204
rect 477552 596164 477558 596176
rect 477678 596164 477684 596176
rect 477736 596164 477742 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 11698 594844 11704 594856
rect 3384 594816 11704 594844
rect 3384 594804 3390 594816
rect 11698 594804 11704 594816
rect 11756 594804 11762 594856
rect 482278 592016 482284 592068
rect 482336 592056 482342 592068
rect 579890 592056 579896 592068
rect 482336 592028 579896 592056
rect 482336 592016 482342 592028
rect 579890 592016 579896 592028
rect 579948 592016 579954 592068
rect 72878 589336 72884 589348
rect 72839 589308 72884 589336
rect 72878 589296 72884 589308
rect 72936 589296 72942 589348
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 413005 589339 413063 589345
rect 413005 589305 413017 589339
rect 413051 589336 413063 589339
rect 413094 589336 413100 589348
rect 413051 589308 413100 589336
rect 413051 589305 413063 589308
rect 413005 589299 413063 589305
rect 413094 589296 413100 589308
rect 413152 589296 413158 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 542725 589339 542783 589345
rect 542725 589305 542737 589339
rect 542771 589336 542783 589339
rect 542814 589336 542820 589348
rect 542771 589308 542820 589336
rect 542771 589305 542783 589308
rect 542725 589299 542783 589305
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 8018 589268 8024 589280
rect 7979 589240 8024 589268
rect 8018 589228 8024 589240
rect 8076 589228 8082 589280
rect 137738 589268 137744 589280
rect 137699 589240 137744 589268
rect 137738 589228 137744 589240
rect 137796 589228 137802 589280
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 284018 589268 284024 589280
rect 283979 589240 284024 589268
rect 284018 589228 284024 589240
rect 284076 589228 284082 589280
rect 347777 589271 347835 589277
rect 347777 589237 347789 589271
rect 347823 589268 347835 589271
rect 347866 589268 347872 589280
rect 347823 589240 347872 589268
rect 347823 589237 347835 589240
rect 347777 589231 347835 589237
rect 347866 589228 347872 589240
rect 347924 589228 347930 589280
rect 364337 589271 364395 589277
rect 364337 589237 364349 589271
rect 364383 589268 364395 589271
rect 364426 589268 364432 589280
rect 364383 589240 364432 589268
rect 364383 589237 364395 589240
rect 364337 589231 364395 589237
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 477497 589271 477555 589277
rect 477497 589237 477509 589271
rect 477543 589268 477555 589271
rect 477586 589268 477592 589280
rect 477543 589240 477592 589268
rect 477543 589237 477555 589240
rect 477497 589231 477555 589237
rect 477586 589228 477592 589240
rect 477644 589228 477650 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 413094 582468 413100 582480
rect 413020 582440 413100 582468
rect 72694 582360 72700 582412
rect 72752 582400 72758 582412
rect 72878 582400 72884 582412
rect 72752 582372 72884 582400
rect 72752 582360 72758 582372
rect 72878 582360 72884 582372
rect 72936 582360 72942 582412
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 413020 582344 413048 582440
rect 413094 582428 413100 582440
rect 413152 582428 413158 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 413002 582292 413008 582344
rect 413060 582292 413066 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 8018 579748 8024 579760
rect 7979 579720 8024 579748
rect 8018 579708 8024 579720
rect 8076 579708 8082 579760
rect 137738 579748 137744 579760
rect 137699 579720 137744 579748
rect 137738 579708 137744 579720
rect 137796 579708 137802 579760
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 284018 579748 284024 579760
rect 283979 579720 284024 579748
rect 284018 579708 284024 579720
rect 284076 579708 284082 579760
rect 347774 579640 347780 579692
rect 347832 579680 347838 579692
rect 364334 579680 364340 579692
rect 347832 579652 347877 579680
rect 364295 579652 364340 579680
rect 347832 579640 347838 579652
rect 364334 579640 364340 579652
rect 364392 579640 364398 579692
rect 477494 579680 477500 579692
rect 477455 579652 477500 579680
rect 477494 579640 477500 579652
rect 477552 579640 477558 579692
rect 489178 579640 489184 579692
rect 489236 579680 489242 579692
rect 580166 579680 580172 579692
rect 489236 579652 580172 579680
rect 489236 579640 489242 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 7926 579572 7932 579624
rect 7984 579612 7990 579624
rect 8110 579612 8116 579624
rect 7984 579584 8116 579612
rect 7984 579572 7990 579584
rect 8110 579572 8116 579584
rect 8168 579572 8174 579624
rect 72605 579615 72663 579621
rect 72605 579581 72617 579615
rect 72651 579612 72663 579615
rect 72694 579612 72700 579624
rect 72651 579584 72700 579612
rect 72651 579581 72663 579584
rect 72605 579575 72663 579581
rect 72694 579572 72700 579584
rect 72752 579572 72758 579624
rect 137557 579615 137615 579621
rect 137557 579581 137569 579615
rect 137603 579612 137615 579615
rect 137646 579612 137652 579624
rect 137603 579584 137652 579612
rect 137603 579581 137615 579584
rect 137557 579575 137615 579581
rect 137646 579572 137652 579584
rect 137704 579572 137710 579624
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 283926 579572 283932 579624
rect 283984 579612 283990 579624
rect 284110 579612 284116 579624
rect 283984 579584 284116 579612
rect 283984 579572 283990 579584
rect 284110 579572 284116 579584
rect 284168 579572 284174 579624
rect 72602 569956 72608 569968
rect 72563 569928 72608 569956
rect 72602 569916 72608 569928
rect 72660 569916 72666 569968
rect 137554 569956 137560 569968
rect 137515 569928 137560 569956
rect 137554 569916 137560 569928
rect 137612 569916 137618 569968
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 347866 569888 347872 569900
rect 347827 569860 347872 569888
rect 347866 569848 347872 569860
rect 347924 569848 347930 569900
rect 364426 569888 364432 569900
rect 364387 569860 364432 569888
rect 364426 569848 364432 569860
rect 364484 569848 364490 569900
rect 477586 569888 477592 569900
rect 477547 569860 477592 569888
rect 477586 569848 477592 569860
rect 477644 569848 477650 569900
rect 494146 569888 494152 569900
rect 494107 569860 494152 569888
rect 494146 569848 494152 569860
rect 494204 569848 494210 569900
rect 4062 567264 4068 567316
rect 4120 567304 4126 567316
rect 10318 567304 10324 567316
rect 4120 567276 10324 567304
rect 4120 567264 4126 567276
rect 10318 567264 10324 567276
rect 10376 567264 10382 567316
rect 412726 563116 412732 563168
rect 412784 563116 412790 563168
rect 429286 563116 429292 563168
rect 429344 563116 429350 563168
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 72602 563048 72608 563100
rect 72660 563048 72666 563100
rect 137554 563048 137560 563100
rect 137612 563048 137618 563100
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 347869 563091 347927 563097
rect 347869 563057 347881 563091
rect 347915 563088 347927 563091
rect 348050 563088 348056 563100
rect 347915 563060 348056 563088
rect 347915 563057 347927 563060
rect 347869 563051 347927 563057
rect 348050 563048 348056 563060
rect 348108 563048 348114 563100
rect 364429 563091 364487 563097
rect 364429 563057 364441 563091
rect 364475 563088 364487 563091
rect 364610 563088 364616 563100
rect 364475 563060 364616 563088
rect 364475 563057 364487 563060
rect 364429 563051 364487 563057
rect 364610 563048 364616 563060
rect 364668 563048 364674 563100
rect 7926 562912 7932 562964
rect 7984 562952 7990 562964
rect 8110 562952 8116 562964
rect 7984 562924 8116 562952
rect 7984 562912 7990 562924
rect 8110 562912 8116 562924
rect 8168 562912 8174 562964
rect 72620 562952 72648 563048
rect 72694 562952 72700 562964
rect 72620 562924 72700 562952
rect 72694 562912 72700 562924
rect 72752 562912 72758 562964
rect 137572 562952 137600 563048
rect 137646 562952 137652 562964
rect 137572 562924 137652 562952
rect 137646 562912 137652 562924
rect 137704 562912 137710 562964
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 412744 563032 412772 563116
rect 429304 563032 429332 563116
rect 477589 563091 477647 563097
rect 477589 563057 477601 563091
rect 477635 563088 477647 563091
rect 477770 563088 477776 563100
rect 477635 563060 477776 563088
rect 477635 563057 477647 563060
rect 477589 563051 477647 563057
rect 477770 563048 477776 563060
rect 477828 563048 477834 563100
rect 494149 563091 494207 563097
rect 494149 563057 494161 563091
rect 494195 563088 494207 563091
rect 494330 563088 494336 563100
rect 494195 563060 494336 563088
rect 494195 563057 494207 563060
rect 494149 563051 494207 563057
rect 494330 563048 494336 563060
rect 494388 563048 494394 563100
rect 542464 563032 542492 563116
rect 559024 563032 559052 563116
rect 412726 562980 412732 563032
rect 412784 562980 412790 563032
rect 429286 562980 429292 563032
rect 429344 562980 429350 563032
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 283926 562912 283932 562964
rect 283984 562952 283990 562964
rect 284110 562952 284116 562964
rect 283984 562924 284116 562952
rect 283984 562912 283990 562924
rect 284110 562912 284116 562924
rect 284168 562912 284174 562964
rect 72694 560232 72700 560244
rect 72655 560204 72700 560232
rect 72694 560192 72700 560204
rect 72752 560192 72758 560244
rect 137646 560232 137652 560244
rect 137607 560204 137652 560232
rect 137646 560192 137652 560204
rect 137704 560192 137710 560244
rect 218974 560232 218980 560244
rect 218935 560204 218980 560232
rect 218974 560192 218980 560204
rect 219032 560192 219038 560244
rect 412726 560232 412732 560244
rect 412687 560204 412732 560232
rect 412726 560192 412732 560204
rect 412784 560192 412790 560244
rect 429286 560232 429292 560244
rect 429247 560204 429292 560232
rect 429286 560192 429292 560204
rect 429344 560192 429350 560244
rect 542446 560232 542452 560244
rect 542407 560204 542452 560232
rect 542446 560192 542452 560204
rect 542504 560192 542510 560244
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 467098 556180 467104 556232
rect 467156 556220 467162 556232
rect 580166 556220 580172 556232
rect 467156 556192 580172 556220
rect 467156 556180 467162 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 72697 550647 72755 550653
rect 72697 550613 72709 550647
rect 72743 550644 72755 550647
rect 72878 550644 72884 550656
rect 72743 550616 72884 550644
rect 72743 550613 72755 550616
rect 72697 550607 72755 550613
rect 72878 550604 72884 550616
rect 72936 550604 72942 550656
rect 137649 550647 137707 550653
rect 137649 550613 137661 550647
rect 137695 550644 137707 550647
rect 137830 550644 137836 550656
rect 137695 550616 137836 550644
rect 137695 550613 137707 550616
rect 137649 550607 137707 550613
rect 137830 550604 137836 550616
rect 137888 550604 137894 550656
rect 218977 550647 219035 550653
rect 218977 550613 218989 550647
rect 219023 550644 219035 550647
rect 219158 550644 219164 550656
rect 219023 550616 219164 550644
rect 219023 550613 219035 550616
rect 218977 550607 219035 550613
rect 219158 550604 219164 550616
rect 219216 550604 219222 550656
rect 347866 550604 347872 550656
rect 347924 550644 347930 550656
rect 348142 550644 348148 550656
rect 347924 550616 348148 550644
rect 347924 550604 347930 550616
rect 348142 550604 348148 550616
rect 348200 550604 348206 550656
rect 364426 550604 364432 550656
rect 364484 550644 364490 550656
rect 364702 550644 364708 550656
rect 364484 550616 364708 550644
rect 364484 550604 364490 550616
rect 364702 550604 364708 550616
rect 364760 550604 364766 550656
rect 412729 550647 412787 550653
rect 412729 550613 412741 550647
rect 412775 550644 412787 550647
rect 412910 550644 412916 550656
rect 412775 550616 412916 550644
rect 412775 550613 412787 550616
rect 412729 550607 412787 550613
rect 412910 550604 412916 550616
rect 412968 550604 412974 550656
rect 429289 550647 429347 550653
rect 429289 550613 429301 550647
rect 429335 550644 429347 550647
rect 429470 550644 429476 550656
rect 429335 550616 429476 550644
rect 429335 550613 429347 550616
rect 429289 550607 429347 550613
rect 429470 550604 429476 550616
rect 429528 550604 429534 550656
rect 477586 550604 477592 550656
rect 477644 550644 477650 550656
rect 477862 550644 477868 550656
rect 477644 550616 477868 550644
rect 477644 550604 477650 550616
rect 477862 550604 477868 550616
rect 477920 550604 477926 550656
rect 494146 550604 494152 550656
rect 494204 550644 494210 550656
rect 494422 550644 494428 550656
rect 494204 550616 494428 550644
rect 494204 550604 494210 550616
rect 494422 550604 494428 550616
rect 494480 550604 494486 550656
rect 542449 550647 542507 550653
rect 542449 550613 542461 550647
rect 542495 550644 542507 550647
rect 542630 550644 542636 550656
rect 542495 550616 542636 550644
rect 542495 550613 542507 550616
rect 542449 550607 542507 550613
rect 542630 550604 542636 550616
rect 542688 550604 542694 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559190 550644 559196 550656
rect 559055 550616 559196 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559190 550604 559196 550616
rect 559248 550604 559254 550656
rect 8018 550576 8024 550588
rect 7979 550548 8024 550576
rect 8018 550536 8024 550548
rect 8076 550536 8082 550588
rect 154298 550576 154304 550588
rect 154259 550548 154304 550576
rect 154298 550536 154304 550548
rect 154356 550536 154362 550588
rect 284018 550576 284024 550588
rect 283979 550548 284024 550576
rect 284018 550536 284024 550548
rect 284076 550536 284082 550588
rect 480898 545096 480904 545148
rect 480956 545136 480962 545148
rect 579890 545136 579896 545148
rect 480956 545108 579896 545136
rect 480956 545096 480962 545108
rect 579890 545096 579896 545108
rect 579948 545096 579954 545148
rect 348142 543844 348148 543856
rect 348068 543816 348148 543844
rect 8021 543779 8079 543785
rect 8021 543745 8033 543779
rect 8067 543776 8079 543779
rect 8202 543776 8208 543788
rect 8067 543748 8208 543776
rect 8067 543745 8079 543748
rect 8021 543739 8079 543745
rect 8202 543736 8208 543748
rect 8260 543736 8266 543788
rect 154301 543779 154359 543785
rect 154301 543745 154313 543779
rect 154347 543776 154359 543779
rect 154482 543776 154488 543788
rect 154347 543748 154488 543776
rect 154347 543745 154359 543748
rect 154301 543739 154359 543745
rect 154482 543736 154488 543748
rect 154540 543736 154546 543788
rect 284021 543779 284079 543785
rect 284021 543745 284033 543779
rect 284067 543776 284079 543779
rect 284202 543776 284208 543788
rect 284067 543748 284208 543776
rect 284067 543745 284079 543748
rect 284021 543739 284079 543745
rect 284202 543736 284208 543748
rect 284260 543736 284266 543788
rect 348068 543720 348096 543816
rect 348142 543804 348148 543816
rect 348200 543804 348206 543856
rect 364702 543844 364708 543856
rect 364628 543816 364708 543844
rect 364628 543720 364656 543816
rect 364702 543804 364708 543816
rect 364760 543804 364766 543856
rect 477862 543844 477868 543856
rect 477788 543816 477868 543844
rect 477788 543720 477816 543816
rect 477862 543804 477868 543816
rect 477920 543804 477926 543856
rect 494422 543844 494428 543856
rect 494348 543816 494428 543844
rect 494348 543720 494376 543816
rect 494422 543804 494428 543816
rect 494480 543804 494486 543856
rect 348050 543668 348056 543720
rect 348108 543668 348114 543720
rect 364610 543668 364616 543720
rect 364668 543668 364674 543720
rect 477770 543668 477776 543720
rect 477828 543668 477834 543720
rect 494330 543668 494336 543720
rect 494388 543668 494394 543720
rect 72694 543600 72700 543652
rect 72752 543640 72758 543652
rect 72878 543640 72884 543652
rect 72752 543612 72884 543640
rect 72752 543600 72758 543612
rect 72878 543600 72884 543612
rect 72936 543600 72942 543652
rect 137646 543600 137652 543652
rect 137704 543640 137710 543652
rect 137830 543640 137836 543652
rect 137704 543612 137836 543640
rect 137704 543600 137710 543612
rect 137830 543600 137836 543612
rect 137888 543600 137894 543652
rect 218974 543600 218980 543652
rect 219032 543640 219038 543652
rect 219158 543640 219164 543652
rect 219032 543612 219164 543640
rect 219032 543600 219038 543612
rect 219158 543600 219164 543612
rect 219216 543600 219222 543652
rect 412726 543600 412732 543652
rect 412784 543640 412790 543652
rect 412910 543640 412916 543652
rect 412784 543612 412916 543640
rect 412784 543600 412790 543612
rect 412910 543600 412916 543612
rect 412968 543600 412974 543652
rect 429286 543600 429292 543652
rect 429344 543640 429350 543652
rect 429470 543640 429476 543652
rect 429344 543612 429476 543640
rect 429344 543600 429350 543612
rect 429470 543600 429476 543612
rect 429528 543600 429534 543652
rect 542446 543600 542452 543652
rect 542504 543640 542510 543652
rect 542630 543640 542636 543652
rect 542504 543612 542636 543640
rect 542504 543600 542510 543612
rect 542630 543600 542636 543612
rect 542688 543600 542694 543652
rect 559006 543600 559012 543652
rect 559064 543640 559070 543652
rect 559190 543640 559196 543652
rect 559064 543612 559196 543640
rect 559064 543600 559070 543612
rect 559190 543600 559196 543612
rect 559248 543600 559254 543652
rect 72694 534012 72700 534064
rect 72752 534052 72758 534064
rect 72878 534052 72884 534064
rect 72752 534024 72884 534052
rect 72752 534012 72758 534024
rect 72878 534012 72884 534024
rect 72936 534012 72942 534064
rect 137646 534012 137652 534064
rect 137704 534052 137710 534064
rect 137830 534052 137836 534064
rect 137704 534024 137836 534052
rect 137704 534012 137710 534024
rect 137830 534012 137836 534024
rect 137888 534012 137894 534064
rect 218974 534012 218980 534064
rect 219032 534052 219038 534064
rect 219158 534052 219164 534064
rect 219032 534024 219164 534052
rect 219032 534012 219038 534024
rect 219158 534012 219164 534024
rect 219216 534012 219222 534064
rect 485038 532720 485044 532772
rect 485096 532760 485102 532772
rect 580166 532760 580172 532772
rect 485096 532732 580172 532760
rect 485096 532720 485102 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 154206 531292 154212 531344
rect 154264 531332 154270 531344
rect 154298 531332 154304 531344
rect 154264 531304 154304 531332
rect 154264 531292 154270 531304
rect 154298 531292 154304 531304
rect 154356 531292 154362 531344
rect 347866 531292 347872 531344
rect 347924 531332 347930 531344
rect 348142 531332 348148 531344
rect 347924 531304 348148 531332
rect 347924 531292 347930 531304
rect 348142 531292 348148 531304
rect 348200 531292 348206 531344
rect 364426 531292 364432 531344
rect 364484 531332 364490 531344
rect 364702 531332 364708 531344
rect 364484 531304 364708 531332
rect 364484 531292 364490 531304
rect 364702 531292 364708 531304
rect 364760 531292 364766 531344
rect 477586 531292 477592 531344
rect 477644 531332 477650 531344
rect 477862 531332 477868 531344
rect 477644 531304 477868 531332
rect 477644 531292 477650 531304
rect 477862 531292 477868 531304
rect 477920 531292 477926 531344
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 72786 524464 72792 524476
rect 72747 524436 72792 524464
rect 72786 524424 72792 524436
rect 72844 524424 72850 524476
rect 137738 524464 137744 524476
rect 137699 524436 137744 524464
rect 137738 524424 137744 524436
rect 137796 524424 137802 524476
rect 154298 524424 154304 524476
rect 154356 524424 154362 524476
rect 219066 524464 219072 524476
rect 219027 524436 219072 524464
rect 219066 524424 219072 524436
rect 219124 524424 219130 524476
rect 8110 524288 8116 524340
rect 8168 524328 8174 524340
rect 8294 524328 8300 524340
rect 8168 524300 8300 524328
rect 8168 524288 8174 524300
rect 8294 524288 8300 524300
rect 8352 524288 8358 524340
rect 154316 524328 154344 524424
rect 154390 524328 154396 524340
rect 154316 524300 154396 524328
rect 154390 524288 154396 524300
rect 154448 524288 154454 524340
rect 284110 524288 284116 524340
rect 284168 524328 284174 524340
rect 284294 524328 284300 524340
rect 284168 524300 284300 524328
rect 284168 524288 284174 524300
rect 284294 524288 284300 524300
rect 284352 524288 284358 524340
rect 72786 521676 72792 521688
rect 72747 521648 72792 521676
rect 72786 521636 72792 521648
rect 72844 521636 72850 521688
rect 137738 521676 137744 521688
rect 137699 521648 137744 521676
rect 137738 521636 137744 521648
rect 137796 521636 137802 521688
rect 219066 521676 219072 521688
rect 219027 521648 219072 521676
rect 219066 521636 219072 521648
rect 219124 521636 219130 521688
rect 347958 521636 347964 521688
rect 348016 521676 348022 521688
rect 348142 521676 348148 521688
rect 348016 521648 348148 521676
rect 348016 521636 348022 521648
rect 348142 521636 348148 521648
rect 348200 521636 348206 521688
rect 364518 521636 364524 521688
rect 364576 521676 364582 521688
rect 364702 521676 364708 521688
rect 364576 521648 364708 521676
rect 364576 521636 364582 521648
rect 364702 521636 364708 521648
rect 364760 521636 364766 521688
rect 477678 521636 477684 521688
rect 477736 521676 477742 521688
rect 477862 521676 477868 521688
rect 477736 521648 477868 521676
rect 477736 521636 477742 521648
rect 477862 521636 477868 521648
rect 477920 521636 477926 521688
rect 494238 521636 494244 521688
rect 494296 521676 494302 521688
rect 494422 521676 494428 521688
rect 494296 521648 494428 521676
rect 494296 521636 494302 521648
rect 494422 521636 494428 521648
rect 494480 521636 494486 521688
rect 284110 516060 284116 516112
rect 284168 516100 284174 516112
rect 291102 516100 291108 516112
rect 284168 516072 291108 516100
rect 284168 516060 284174 516072
rect 291102 516060 291108 516072
rect 291160 516060 291166 516112
rect 106182 515720 106188 515772
rect 106240 515760 106246 515772
rect 196802 515760 196808 515772
rect 106240 515732 196808 515760
rect 106240 515720 106246 515732
rect 196802 515720 196808 515732
rect 196860 515720 196866 515772
rect 385494 515720 385500 515772
rect 385552 515760 385558 515772
rect 462314 515760 462320 515772
rect 385552 515732 462320 515760
rect 385552 515720 385558 515732
rect 462314 515720 462320 515732
rect 462372 515720 462378 515772
rect 89622 515652 89628 515704
rect 89680 515692 89686 515704
rect 185026 515692 185032 515704
rect 89680 515664 185032 515692
rect 89680 515652 89686 515664
rect 185026 515652 185032 515664
rect 185084 515652 185090 515704
rect 397270 515652 397276 515704
rect 397328 515692 397334 515704
rect 477678 515692 477684 515704
rect 397328 515664 477684 515692
rect 397328 515652 397334 515664
rect 477678 515652 477684 515664
rect 477736 515652 477742 515704
rect 72786 515584 72792 515636
rect 72844 515624 72850 515636
rect 173250 515624 173256 515636
rect 72844 515596 173256 515624
rect 72844 515584 72850 515596
rect 173250 515584 173256 515596
rect 173308 515584 173314 515636
rect 202782 515584 202788 515636
rect 202840 515624 202846 515636
rect 243998 515624 244004 515636
rect 202840 515596 244004 515624
rect 202840 515584 202846 515596
rect 243998 515584 244004 515596
rect 244056 515584 244062 515636
rect 409046 515584 409052 515636
rect 409104 515624 409110 515636
rect 494238 515624 494244 515636
rect 409104 515596 494244 515624
rect 409104 515584 409110 515596
rect 494238 515584 494244 515596
rect 494296 515584 494302 515636
rect 41322 515516 41328 515568
rect 41380 515556 41386 515568
rect 161474 515556 161480 515568
rect 41380 515528 161480 515556
rect 41380 515516 41386 515528
rect 161474 515516 161480 515528
rect 161532 515516 161538 515568
rect 171042 515516 171048 515568
rect 171100 515556 171106 515568
rect 232222 515556 232228 515568
rect 171100 515528 232228 515556
rect 171100 515516 171106 515528
rect 232222 515516 232228 515528
rect 232280 515516 232286 515568
rect 350074 515516 350080 515568
rect 350132 515556 350138 515568
rect 397454 515556 397460 515568
rect 350132 515528 397460 515556
rect 350132 515516 350138 515528
rect 397454 515516 397460 515528
rect 397512 515516 397518 515568
rect 420822 515516 420828 515568
rect 420880 515556 420886 515568
rect 527174 515556 527180 515568
rect 420880 515528 527180 515556
rect 420880 515516 420886 515528
rect 527174 515516 527180 515528
rect 527232 515516 527238 515568
rect 24762 515448 24768 515500
rect 24820 515488 24826 515500
rect 149698 515488 149704 515500
rect 24820 515460 149704 515488
rect 24820 515448 24826 515460
rect 149698 515448 149704 515460
rect 149756 515448 149762 515500
rect 154390 515448 154396 515500
rect 154448 515488 154454 515500
rect 220446 515488 220452 515500
rect 154448 515460 220452 515488
rect 154448 515448 154454 515460
rect 220446 515448 220452 515460
rect 220504 515448 220510 515500
rect 235902 515448 235908 515500
rect 235960 515488 235966 515500
rect 267550 515488 267556 515500
rect 235960 515460 267556 515488
rect 235960 515448 235966 515460
rect 267550 515448 267556 515460
rect 267608 515448 267614 515500
rect 326522 515448 326528 515500
rect 326580 515488 326586 515500
rect 347958 515488 347964 515500
rect 326580 515460 347964 515488
rect 326580 515448 326586 515460
rect 347958 515448 347964 515460
rect 348016 515448 348022 515500
rect 361850 515448 361856 515500
rect 361908 515488 361914 515500
rect 412910 515488 412916 515500
rect 361908 515460 412916 515488
rect 361908 515448 361914 515460
rect 412910 515448 412916 515460
rect 412968 515448 412974 515500
rect 432598 515448 432604 515500
rect 432656 515488 432662 515500
rect 542630 515488 542636 515500
rect 432656 515460 542636 515488
rect 432656 515448 432662 515460
rect 542630 515448 542636 515460
rect 542688 515448 542694 515500
rect 8110 515380 8116 515432
rect 8168 515420 8174 515432
rect 137922 515420 137928 515432
rect 8168 515392 137928 515420
rect 8168 515380 8174 515392
rect 137922 515380 137928 515392
rect 137980 515380 137986 515432
rect 138014 515380 138020 515432
rect 138072 515420 138078 515432
rect 208578 515420 208584 515432
rect 138072 515392 208584 515420
rect 138072 515380 138078 515392
rect 208578 515380 208584 515392
rect 208636 515380 208642 515432
rect 219066 515380 219072 515432
rect 219124 515420 219130 515432
rect 255774 515420 255780 515432
rect 219124 515392 255780 515420
rect 219124 515380 219130 515392
rect 255774 515380 255780 515392
rect 255832 515380 255838 515432
rect 267642 515380 267648 515432
rect 267700 515420 267706 515432
rect 279326 515420 279332 515432
rect 267700 515392 279332 515420
rect 267700 515380 267706 515392
rect 279326 515380 279332 515392
rect 279384 515380 279390 515432
rect 314746 515380 314752 515432
rect 314804 515420 314810 515432
rect 331214 515420 331220 515432
rect 314804 515392 331220 515420
rect 314804 515380 314810 515392
rect 331214 515380 331220 515392
rect 331272 515380 331278 515432
rect 338298 515380 338304 515432
rect 338356 515420 338362 515432
rect 364518 515420 364524 515432
rect 338356 515392 364524 515420
rect 338356 515380 338362 515392
rect 364518 515380 364524 515392
rect 364576 515380 364582 515432
rect 373626 515380 373632 515432
rect 373684 515420 373690 515432
rect 429470 515420 429476 515432
rect 373684 515392 429476 515420
rect 373684 515380 373690 515392
rect 429470 515380 429476 515392
rect 429528 515380 429534 515432
rect 444374 515380 444380 515432
rect 444432 515420 444438 515432
rect 559190 515420 559196 515432
rect 444432 515392 559196 515420
rect 444432 515380 444438 515392
rect 559190 515380 559196 515392
rect 559248 515380 559254 515432
rect 300762 514836 300768 514888
rect 300820 514876 300826 514888
rect 302970 514876 302976 514888
rect 300820 514848 302976 514876
rect 300820 514836 300826 514848
rect 302970 514836 302976 514848
rect 303028 514836 303034 514888
rect 3234 509260 3240 509312
rect 3292 509300 3298 509312
rect 7558 509300 7564 509312
rect 3292 509272 7564 509300
rect 3292 509260 3298 509272
rect 7558 509260 7564 509272
rect 7616 509260 7622 509312
rect 462958 509260 462964 509312
rect 463016 509300 463022 509312
rect 580166 509300 580172 509312
rect 463016 509272 580172 509300
rect 463016 509260 463022 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 6178 509192 6184 509244
rect 6236 509232 6242 509244
rect 128354 509232 128360 509244
rect 6236 509204 128360 509232
rect 6236 509192 6242 509204
rect 128354 509192 128360 509204
rect 128412 509192 128418 509244
rect 453206 509192 453212 509244
rect 453264 509232 453270 509244
rect 476758 509232 476764 509244
rect 453264 509204 476764 509232
rect 453264 509192 453270 509204
rect 476758 509192 476764 509204
rect 476816 509192 476822 509244
rect 3418 502256 3424 502308
rect 3476 502296 3482 502308
rect 128354 502296 128360 502308
rect 3476 502268 128360 502296
rect 3476 502256 3482 502268
rect 128354 502256 128360 502268
rect 128412 502256 128418 502308
rect 453390 502256 453396 502308
rect 453448 502296 453454 502308
rect 580258 502296 580264 502308
rect 453448 502268 580264 502296
rect 453448 502256 453454 502268
rect 580258 502256 580264 502268
rect 580316 502256 580322 502308
rect 460198 498176 460204 498228
rect 460256 498216 460262 498228
rect 580166 498216 580172 498228
rect 460256 498188 580172 498216
rect 460256 498176 460262 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 453942 495388 453948 495440
rect 454000 495428 454006 495440
rect 483658 495428 483664 495440
rect 454000 495400 483664 495428
rect 454000 495388 454006 495400
rect 483658 495388 483664 495400
rect 483716 495388 483722 495440
rect 453758 488452 453764 488504
rect 453816 488492 453822 488504
rect 475378 488492 475384 488504
rect 453816 488464 475384 488492
rect 453816 488452 453822 488464
rect 475378 488452 475384 488464
rect 475436 488452 475442 488504
rect 456058 485800 456064 485852
rect 456116 485840 456122 485852
rect 580166 485840 580172 485852
rect 456116 485812 580172 485840
rect 456116 485800 456122 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 8938 485732 8944 485784
rect 8996 485772 9002 485784
rect 128354 485772 128360 485784
rect 8996 485744 128360 485772
rect 8996 485732 9002 485744
rect 128354 485732 128360 485744
rect 128412 485732 128418 485784
rect 453758 481584 453764 481636
rect 453816 481624 453822 481636
rect 580350 481624 580356 481636
rect 453816 481596 580356 481624
rect 453816 481584 453822 481596
rect 580350 481584 580356 481596
rect 580408 481584 580414 481636
rect 3510 478796 3516 478848
rect 3568 478836 3574 478848
rect 128354 478836 128360 478848
rect 3568 478808 128360 478836
rect 3568 478796 3574 478808
rect 128354 478796 128360 478808
rect 128412 478796 128418 478848
rect 453942 473288 453948 473340
rect 454000 473328 454006 473340
rect 479518 473328 479524 473340
rect 454000 473300 479524 473328
rect 454000 473288 454006 473300
rect 479518 473288 479524 473300
rect 479576 473288 479582 473340
rect 11698 470500 11704 470552
rect 11756 470540 11762 470552
rect 128354 470540 128360 470552
rect 11756 470512 128360 470540
rect 11756 470500 11762 470512
rect 128354 470500 128360 470512
rect 128412 470500 128418 470552
rect 452746 466352 452752 466404
rect 452804 466392 452810 466404
rect 471238 466392 471244 466404
rect 452804 466364 471244 466392
rect 452804 466352 452810 466364
rect 471238 466352 471244 466364
rect 471296 466352 471302 466404
rect 10318 463632 10324 463684
rect 10376 463672 10382 463684
rect 128354 463672 128360 463684
rect 10376 463644 128360 463672
rect 10376 463632 10382 463644
rect 128354 463632 128360 463644
rect 128412 463632 128418 463684
rect 542998 462340 543004 462392
rect 543056 462380 543062 462392
rect 580166 462380 580172 462392
rect 543056 462352 580172 462380
rect 543056 462340 543062 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 453390 459484 453396 459536
rect 453448 459524 453454 459536
rect 482278 459524 482284 459536
rect 453448 459496 482284 459524
rect 453448 459484 453454 459496
rect 482278 459484 482284 459496
rect 482336 459484 482342 459536
rect 3602 455336 3608 455388
rect 3660 455376 3666 455388
rect 128354 455376 128360 455388
rect 3660 455348 128360 455376
rect 3660 455336 3666 455348
rect 128354 455336 128360 455348
rect 128412 455336 128418 455388
rect 453942 452548 453948 452600
rect 454000 452588 454006 452600
rect 489178 452588 489184 452600
rect 454000 452560 489184 452588
rect 454000 452548 454006 452560
rect 489178 452548 489184 452560
rect 489236 452548 489242 452600
rect 3694 448468 3700 448520
rect 3752 448508 3758 448520
rect 128354 448508 128360 448520
rect 3752 448480 128360 448508
rect 3752 448468 3758 448480
rect 128354 448468 128360 448480
rect 128412 448468 128418 448520
rect 453666 445680 453672 445732
rect 453724 445720 453730 445732
rect 467098 445720 467104 445732
rect 453724 445692 467104 445720
rect 453724 445680 453730 445692
rect 467098 445680 467104 445692
rect 467156 445680 467162 445732
rect 7558 440172 7564 440224
rect 7616 440212 7622 440224
rect 128354 440212 128360 440224
rect 7616 440184 128360 440212
rect 7616 440172 7622 440184
rect 128354 440172 128360 440184
rect 128412 440172 128418 440224
rect 453298 438880 453304 438932
rect 453356 438920 453362 438932
rect 579890 438920 579896 438932
rect 453356 438892 579896 438920
rect 453356 438880 453362 438892
rect 579890 438880 579896 438892
rect 579948 438880 579954 438932
rect 453758 438812 453764 438864
rect 453816 438852 453822 438864
rect 480898 438852 480904 438864
rect 453816 438824 480904 438852
rect 453816 438812 453822 438824
rect 480898 438812 480904 438824
rect 480956 438812 480962 438864
rect 3418 433236 3424 433288
rect 3476 433276 3482 433288
rect 128354 433276 128360 433288
rect 3476 433248 128360 433276
rect 3476 433236 3482 433248
rect 128354 433236 128360 433248
rect 128412 433236 128418 433288
rect 453942 430516 453948 430568
rect 454000 430556 454006 430568
rect 485038 430556 485044 430568
rect 454000 430528 485044 430556
rect 454000 430516 454006 430528
rect 485038 430516 485044 430528
rect 485096 430516 485102 430568
rect 3786 425008 3792 425060
rect 3844 425048 3850 425060
rect 128354 425048 128360 425060
rect 3844 425020 128360 425048
rect 3844 425008 3850 425020
rect 128354 425008 128360 425020
rect 128412 425008 128418 425060
rect 453942 423580 453948 423632
rect 454000 423620 454006 423632
rect 462958 423620 462964 423632
rect 454000 423592 462964 423620
rect 454000 423580 454006 423592
rect 462958 423580 462964 423592
rect 463016 423580 463022 423632
rect 3510 418072 3516 418124
rect 3568 418112 3574 418124
rect 128354 418112 128360 418124
rect 3568 418084 128360 418112
rect 3568 418072 3574 418084
rect 128354 418072 128360 418084
rect 128412 418072 128418 418124
rect 453942 416372 453948 416424
rect 454000 416412 454006 416424
rect 460198 416412 460204 416424
rect 454000 416384 460204 416412
rect 454000 416372 454006 416384
rect 460198 416372 460204 416384
rect 460256 416372 460262 416424
rect 3602 409776 3608 409828
rect 3660 409816 3666 409828
rect 128354 409816 128360 409828
rect 3660 409788 128360 409816
rect 3660 409776 3666 409788
rect 128354 409776 128360 409788
rect 128412 409776 128418 409828
rect 453390 409368 453396 409420
rect 453448 409408 453454 409420
rect 456058 409408 456064 409420
rect 453448 409380 456064 409408
rect 453448 409368 453454 409380
rect 456058 409368 456064 409380
rect 456116 409368 456122 409420
rect 3418 402908 3424 402960
rect 3476 402948 3482 402960
rect 128354 402948 128360 402960
rect 3476 402920 128360 402948
rect 3476 402908 3482 402920
rect 128354 402908 128360 402920
rect 128412 402908 128418 402960
rect 453942 402908 453948 402960
rect 454000 402948 454006 402960
rect 542998 402948 543004 402960
rect 454000 402920 543004 402948
rect 454000 402908 454006 402920
rect 542998 402908 543004 402920
rect 543056 402908 543062 402960
rect 453758 395972 453764 396024
rect 453816 396012 453822 396024
rect 580258 396012 580264 396024
rect 453816 395984 580264 396012
rect 453816 395972 453822 395984
rect 580258 395972 580264 395984
rect 580316 395972 580322 396024
rect 3418 394612 3424 394664
rect 3476 394652 3482 394664
rect 128354 394652 128360 394664
rect 3476 394624 128360 394652
rect 3476 394612 3482 394624
rect 128354 394612 128360 394624
rect 128412 394612 128418 394664
rect 460198 391960 460204 392012
rect 460256 392000 460262 392012
rect 580166 392000 580172 392012
rect 460256 391972 580172 392000
rect 460256 391960 460262 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 128998 380848 129004 380860
rect 3292 380820 129004 380848
rect 3292 380808 3298 380820
rect 128998 380808 129004 380820
rect 129056 380808 129062 380860
rect 453942 380808 453948 380860
rect 454000 380848 454006 380860
rect 578878 380848 578884 380860
rect 454000 380820 578884 380848
rect 454000 380808 454006 380820
rect 578878 380808 578884 380820
rect 578936 380808 578942 380860
rect 453390 373940 453396 373992
rect 453448 373980 453454 373992
rect 580350 373980 580356 373992
rect 453448 373952 580356 373980
rect 453448 373940 453454 373952
rect 580350 373940 580356 373952
rect 580408 373940 580414 373992
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 128998 367044 129004 367056
rect 3200 367016 129004 367044
rect 3200 367004 3206 367016
rect 128998 367004 129004 367016
rect 129056 367004 129062 367056
rect 453942 366664 453948 366716
rect 454000 366704 454006 366716
rect 460198 366704 460204 366716
rect 454000 366676 460204 366704
rect 454000 366664 454006 366676
rect 460198 366664 460204 366676
rect 460256 366664 460262 366716
rect 453942 360136 453948 360188
rect 454000 360176 454006 360188
rect 580258 360176 580264 360188
rect 454000 360148 580264 360176
rect 454000 360136 454006 360148
rect 580258 360136 580264 360148
rect 580316 360136 580322 360188
rect 453758 353200 453764 353252
rect 453816 353240 453822 353252
rect 580258 353240 580264 353252
rect 453816 353212 580264 353240
rect 453816 353200 453822 353212
rect 580258 353200 580264 353212
rect 580316 353200 580322 353252
rect 3418 347760 3424 347812
rect 3476 347800 3482 347812
rect 128354 347800 128360 347812
rect 3476 347772 128360 347800
rect 3476 347760 3482 347772
rect 128354 347760 128360 347772
rect 128412 347760 128418 347812
rect 453942 345652 453948 345704
rect 454000 345692 454006 345704
rect 580166 345692 580172 345704
rect 454000 345664 580172 345692
rect 454000 345652 454006 345664
rect 580166 345652 580172 345664
rect 580224 345652 580230 345704
rect 3510 338036 3516 338088
rect 3568 338076 3574 338088
rect 129274 338076 129280 338088
rect 3568 338048 129280 338076
rect 3568 338036 3574 338048
rect 129274 338036 129280 338048
rect 129332 338036 129338 338088
rect 8938 332596 8944 332648
rect 8996 332636 9002 332648
rect 128354 332636 128360 332648
rect 8996 332608 128360 332636
rect 8996 332596 9002 332608
rect 128354 332596 128360 332608
rect 128412 332596 128418 332648
rect 7558 324300 7564 324352
rect 7616 324340 7622 324352
rect 128354 324340 128360 324352
rect 7616 324312 128360 324340
rect 7616 324300 7622 324312
rect 128354 324300 128360 324312
rect 128412 324300 128418 324352
rect 3510 324232 3516 324284
rect 3568 324272 3574 324284
rect 128998 324272 129004 324284
rect 3568 324244 129004 324272
rect 3568 324232 3574 324244
rect 128998 324232 129004 324244
rect 129056 324232 129062 324284
rect 453482 322872 453488 322924
rect 453540 322912 453546 322924
rect 580166 322912 580172 322924
rect 453540 322884 580172 322912
rect 453540 322872 453546 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 453390 311788 453396 311840
rect 453448 311828 453454 311840
rect 580166 311828 580172 311840
rect 453448 311800 580172 311828
rect 453448 311788 453454 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 11698 309136 11704 309188
rect 11756 309176 11762 309188
rect 128354 309176 128360 309188
rect 11756 309148 128360 309176
rect 11756 309136 11762 309148
rect 128354 309136 128360 309148
rect 128412 309136 128418 309188
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 129182 309108 129188 309120
rect 3384 309080 129188 309108
rect 3384 309068 3390 309080
rect 129182 309068 129188 309080
rect 129240 309068 129246 309120
rect 453666 302336 453672 302388
rect 453724 302376 453730 302388
rect 456058 302376 456064 302388
rect 453724 302348 456064 302376
rect 453724 302336 453730 302348
rect 456058 302336 456064 302348
rect 456116 302336 456122 302388
rect 6178 302200 6184 302252
rect 6236 302240 6242 302252
rect 128354 302240 128360 302252
rect 6236 302212 128360 302240
rect 6236 302200 6242 302212
rect 128354 302200 128360 302212
rect 128412 302200 128418 302252
rect 453298 299412 453304 299464
rect 453356 299452 453362 299464
rect 579798 299452 579804 299464
rect 453356 299424 579804 299452
rect 453356 299412 453362 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 13078 287036 13084 287088
rect 13136 287076 13142 287088
rect 128354 287076 128360 287088
rect 13136 287048 128360 287076
rect 13136 287036 13142 287048
rect 128354 287036 128360 287048
rect 128412 287036 128418 287088
rect 453942 280168 453948 280220
rect 454000 280208 454006 280220
rect 461578 280208 461584 280220
rect 454000 280180 461584 280208
rect 454000 280168 454006 280180
rect 461578 280168 461584 280180
rect 461636 280168 461642 280220
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 129090 280140 129096 280152
rect 3476 280112 129096 280140
rect 3476 280100 3482 280112
rect 129090 280100 129096 280112
rect 129148 280100 129154 280152
rect 3418 277992 3424 278044
rect 3476 278032 3482 278044
rect 128262 278032 128268 278044
rect 3476 278004 128268 278032
rect 3476 277992 3482 278004
rect 128262 277992 128268 278004
rect 128320 277992 128326 278044
rect 453574 275952 453580 276004
rect 453632 275992 453638 276004
rect 580166 275992 580172 276004
rect 453632 275964 580172 275992
rect 453632 275952 453638 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3510 266024 3516 266076
rect 3568 266064 3574 266076
rect 8938 266064 8944 266076
rect 3568 266036 8944 266064
rect 3568 266024 3574 266036
rect 8938 266024 8944 266036
rect 8996 266024 9002 266076
rect 453482 264868 453488 264920
rect 453540 264908 453546 264920
rect 580166 264908 580172 264920
rect 453540 264880 580172 264908
rect 453540 264868 453546 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 8938 263576 8944 263628
rect 8996 263616 9002 263628
rect 128354 263616 128360 263628
rect 8996 263588 128360 263616
rect 8996 263576 9002 263588
rect 128354 263576 128360 263588
rect 128412 263576 128418 263628
rect 453942 259428 453948 259480
rect 454000 259468 454006 259480
rect 471238 259468 471244 259480
rect 454000 259440 471244 259468
rect 454000 259428 454006 259440
rect 471238 259428 471244 259440
rect 471296 259428 471302 259480
rect 10318 256708 10324 256760
rect 10376 256748 10382 256760
rect 128354 256748 128360 256760
rect 10376 256720 128360 256748
rect 10376 256708 10382 256720
rect 128354 256708 128360 256720
rect 128412 256708 128418 256760
rect 456058 252492 456064 252544
rect 456116 252532 456122 252544
rect 579798 252532 579804 252544
rect 456116 252504 579804 252532
rect 456116 252492 456122 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3510 251608 3516 251660
rect 3568 251648 3574 251660
rect 7558 251648 7564 251660
rect 3568 251620 7564 251648
rect 3568 251608 3574 251620
rect 7558 251608 7564 251620
rect 7616 251608 7622 251660
rect 453022 251200 453028 251252
rect 453080 251240 453086 251252
rect 457438 251240 457444 251252
rect 453080 251212 457444 251240
rect 453080 251200 453086 251212
rect 457438 251200 457444 251212
rect 457496 251200 457502 251252
rect 15838 241476 15844 241528
rect 15896 241516 15902 241528
rect 128354 241516 128360 241528
rect 15896 241488 128360 241516
rect 15896 241476 15902 241488
rect 128354 241476 128360 241488
rect 128412 241476 128418 241528
rect 453942 237396 453948 237448
rect 454000 237436 454006 237448
rect 469858 237436 469864 237448
rect 454000 237408 469864 237436
rect 454000 237396 454006 237408
rect 469858 237396 469864 237408
rect 469916 237396 469922 237448
rect 3510 237328 3516 237380
rect 3568 237368 3574 237380
rect 128998 237368 129004 237380
rect 3568 237340 129004 237368
rect 3568 237328 3574 237340
rect 128998 237328 129004 237340
rect 129056 237328 129062 237380
rect 14458 233248 14464 233300
rect 14516 233288 14522 233300
rect 128354 233288 128360 233300
rect 14516 233260 128360 233288
rect 14516 233248 14522 233260
rect 128354 233248 128360 233260
rect 128412 233248 128418 233300
rect 453114 230460 453120 230512
rect 453172 230500 453178 230512
rect 473998 230500 474004 230512
rect 453172 230472 474004 230500
rect 453172 230460 453178 230472
rect 473998 230460 474004 230472
rect 474056 230460 474062 230512
rect 453390 229032 453396 229084
rect 453448 229072 453454 229084
rect 580166 229072 580172 229084
rect 453448 229044 580172 229072
rect 453448 229032 453454 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 11698 223564 11704 223576
rect 3200 223536 11704 223564
rect 3200 223524 3206 223536
rect 11698 223524 11704 223536
rect 11756 223524 11762 223576
rect 11698 218016 11704 218068
rect 11756 218056 11762 218068
rect 128354 218056 128360 218068
rect 11756 218028 128360 218056
rect 11756 218016 11762 218028
rect 128354 218016 128360 218028
rect 128412 218016 128418 218068
rect 453298 217948 453304 218000
rect 453356 217988 453362 218000
rect 580166 217988 580172 218000
rect 453356 217960 580172 217988
rect 453356 217948 453362 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 453758 216792 453764 216844
rect 453816 216832 453822 216844
rect 456058 216832 456064 216844
rect 453816 216804 456064 216832
rect 453816 216792 453822 216804
rect 456058 216792 456064 216804
rect 456116 216792 456122 216844
rect 7558 211148 7564 211200
rect 7616 211188 7622 211200
rect 128354 211188 128360 211200
rect 7616 211160 128360 211188
rect 7616 211148 7622 211160
rect 128354 211148 128360 211160
rect 128412 211148 128418 211200
rect 453942 209788 453948 209840
rect 454000 209828 454006 209840
rect 478138 209828 478144 209840
rect 454000 209800 478144 209828
rect 454000 209788 454006 209800
rect 478138 209788 478144 209800
rect 478196 209788 478202 209840
rect 3142 208156 3148 208208
rect 3200 208196 3206 208208
rect 6178 208196 6184 208208
rect 3200 208168 6184 208196
rect 3200 208156 3206 208168
rect 6178 208156 6184 208168
rect 6236 208156 6242 208208
rect 461578 205572 461584 205624
rect 461636 205612 461642 205624
rect 579798 205612 579804 205624
rect 461636 205584 579804 205612
rect 461636 205572 461642 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 6178 194556 6184 194608
rect 6236 194596 6242 194608
rect 128630 194596 128636 194608
rect 6236 194568 128636 194596
rect 6236 194556 6242 194568
rect 128630 194556 128636 194568
rect 128688 194556 128694 194608
rect 453942 194556 453948 194608
rect 454000 194596 454006 194608
rect 483658 194596 483664 194608
rect 454000 194568 483664 194596
rect 454000 194556 454006 194568
rect 483658 194556 483664 194568
rect 483716 194556 483722 194608
rect 2866 194488 2872 194540
rect 2924 194528 2930 194540
rect 129366 194528 129372 194540
rect 2924 194500 129372 194528
rect 2924 194488 2930 194500
rect 129366 194488 129372 194500
rect 129424 194488 129430 194540
rect 303890 190340 303896 190392
rect 303948 190380 303954 190392
rect 304810 190380 304816 190392
rect 303948 190352 304816 190380
rect 303948 190340 303954 190352
rect 304810 190340 304816 190352
rect 304868 190340 304874 190392
rect 168650 190272 168656 190324
rect 168708 190312 168714 190324
rect 169570 190312 169576 190324
rect 168708 190284 169576 190312
rect 168708 190272 168714 190284
rect 169570 190272 169576 190284
rect 169628 190272 169634 190324
rect 201586 190204 201592 190256
rect 201644 190244 201650 190256
rect 204898 190244 204904 190256
rect 201644 190216 204904 190244
rect 201644 190204 201650 190216
rect 204898 190204 204904 190216
rect 204956 190204 204962 190256
rect 332778 190204 332784 190256
rect 332836 190244 332842 190256
rect 333882 190244 333888 190256
rect 332836 190216 333888 190244
rect 332836 190204 332842 190216
rect 333882 190204 333888 190216
rect 333940 190204 333946 190256
rect 375650 190204 375656 190256
rect 375708 190244 375714 190256
rect 376662 190244 376668 190256
rect 375708 190216 376668 190244
rect 375708 190204 375714 190216
rect 376662 190204 376668 190216
rect 376720 190204 376726 190256
rect 392118 190204 392124 190256
rect 392176 190244 392182 190256
rect 393130 190244 393136 190256
rect 392176 190216 393136 190244
rect 392176 190204 392182 190216
rect 393130 190204 393136 190216
rect 393188 190204 393194 190256
rect 416866 190204 416872 190256
rect 416924 190244 416930 190256
rect 417970 190244 417976 190256
rect 416924 190216 417976 190244
rect 416924 190204 416930 190216
rect 417970 190204 417976 190216
rect 418028 190204 418034 190256
rect 434990 190204 434996 190256
rect 435048 190244 435054 190256
rect 435910 190244 435916 190256
rect 435048 190216 435916 190244
rect 435048 190204 435054 190216
rect 435910 190204 435916 190216
rect 435968 190204 435974 190256
rect 281626 190136 281632 190188
rect 281684 190176 281690 190188
rect 282730 190176 282736 190188
rect 281684 190148 282736 190176
rect 281684 190136 281690 190148
rect 282730 190136 282736 190148
rect 282788 190136 282794 190188
rect 408586 190136 408592 190188
rect 408644 190176 408650 190188
rect 409690 190176 409696 190188
rect 408644 190148 409696 190176
rect 408644 190136 408650 190148
rect 409690 190136 409696 190148
rect 409748 190136 409754 190188
rect 441614 190136 441620 190188
rect 441672 190176 441678 190188
rect 442810 190176 442816 190188
rect 441672 190148 442816 190176
rect 441672 190136 441678 190148
rect 442810 190136 442816 190148
rect 442868 190136 442874 190188
rect 154666 190068 154672 190120
rect 154724 190108 154730 190120
rect 155770 190108 155776 190120
rect 154724 190080 155776 190108
rect 154724 190068 154730 190080
rect 155770 190068 155776 190080
rect 155828 190068 155834 190120
rect 164510 190068 164516 190120
rect 164568 190108 164574 190120
rect 165430 190108 165436 190120
rect 164568 190080 165436 190108
rect 164568 190068 164574 190080
rect 165430 190068 165436 190080
rect 165488 190068 165494 190120
rect 244550 190068 244556 190120
rect 244608 190108 244614 190120
rect 245470 190108 245476 190120
rect 244608 190080 245476 190108
rect 244608 190068 244614 190080
rect 245470 190068 245476 190080
rect 245528 190068 245534 190120
rect 253566 190068 253572 190120
rect 253624 190108 253630 190120
rect 257338 190108 257344 190120
rect 253624 190080 257344 190108
rect 253624 190068 253630 190080
rect 257338 190068 257344 190080
rect 257396 190068 257402 190120
rect 316218 190068 316224 190120
rect 316276 190108 316282 190120
rect 317230 190108 317236 190120
rect 316276 190080 317236 190108
rect 316276 190068 316282 190080
rect 317230 190068 317236 190080
rect 317288 190068 317294 190120
rect 345106 190068 345112 190120
rect 345164 190108 345170 190120
rect 346210 190108 346216 190120
rect 345164 190080 346216 190108
rect 345164 190068 345170 190080
rect 346210 190068 346216 190080
rect 346268 190068 346274 190120
rect 353386 190068 353392 190120
rect 353444 190108 353450 190120
rect 354490 190108 354496 190120
rect 353444 190080 354496 190108
rect 353444 190068 353450 190080
rect 354490 190068 354496 190080
rect 354548 190068 354554 190120
rect 433334 190068 433340 190120
rect 433392 190108 433398 190120
rect 434530 190108 434536 190120
rect 433392 190080 434536 190108
rect 433392 190068 433398 190080
rect 434530 190068 434536 190080
rect 434588 190068 434594 190120
rect 226334 190000 226340 190052
rect 226392 190040 226398 190052
rect 227530 190040 227536 190052
rect 226392 190012 227536 190040
rect 226392 190000 226398 190012
rect 227530 190000 227536 190012
rect 227588 190000 227594 190052
rect 369854 190000 369860 190052
rect 369912 190040 369918 190052
rect 371050 190040 371056 190052
rect 369912 190012 371056 190040
rect 369912 190000 369918 190012
rect 371050 190000 371056 190012
rect 371108 190000 371114 190052
rect 162854 189932 162860 189984
rect 162912 189972 162918 189984
rect 164050 189972 164056 189984
rect 162912 189944 164056 189972
rect 162912 189932 162918 189944
rect 164050 189932 164056 189944
rect 164108 189932 164114 189984
rect 237926 189932 237932 189984
rect 237984 189972 237990 189984
rect 238662 189972 238668 189984
rect 237984 189944 238668 189972
rect 237984 189932 237990 189944
rect 238662 189932 238668 189944
rect 238720 189932 238726 189984
rect 269206 189932 269212 189984
rect 269264 189972 269270 189984
rect 270310 189972 270316 189984
rect 269264 189944 270316 189972
rect 269264 189932 269270 189944
rect 270310 189932 270316 189944
rect 270368 189932 270374 189984
rect 329466 189932 329472 189984
rect 329524 189972 329530 189984
rect 331858 189972 331864 189984
rect 329524 189944 331864 189972
rect 329524 189932 329530 189944
rect 331858 189932 331864 189944
rect 331916 189932 331922 189984
rect 340966 189932 340972 189984
rect 341024 189972 341030 189984
rect 342070 189972 342076 189984
rect 341024 189944 342076 189972
rect 341024 189932 341030 189944
rect 342070 189932 342076 189944
rect 342128 189932 342134 189984
rect 357526 189932 357532 189984
rect 357584 189972 357590 189984
rect 358630 189972 358636 189984
rect 357584 189944 358636 189972
rect 357584 189932 357590 189944
rect 358630 189932 358636 189944
rect 358688 189932 358694 189984
rect 373166 189932 373172 189984
rect 373224 189972 373230 189984
rect 373902 189972 373908 189984
rect 373224 189944 373908 189972
rect 373224 189932 373230 189944
rect 373902 189932 373908 189944
rect 373960 189932 373966 189984
rect 429194 189932 429200 189984
rect 429252 189972 429258 189984
rect 430390 189972 430396 189984
rect 429252 189944 430396 189972
rect 429252 189932 429258 189944
rect 430390 189932 430396 189944
rect 430448 189932 430454 189984
rect 445754 189932 445760 189984
rect 445812 189972 445818 189984
rect 446950 189972 446956 189984
rect 445812 189944 446956 189972
rect 445812 189932 445818 189944
rect 446950 189932 446956 189944
rect 447008 189932 447014 189984
rect 310514 189864 310520 189916
rect 310572 189904 310578 189916
rect 315298 189904 315304 189916
rect 310572 189876 315304 189904
rect 310572 189864 310578 189876
rect 315298 189864 315304 189876
rect 315356 189864 315362 189916
rect 382274 189864 382280 189916
rect 382332 189904 382338 189916
rect 387058 189904 387064 189916
rect 382332 189876 387064 189904
rect 382332 189864 382338 189876
rect 387058 189864 387064 189876
rect 387116 189864 387122 189916
rect 158714 189796 158720 189848
rect 158772 189836 158778 189848
rect 159910 189836 159916 189848
rect 158772 189808 159916 189836
rect 158772 189796 158778 189808
rect 159910 189796 159916 189808
rect 159968 189796 159974 189848
rect 178494 189796 178500 189848
rect 178552 189836 178558 189848
rect 188338 189836 188344 189848
rect 178552 189808 188344 189836
rect 178552 189796 178558 189808
rect 188338 189796 188344 189808
rect 188396 189796 188402 189848
rect 240410 189796 240416 189848
rect 240468 189836 240474 189848
rect 255958 189836 255964 189848
rect 240468 189808 255964 189836
rect 240468 189796 240474 189808
rect 255958 189796 255964 189808
rect 256016 189796 256022 189848
rect 257706 189796 257712 189848
rect 257764 189836 257770 189848
rect 301498 189836 301504 189848
rect 257764 189808 301504 189836
rect 257764 189796 257770 189808
rect 301498 189796 301504 189808
rect 301556 189796 301562 189848
rect 349246 189796 349252 189848
rect 349304 189836 349310 189848
rect 384298 189836 384304 189848
rect 349304 189808 384304 189836
rect 349304 189796 349310 189808
rect 384298 189796 384304 189808
rect 384356 189796 384362 189848
rect 411070 189796 411076 189848
rect 411128 189836 411134 189848
rect 451918 189836 451924 189848
rect 411128 189808 451924 189836
rect 411128 189796 411134 189808
rect 451918 189796 451924 189808
rect 451976 189796 451982 189848
rect 180978 189728 180984 189780
rect 181036 189768 181042 189780
rect 192478 189768 192484 189780
rect 181036 189740 192484 189768
rect 181036 189728 181042 189740
rect 192478 189728 192484 189740
rect 192536 189728 192542 189780
rect 195882 189728 195888 189780
rect 195940 189768 195946 189780
rect 213178 189768 213184 189780
rect 195940 189740 213184 189768
rect 195940 189728 195946 189740
rect 213178 189728 213184 189740
rect 213236 189728 213242 189780
rect 223114 189728 223120 189780
rect 223172 189768 223178 189780
rect 242158 189768 242164 189780
rect 223172 189740 242164 189768
rect 223172 189728 223178 189740
rect 242158 189728 242164 189740
rect 242216 189728 242222 189780
rect 275002 189728 275008 189780
rect 275060 189768 275066 189780
rect 280798 189768 280804 189780
rect 275060 189740 280804 189768
rect 275060 189728 275066 189740
rect 280798 189728 280804 189740
rect 280856 189728 280862 189780
rect 294782 189728 294788 189780
rect 294840 189768 294846 189780
rect 352558 189768 352564 189780
rect 294840 189740 352564 189768
rect 294840 189728 294846 189740
rect 352558 189728 352564 189740
rect 352616 189728 352622 189780
rect 383838 189728 383844 189780
rect 383896 189768 383902 189780
rect 485774 189768 485780 189780
rect 383896 189740 485780 189768
rect 383896 189728 383902 189740
rect 485774 189728 485780 189740
rect 485832 189728 485838 189780
rect 229646 189660 229652 189712
rect 229704 189700 229710 189712
rect 230382 189700 230388 189712
rect 229704 189672 230388 189700
rect 229704 189660 229710 189672
rect 230382 189660 230388 189672
rect 230440 189660 230446 189712
rect 309686 189660 309692 189712
rect 309744 189700 309750 189712
rect 310422 189700 310428 189712
rect 309744 189672 310428 189700
rect 309744 189660 309750 189672
rect 310422 189660 310428 189672
rect 310480 189660 310486 189712
rect 222286 189456 222292 189508
rect 222344 189496 222350 189508
rect 223482 189496 223488 189508
rect 222344 189468 223488 189496
rect 222344 189456 222350 189468
rect 223482 189456 223488 189468
rect 223540 189456 223546 189508
rect 250254 189456 250260 189508
rect 250312 189496 250318 189508
rect 251082 189496 251088 189508
rect 250312 189468 251088 189496
rect 250312 189456 250318 189468
rect 251082 189456 251088 189468
rect 251140 189456 251146 189508
rect 285766 189456 285772 189508
rect 285824 189496 285830 189508
rect 286962 189496 286968 189508
rect 285824 189468 286968 189496
rect 285824 189456 285830 189468
rect 286962 189456 286968 189468
rect 287020 189456 287026 189508
rect 322014 189456 322020 189508
rect 322072 189496 322078 189508
rect 322842 189496 322848 189508
rect 322072 189468 322848 189496
rect 322072 189456 322078 189468
rect 322842 189456 322848 189468
rect 322900 189456 322906 189508
rect 330294 189456 330300 189508
rect 330352 189496 330358 189508
rect 331122 189496 331128 189508
rect 330352 189468 331128 189496
rect 330352 189456 330358 189468
rect 331122 189456 331128 189468
rect 331180 189456 331186 189508
rect 182634 189388 182640 189440
rect 182692 189428 182698 189440
rect 183462 189428 183468 189440
rect 182692 189400 183468 189428
rect 182692 189388 182698 189400
rect 183462 189388 183468 189400
rect 183520 189388 183526 189440
rect 203242 189388 203248 189440
rect 203300 189428 203306 189440
rect 204162 189428 204168 189440
rect 203300 189400 204168 189428
rect 203300 189388 203306 189400
rect 204162 189388 204168 189400
rect 204220 189388 204226 189440
rect 219802 189388 219808 189440
rect 219860 189428 219866 189440
rect 220630 189428 220636 189440
rect 219860 189400 220636 189428
rect 219860 189388 219866 189400
rect 220630 189388 220636 189400
rect 220688 189388 220694 189440
rect 283282 189388 283288 189440
rect 283340 189428 283346 189440
rect 284202 189428 284208 189440
rect 283340 189400 284208 189428
rect 283340 189388 283346 189400
rect 284202 189388 284208 189400
rect 284260 189388 284266 189440
rect 293954 189388 293960 189440
rect 294012 189428 294018 189440
rect 295242 189428 295248 189440
rect 294012 189400 295248 189428
rect 294012 189388 294018 189400
rect 295242 189388 295248 189400
rect 295300 189388 295306 189440
rect 328638 189388 328644 189440
rect 328696 189428 328702 189440
rect 329742 189428 329748 189440
rect 328696 189400 329748 189428
rect 328696 189388 328702 189400
rect 329742 189388 329748 189400
rect 329800 189388 329806 189440
rect 389634 189388 389640 189440
rect 389692 189428 389698 189440
rect 390462 189428 390468 189440
rect 389692 189400 390468 189428
rect 389692 189388 389698 189400
rect 390462 189388 390468 189400
rect 390520 189388 390526 189440
rect 156230 189320 156236 189372
rect 156288 189360 156294 189372
rect 157242 189360 157248 189372
rect 156288 189332 157248 189360
rect 156288 189320 156294 189332
rect 157242 189320 157248 189332
rect 157300 189320 157306 189372
rect 172790 189320 172796 189372
rect 172848 189360 172854 189372
rect 173802 189360 173808 189372
rect 172848 189332 173808 189360
rect 172848 189320 172854 189332
rect 173802 189320 173808 189332
rect 173860 189320 173866 189372
rect 197538 189320 197544 189372
rect 197596 189360 197602 189372
rect 198642 189360 198648 189372
rect 197596 189332 198648 189360
rect 197596 189320 197602 189332
rect 198642 189320 198648 189332
rect 198700 189320 198706 189372
rect 214006 189320 214012 189372
rect 214064 189360 214070 189372
rect 215202 189360 215208 189372
rect 214064 189332 215208 189360
rect 214064 189320 214070 189332
rect 215202 189320 215208 189332
rect 215260 189320 215266 189372
rect 236270 189320 236276 189372
rect 236328 189360 236334 189372
rect 237282 189360 237288 189372
rect 236328 189332 237288 189360
rect 236328 189320 236334 189332
rect 237282 189320 237288 189332
rect 237340 189320 237346 189372
rect 261018 189320 261024 189372
rect 261076 189360 261082 189372
rect 262122 189360 262128 189372
rect 261076 189332 262128 189360
rect 261076 189320 261082 189332
rect 262122 189320 262128 189332
rect 262180 189320 262186 189372
rect 277486 189320 277492 189372
rect 277544 189360 277550 189372
rect 278682 189360 278688 189372
rect 277544 189332 278688 189360
rect 277544 189320 277550 189332
rect 278682 189320 278688 189332
rect 278740 189320 278746 189372
rect 299750 189320 299756 189372
rect 299808 189360 299814 189372
rect 300762 189360 300768 189372
rect 299808 189332 300768 189360
rect 299808 189320 299814 189332
rect 300762 189320 300768 189332
rect 300820 189320 300826 189372
rect 371510 189320 371516 189372
rect 371568 189360 371574 189372
rect 372522 189360 372528 189372
rect 371568 189332 372528 189360
rect 371568 189320 371574 189332
rect 372522 189320 372528 189332
rect 372580 189320 372586 189372
rect 412726 189320 412732 189372
rect 412784 189360 412790 189372
rect 413922 189360 413928 189372
rect 412784 189332 413928 189360
rect 412784 189320 412790 189332
rect 413922 189320 413928 189332
rect 413980 189320 413986 189372
rect 175274 189252 175280 189304
rect 175332 189292 175338 189304
rect 176562 189292 176568 189304
rect 175332 189264 176568 189292
rect 175332 189252 175338 189264
rect 176562 189252 176568 189264
rect 176620 189252 176626 189304
rect 185118 189252 185124 189304
rect 185176 189292 185182 189304
rect 186222 189292 186228 189304
rect 185176 189264 186228 189292
rect 185176 189252 185182 189264
rect 186222 189252 186228 189264
rect 186280 189252 186286 189304
rect 193398 189252 193404 189304
rect 193456 189292 193462 189304
rect 194502 189292 194508 189304
rect 193456 189264 194508 189292
rect 193456 189252 193462 189264
rect 194502 189252 194508 189264
rect 194560 189252 194566 189304
rect 205726 189252 205732 189304
rect 205784 189292 205790 189304
rect 206922 189292 206928 189304
rect 205784 189264 206928 189292
rect 205784 189252 205790 189264
rect 206922 189252 206928 189264
rect 206980 189252 206986 189304
rect 209866 189252 209872 189304
rect 209924 189292 209930 189304
rect 211062 189292 211068 189304
rect 209924 189264 211068 189292
rect 209924 189252 209930 189264
rect 211062 189252 211068 189264
rect 211120 189252 211126 189304
rect 221458 189252 221464 189304
rect 221516 189292 221522 189304
rect 222838 189292 222844 189304
rect 221516 189264 222844 189292
rect 221516 189252 221522 189264
rect 222838 189252 222844 189264
rect 222896 189252 222902 189304
rect 223850 189252 223856 189304
rect 223908 189292 223914 189304
rect 224862 189292 224868 189304
rect 223908 189264 224868 189292
rect 223908 189252 223914 189264
rect 224862 189252 224868 189264
rect 224920 189252 224926 189304
rect 230474 189252 230480 189304
rect 230532 189292 230538 189304
rect 231762 189292 231768 189304
rect 230532 189264 231768 189292
rect 230532 189252 230538 189264
rect 231762 189252 231768 189264
rect 231820 189252 231826 189304
rect 234614 189252 234620 189304
rect 234672 189292 234678 189304
rect 235902 189292 235908 189304
rect 234672 189264 235908 189292
rect 234672 189252 234678 189264
rect 235902 189252 235908 189264
rect 235960 189252 235966 189304
rect 238754 189252 238760 189304
rect 238812 189292 238818 189304
rect 240042 189292 240048 189304
rect 238812 189264 240048 189292
rect 238812 189252 238818 189264
rect 240042 189252 240048 189264
rect 240100 189252 240106 189304
rect 248598 189252 248604 189304
rect 248656 189292 248662 189304
rect 249702 189292 249708 189304
rect 248656 189264 249708 189292
rect 248656 189252 248662 189264
rect 249702 189252 249708 189264
rect 249760 189252 249766 189304
rect 265158 189252 265164 189304
rect 265216 189292 265222 189304
rect 266262 189292 266268 189304
rect 265216 189264 266268 189292
rect 265216 189252 265222 189264
rect 266262 189252 266268 189264
rect 266320 189252 266326 189304
rect 270862 189252 270868 189304
rect 270920 189292 270926 189304
rect 271966 189292 271972 189304
rect 270920 189264 271972 189292
rect 270920 189252 270926 189264
rect 271966 189252 271972 189264
rect 272024 189252 272030 189304
rect 302234 189252 302240 189304
rect 302292 189292 302298 189304
rect 303522 189292 303528 189304
rect 302292 189264 303528 189292
rect 302292 189252 302298 189264
rect 303522 189252 303528 189264
rect 303580 189252 303586 189304
rect 306374 189252 306380 189304
rect 306432 189292 306438 189304
rect 307662 189292 307668 189304
rect 306432 189264 307668 189292
rect 306432 189252 306438 189264
rect 307662 189252 307668 189264
rect 307720 189252 307726 189304
rect 312170 189252 312176 189304
rect 312228 189292 312234 189304
rect 313182 189292 313188 189304
rect 312228 189264 313188 189292
rect 312228 189252 312234 189264
rect 313182 189252 313188 189264
rect 313240 189252 313246 189304
rect 320358 189252 320364 189304
rect 320416 189292 320422 189304
rect 321462 189292 321468 189304
rect 320416 189264 321468 189292
rect 320416 189252 320422 189264
rect 321462 189252 321468 189264
rect 321520 189252 321526 189304
rect 336918 189252 336924 189304
rect 336976 189292 336982 189304
rect 338022 189292 338028 189304
rect 336976 189264 338028 189292
rect 336976 189252 336982 189264
rect 338022 189252 338028 189264
rect 338080 189252 338086 189304
rect 365714 189252 365720 189304
rect 365772 189292 365778 189304
rect 367002 189292 367008 189304
rect 365772 189264 367008 189292
rect 365772 189252 365778 189264
rect 367002 189252 367008 189264
rect 367060 189252 367066 189304
rect 373994 189252 374000 189304
rect 374052 189292 374058 189304
rect 375282 189292 375288 189304
rect 374052 189264 375288 189292
rect 374052 189252 374058 189264
rect 375282 189252 375288 189264
rect 375340 189252 375346 189304
rect 378134 189252 378140 189304
rect 378192 189292 378198 189304
rect 379422 189292 379428 189304
rect 378192 189264 379428 189292
rect 378192 189252 378198 189264
rect 379422 189252 379428 189264
rect 379480 189252 379486 189304
rect 425146 189252 425152 189304
rect 425204 189292 425210 189304
rect 426342 189292 426348 189304
rect 425204 189264 426348 189292
rect 425204 189252 425210 189264
rect 426342 189252 426348 189264
rect 426400 189252 426406 189304
rect 437474 189252 437480 189304
rect 437532 189292 437538 189304
rect 438762 189292 438768 189304
rect 437532 189264 438768 189292
rect 437532 189252 437538 189264
rect 438762 189252 438768 189264
rect 438820 189252 438826 189304
rect 439130 189252 439136 189304
rect 439188 189292 439194 189304
rect 440050 189292 440056 189304
rect 439188 189264 440056 189292
rect 439188 189252 439194 189264
rect 440050 189252 440056 189264
rect 440108 189252 440114 189304
rect 160370 189116 160376 189168
rect 160428 189156 160434 189168
rect 161382 189156 161388 189168
rect 160428 189128 161388 189156
rect 160428 189116 160434 189128
rect 161382 189116 161388 189128
rect 161440 189116 161446 189168
rect 213546 189116 213552 189168
rect 213604 189156 213610 189168
rect 221458 189156 221464 189168
rect 213604 189128 221464 189156
rect 213604 189116 213610 189128
rect 221458 189116 221464 189128
rect 221516 189116 221522 189168
rect 307202 189116 307208 189168
rect 307260 189156 307266 189168
rect 309778 189156 309784 189168
rect 307260 189128 309784 189156
rect 307260 189116 307266 189128
rect 309778 189116 309784 189128
rect 309836 189116 309842 189168
rect 378962 189116 378968 189168
rect 379020 189156 379026 189168
rect 381538 189156 381544 189168
rect 379020 189128 381544 189156
rect 379020 189116 379026 189128
rect 381538 189116 381544 189128
rect 381596 189116 381602 189168
rect 157886 189048 157892 189100
rect 157944 189088 157950 189100
rect 158622 189088 158628 189100
rect 157944 189060 158628 189088
rect 157944 189048 157950 189060
rect 158622 189048 158628 189060
rect 158680 189048 158686 189100
rect 166166 189048 166172 189100
rect 166224 189088 166230 189100
rect 166902 189088 166908 189100
rect 166224 189060 166908 189088
rect 166224 189048 166230 189060
rect 166902 189048 166908 189060
rect 166960 189048 166966 189100
rect 166994 189048 167000 189100
rect 167052 189088 167058 189100
rect 168190 189088 168196 189100
rect 167052 189060 168196 189088
rect 167052 189048 167058 189060
rect 168190 189048 168196 189060
rect 168248 189048 168254 189100
rect 171134 189048 171140 189100
rect 171192 189088 171198 189100
rect 172422 189088 172428 189100
rect 171192 189060 172428 189088
rect 171192 189048 171198 189060
rect 172422 189048 172428 189060
rect 172480 189048 172486 189100
rect 174446 189048 174452 189100
rect 174504 189088 174510 189100
rect 175182 189088 175188 189100
rect 174504 189060 175188 189088
rect 174504 189048 174510 189060
rect 175182 189048 175188 189060
rect 175240 189048 175246 189100
rect 176930 189048 176936 189100
rect 176988 189088 176994 189100
rect 177850 189088 177856 189100
rect 176988 189060 177856 189088
rect 176988 189048 176994 189060
rect 177850 189048 177856 189060
rect 177908 189048 177914 189100
rect 186774 189048 186780 189100
rect 186832 189088 186838 189100
rect 187510 189088 187516 189100
rect 186832 189060 187516 189088
rect 186832 189048 186838 189060
rect 187510 189048 187516 189060
rect 187568 189048 187574 189100
rect 189258 189048 189264 189100
rect 189316 189088 189322 189100
rect 190270 189088 190276 189100
rect 189316 189060 190276 189088
rect 189316 189048 189322 189060
rect 190270 189048 190276 189060
rect 190328 189048 190334 189100
rect 190914 189048 190920 189100
rect 190972 189088 190978 189100
rect 191742 189088 191748 189100
rect 190972 189060 191748 189088
rect 190972 189048 190978 189060
rect 191742 189048 191748 189060
rect 191800 189048 191806 189100
rect 195054 189048 195060 189100
rect 195112 189088 195118 189100
rect 195882 189088 195888 189100
rect 195112 189060 195888 189088
rect 195112 189048 195118 189060
rect 195882 189048 195888 189060
rect 195940 189048 195946 189100
rect 199194 189048 199200 189100
rect 199252 189088 199258 189100
rect 200758 189088 200764 189100
rect 199252 189060 200764 189088
rect 199252 189048 199258 189060
rect 200758 189048 200764 189060
rect 200816 189048 200822 189100
rect 207382 189048 207388 189100
rect 207440 189088 207446 189100
rect 208302 189088 208308 189100
rect 207440 189060 208308 189088
rect 207440 189048 207446 189060
rect 208302 189048 208308 189060
rect 208360 189048 208366 189100
rect 211522 189048 211528 189100
rect 211580 189088 211586 189100
rect 212350 189088 212356 189100
rect 211580 189060 212356 189088
rect 211580 189048 211586 189060
rect 212350 189048 212356 189060
rect 212408 189048 212414 189100
rect 215662 189048 215668 189100
rect 215720 189088 215726 189100
rect 216582 189088 216588 189100
rect 215720 189060 216588 189088
rect 215720 189048 215726 189060
rect 216582 189048 216588 189060
rect 216640 189048 216646 189100
rect 218146 189048 218152 189100
rect 218204 189088 218210 189100
rect 219342 189088 219348 189100
rect 218204 189060 219348 189088
rect 218204 189048 218210 189060
rect 219342 189048 219348 189060
rect 219400 189048 219406 189100
rect 227990 189048 227996 189100
rect 228048 189088 228054 189100
rect 229002 189088 229008 189100
rect 228048 189060 229008 189088
rect 228048 189048 228054 189060
rect 229002 189048 229008 189060
rect 229060 189048 229066 189100
rect 232130 189048 232136 189100
rect 232188 189088 232194 189100
rect 233050 189088 233056 189100
rect 232188 189060 233056 189088
rect 232188 189048 232194 189060
rect 233050 189048 233056 189060
rect 233108 189048 233114 189100
rect 242894 189048 242900 189100
rect 242952 189088 242958 189100
rect 244182 189088 244188 189100
rect 242952 189060 244188 189088
rect 242952 189048 242958 189060
rect 244182 189048 244188 189060
rect 244240 189048 244246 189100
rect 246114 189048 246120 189100
rect 246172 189088 246178 189100
rect 246942 189088 246948 189100
rect 246172 189060 246948 189088
rect 246172 189048 246178 189060
rect 246942 189048 246948 189060
rect 247000 189048 247006 189100
rect 256878 189048 256884 189100
rect 256936 189088 256942 189100
rect 257982 189088 257988 189100
rect 256936 189060 257988 189088
rect 256936 189048 256942 189060
rect 257982 189048 257988 189060
rect 258040 189048 258046 189100
rect 258534 189048 258540 189100
rect 258592 189088 258598 189100
rect 259270 189088 259276 189100
rect 258592 189060 259276 189088
rect 258592 189048 258598 189060
rect 259270 189048 259276 189060
rect 259328 189048 259334 189100
rect 262674 189048 262680 189100
rect 262732 189088 262738 189100
rect 263502 189088 263508 189100
rect 262732 189060 263508 189088
rect 262732 189048 262738 189060
rect 263502 189048 263508 189060
rect 263560 189048 263566 189100
rect 266814 189048 266820 189100
rect 266872 189088 266878 189100
rect 267550 189088 267556 189100
rect 266872 189060 267556 189088
rect 266872 189048 266878 189060
rect 267550 189048 267556 189060
rect 267608 189048 267614 189100
rect 273346 189048 273352 189100
rect 273404 189088 273410 189100
rect 274542 189088 274548 189100
rect 273404 189060 274548 189088
rect 273404 189048 273410 189060
rect 274542 189048 274548 189060
rect 274600 189048 274606 189100
rect 279142 189048 279148 189100
rect 279200 189088 279206 189100
rect 279970 189088 279976 189100
rect 279200 189060 279976 189088
rect 279200 189048 279206 189060
rect 279970 189048 279976 189060
rect 280028 189048 280034 189100
rect 287422 189048 287428 189100
rect 287480 189088 287486 189100
rect 288342 189088 288348 189100
rect 287480 189060 288348 189088
rect 287480 189048 287486 189060
rect 288342 189048 288348 189060
rect 288400 189048 288406 189100
rect 289906 189048 289912 189100
rect 289964 189088 289970 189100
rect 291102 189088 291108 189100
rect 289964 189060 291108 189088
rect 289964 189048 289970 189060
rect 291102 189048 291108 189060
rect 291160 189048 291166 189100
rect 291562 189048 291568 189100
rect 291620 189088 291626 189100
rect 292390 189088 292396 189100
rect 291620 189060 292396 189088
rect 291620 189048 291626 189060
rect 292390 189048 292396 189060
rect 292448 189048 292454 189100
rect 293126 189048 293132 189100
rect 293184 189088 293190 189100
rect 293862 189088 293868 189100
rect 293184 189060 293868 189088
rect 293184 189048 293190 189060
rect 293862 189048 293868 189060
rect 293920 189048 293926 189100
rect 295610 189048 295616 189100
rect 295668 189088 295674 189100
rect 296622 189088 296628 189100
rect 295668 189060 296628 189088
rect 295668 189048 295674 189060
rect 296622 189048 296628 189060
rect 296680 189048 296686 189100
rect 298094 189048 298100 189100
rect 298152 189088 298158 189100
rect 299382 189088 299388 189100
rect 298152 189060 299388 189088
rect 298152 189048 298158 189060
rect 299382 189048 299388 189060
rect 299440 189048 299446 189100
rect 301406 189048 301412 189100
rect 301464 189088 301470 189100
rect 302142 189088 302148 189100
rect 301464 189060 302148 189088
rect 301464 189048 301470 189060
rect 302142 189048 302148 189060
rect 302200 189048 302206 189100
rect 308030 189048 308036 189100
rect 308088 189088 308094 189100
rect 308950 189088 308956 189100
rect 308088 189060 308956 189088
rect 308088 189048 308094 189060
rect 308950 189048 308956 189060
rect 309008 189048 309014 189100
rect 324498 189048 324504 189100
rect 324556 189088 324562 189100
rect 327718 189088 327724 189100
rect 324556 189060 327724 189088
rect 324556 189048 324562 189060
rect 327718 189048 327724 189060
rect 327776 189048 327782 189100
rect 338482 189048 338488 189100
rect 338540 189088 338546 189100
rect 339310 189088 339316 189100
rect 338540 189060 339316 189088
rect 338540 189048 338546 189060
rect 339310 189048 339316 189060
rect 339368 189048 339374 189100
rect 342622 189048 342628 189100
rect 342680 189088 342686 189100
rect 344278 189088 344284 189100
rect 342680 189060 344284 189088
rect 342680 189048 342686 189060
rect 344278 189048 344284 189060
rect 344336 189048 344342 189100
rect 346762 189048 346768 189100
rect 346820 189088 346826 189100
rect 348418 189088 348424 189100
rect 346820 189060 348424 189088
rect 346820 189048 346826 189060
rect 348418 189048 348424 189060
rect 348476 189048 348482 189100
rect 350902 189048 350908 189100
rect 350960 189088 350966 189100
rect 351730 189088 351736 189100
rect 350960 189060 351736 189088
rect 350960 189048 350966 189060
rect 351730 189048 351736 189060
rect 351788 189048 351794 189100
rect 355042 189048 355048 189100
rect 355100 189088 355106 189100
rect 355870 189088 355876 189100
rect 355100 189060 355876 189088
rect 355100 189048 355106 189060
rect 355870 189048 355876 189060
rect 355928 189048 355934 189100
rect 359182 189048 359188 189100
rect 359240 189088 359246 189100
rect 360102 189088 360108 189100
rect 359240 189060 360108 189088
rect 359240 189048 359246 189060
rect 360102 189048 360108 189060
rect 360160 189048 360166 189100
rect 361574 189048 361580 189100
rect 361632 189088 361638 189100
rect 362862 189088 362868 189100
rect 361632 189060 362868 189088
rect 361632 189048 361638 189060
rect 362862 189048 362868 189060
rect 362920 189048 362926 189100
rect 363230 189048 363236 189100
rect 363288 189088 363294 189100
rect 364242 189088 364248 189100
rect 363288 189060 364248 189088
rect 363288 189048 363294 189060
rect 364242 189048 364248 189060
rect 364300 189048 364306 189100
rect 364886 189048 364892 189100
rect 364944 189088 364950 189100
rect 365622 189088 365628 189100
rect 364944 189060 365628 189088
rect 364944 189048 364950 189060
rect 365622 189048 365628 189060
rect 365680 189048 365686 189100
rect 379790 189048 379796 189100
rect 379848 189088 379854 189100
rect 380710 189088 380716 189100
rect 379848 189060 380716 189088
rect 379848 189048 379854 189060
rect 380710 189048 380716 189060
rect 380768 189048 380774 189100
rect 381446 189048 381452 189100
rect 381504 189088 381510 189100
rect 382182 189088 382188 189100
rect 381504 189060 382188 189088
rect 381504 189048 381510 189060
rect 382182 189048 382188 189060
rect 382240 189048 382246 189100
rect 385494 189048 385500 189100
rect 385552 189088 385558 189100
rect 386230 189088 386236 189100
rect 385552 189060 386236 189088
rect 385552 189048 385558 189060
rect 386230 189048 386236 189060
rect 386288 189048 386294 189100
rect 387978 189048 387984 189100
rect 388036 189088 388042 189100
rect 388990 189088 388996 189100
rect 388036 189060 388996 189088
rect 388036 189048 388042 189060
rect 388990 189048 388996 189060
rect 389048 189048 389054 189100
rect 400398 189048 400404 189100
rect 400456 189088 400462 189100
rect 401502 189088 401508 189100
rect 400456 189060 401508 189088
rect 400456 189048 400462 189060
rect 401502 189048 401508 189060
rect 401560 189048 401566 189100
rect 402054 189048 402060 189100
rect 402112 189088 402118 189100
rect 402882 189088 402888 189100
rect 402112 189060 402888 189088
rect 402112 189048 402118 189060
rect 402882 189048 402888 189060
rect 402940 189048 402946 189100
rect 404538 189048 404544 189100
rect 404596 189088 404602 189100
rect 405550 189088 405556 189100
rect 404596 189060 405556 189088
rect 404596 189048 404602 189060
rect 405550 189048 405556 189060
rect 405608 189048 405614 189100
rect 410242 189048 410248 189100
rect 410300 189088 410306 189100
rect 411162 189088 411168 189100
rect 410300 189060 411168 189088
rect 410300 189048 410306 189060
rect 411162 189048 411168 189060
rect 411220 189048 411226 189100
rect 414382 189048 414388 189100
rect 414440 189088 414446 189100
rect 416038 189088 416044 189100
rect 414440 189060 416044 189088
rect 414440 189048 414446 189060
rect 416038 189048 416044 189060
rect 416096 189048 416102 189100
rect 418522 189048 418528 189100
rect 418580 189088 418586 189100
rect 420178 189088 420184 189100
rect 418580 189060 420184 189088
rect 418580 189048 418586 189060
rect 420178 189048 420184 189060
rect 420236 189048 420242 189100
rect 421006 189048 421012 189100
rect 421064 189088 421070 189100
rect 422110 189088 422116 189100
rect 421064 189060 422116 189088
rect 421064 189048 421070 189060
rect 422110 189048 422116 189060
rect 422168 189048 422174 189100
rect 422662 189048 422668 189100
rect 422720 189088 422726 189100
rect 423490 189088 423496 189100
rect 422720 189060 423496 189088
rect 422720 189048 422726 189060
rect 423490 189048 423496 189060
rect 423548 189048 423554 189100
rect 426802 189048 426808 189100
rect 426860 189088 426866 189100
rect 427630 189088 427636 189100
rect 426860 189060 427636 189088
rect 426860 189048 426866 189060
rect 427630 189048 427636 189060
rect 427688 189048 427694 189100
rect 428366 189048 428372 189100
rect 428424 189088 428430 189100
rect 429102 189088 429108 189100
rect 428424 189060 429108 189088
rect 428424 189048 428430 189060
rect 429102 189048 429108 189060
rect 429160 189048 429166 189100
rect 430850 189048 430856 189100
rect 430908 189088 430914 189100
rect 431770 189088 431776 189100
rect 430908 189060 431776 189088
rect 430908 189048 430914 189060
rect 431770 189048 431776 189060
rect 431828 189048 431834 189100
rect 436646 189048 436652 189100
rect 436704 189088 436710 189100
rect 437382 189088 437388 189100
rect 436704 189060 437388 189088
rect 436704 189048 436710 189060
rect 437382 189048 437388 189060
rect 437440 189048 437446 189100
rect 443270 189048 443276 189100
rect 443328 189088 443334 189100
rect 444190 189088 444196 189100
rect 443328 189060 444196 189088
rect 443328 189048 443334 189060
rect 444190 189048 444196 189060
rect 444248 189048 444254 189100
rect 444926 189048 444932 189100
rect 444984 189088 444990 189100
rect 445662 189088 445668 189100
rect 444984 189060 445668 189088
rect 444984 189048 444990 189060
rect 445662 189048 445668 189060
rect 445720 189048 445726 189100
rect 447410 189048 447416 189100
rect 447468 189088 447474 189100
rect 448422 189088 448428 189100
rect 447468 189060 448428 189088
rect 447468 189048 447474 189060
rect 448422 189048 448428 189060
rect 448480 189048 448486 189100
rect 449894 189048 449900 189100
rect 449952 189088 449958 189100
rect 451182 189088 451188 189100
rect 449952 189060 451188 189088
rect 449952 189048 449958 189060
rect 451182 189048 451188 189060
rect 451240 189048 451246 189100
rect 220722 188300 220728 188352
rect 220780 188340 220786 188352
rect 251174 188340 251180 188352
rect 220780 188312 251180 188340
rect 220780 188300 220786 188312
rect 251174 188300 251180 188312
rect 251232 188300 251238 188352
rect 252738 188300 252744 188352
rect 252796 188340 252802 188352
rect 296714 188340 296720 188352
rect 252796 188312 296720 188340
rect 252796 188300 252802 188312
rect 296714 188300 296720 188312
rect 296772 188300 296778 188352
rect 388806 188300 388812 188352
rect 388864 188340 388870 188352
rect 494054 188340 494060 188352
rect 388864 188312 494060 188340
rect 388864 188300 388870 188312
rect 494054 188300 494060 188312
rect 494112 188300 494118 188352
rect 235442 186940 235448 186992
rect 235500 186980 235506 186992
rect 271874 186980 271880 186992
rect 235500 186952 271880 186980
rect 235500 186940 235506 186952
rect 271874 186940 271880 186952
rect 271932 186940 271938 186992
rect 271966 186940 271972 186992
rect 272024 186980 272030 186992
rect 322934 186980 322940 186992
rect 272024 186952 322940 186980
rect 272024 186940 272030 186952
rect 322934 186940 322940 186952
rect 322992 186940 322998 186992
rect 393774 186940 393780 186992
rect 393832 186980 393838 186992
rect 500954 186980 500960 186992
rect 393832 186952 500960 186980
rect 393832 186940 393838 186952
rect 500954 186940 500960 186952
rect 501012 186940 501018 186992
rect 147674 185580 147680 185632
rect 147732 185620 147738 185632
rect 148502 185620 148508 185632
rect 147732 185592 148508 185620
rect 147732 185580 147738 185592
rect 148502 185580 148508 185592
rect 148560 185580 148566 185632
rect 150434 185580 150440 185632
rect 150492 185620 150498 185632
rect 151078 185620 151084 185632
rect 150492 185592 151084 185620
rect 150492 185580 150498 185592
rect 151078 185580 151084 185592
rect 151136 185580 151142 185632
rect 396258 185580 396264 185632
rect 396316 185620 396322 185632
rect 503714 185620 503720 185632
rect 396316 185592 503720 185620
rect 396316 185580 396322 185592
rect 503714 185580 503720 185592
rect 503772 185580 503778 185632
rect 401226 184152 401232 184204
rect 401284 184192 401290 184204
rect 511994 184192 512000 184204
rect 401284 184164 512000 184192
rect 401284 184152 401290 184164
rect 511994 184152 512000 184164
rect 512052 184152 512058 184204
rect 135530 183472 135536 183524
rect 135588 183512 135594 183524
rect 135622 183512 135628 183524
rect 135588 183484 135628 183512
rect 135588 183472 135594 183484
rect 135622 183472 135628 183484
rect 135680 183472 135686 183524
rect 406102 182792 406108 182844
rect 406160 182832 406166 182844
rect 518894 182832 518900 182844
rect 406160 182804 518900 182832
rect 406160 182792 406166 182804
rect 518894 182792 518900 182804
rect 518952 182792 518958 182844
rect 453666 182112 453672 182164
rect 453724 182152 453730 182164
rect 580166 182152 580172 182164
rect 453724 182124 580172 182152
rect 453724 182112 453730 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 142154 181432 142160 181484
rect 142212 181472 142218 181484
rect 142798 181472 142804 181484
rect 142212 181444 142804 181472
rect 142212 181432 142218 181444
rect 142798 181432 142804 181444
rect 142856 181432 142862 181484
rect 367370 181432 367376 181484
rect 367428 181472 367434 181484
rect 462314 181472 462320 181484
rect 367428 181444 462320 181472
rect 367428 181432 367434 181444
rect 462314 181432 462320 181444
rect 462372 181432 462378 181484
rect 146294 180888 146300 180940
rect 146352 180928 146358 180940
rect 146846 180928 146852 180940
rect 146352 180900 146852 180928
rect 146352 180888 146358 180900
rect 146846 180888 146852 180900
rect 146904 180888 146910 180940
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 13078 180792 13084 180804
rect 3292 180764 13084 180792
rect 3292 180752 3298 180764
rect 13078 180752 13084 180764
rect 13136 180752 13142 180804
rect 409690 180072 409696 180124
rect 409748 180112 409754 180124
rect 521654 180112 521660 180124
rect 409748 180084 521660 180112
rect 409748 180072 409754 180084
rect 521654 180072 521660 180084
rect 521712 180072 521718 180124
rect 223482 178644 223488 178696
rect 223540 178684 223546 178696
rect 252554 178684 252560 178696
rect 223540 178656 252560 178684
rect 223540 178644 223546 178656
rect 252554 178644 252560 178656
rect 252612 178644 252618 178696
rect 259270 178644 259276 178696
rect 259328 178684 259334 178696
rect 304994 178684 305000 178696
rect 259328 178656 305000 178684
rect 259328 178644 259334 178656
rect 304994 178644 305000 178656
rect 305052 178644 305058 178696
rect 318610 178644 318616 178696
rect 318668 178684 318674 178696
rect 390554 178684 390560 178696
rect 318668 178656 390560 178684
rect 318668 178644 318674 178656
rect 390554 178644 390560 178656
rect 390612 178644 390618 178696
rect 413830 178644 413836 178696
rect 413888 178684 413894 178696
rect 528554 178684 528560 178696
rect 413888 178656 528560 178684
rect 413888 178644 413894 178656
rect 528554 178644 528560 178656
rect 528612 178644 528618 178696
rect 227530 177284 227536 177336
rect 227588 177324 227594 177336
rect 259454 177324 259460 177336
rect 227588 177296 259460 177324
rect 227588 177284 227594 177296
rect 259454 177284 259460 177296
rect 259512 177284 259518 177336
rect 335170 177284 335176 177336
rect 335228 177324 335234 177336
rect 415394 177324 415400 177336
rect 335228 177296 415400 177324
rect 335228 177284 335234 177296
rect 415394 177284 415400 177296
rect 415452 177284 415458 177336
rect 420178 177284 420184 177336
rect 420236 177324 420242 177336
rect 536834 177324 536840 177336
rect 420236 177296 536840 177324
rect 420236 177284 420242 177296
rect 536834 177284 536840 177296
rect 536892 177284 536898 177336
rect 422110 175924 422116 175976
rect 422168 175964 422174 175976
rect 539594 175964 539600 175976
rect 422168 175936 539600 175964
rect 422168 175924 422174 175936
rect 539594 175924 539600 175936
rect 539652 175924 539658 175976
rect 426250 174496 426256 174548
rect 426308 174536 426314 174548
rect 546494 174536 546500 174548
rect 426308 174508 546500 174536
rect 426308 174496 426314 174508
rect 546494 174496 546500 174508
rect 546552 174496 546558 174548
rect 143902 173884 143908 173936
rect 143960 173924 143966 173936
rect 144178 173924 144184 173936
rect 143960 173896 144184 173924
rect 143960 173884 143966 173896
rect 144178 173884 144184 173896
rect 144236 173884 144242 173936
rect 431770 173136 431776 173188
rect 431828 173176 431834 173188
rect 554774 173176 554780 173188
rect 431828 173148 554780 173176
rect 431828 173136 431834 173148
rect 554774 173136 554780 173148
rect 554832 173136 554838 173188
rect 434530 171776 434536 171828
rect 434588 171816 434594 171828
rect 557534 171816 557540 171828
rect 434588 171788 557540 171816
rect 434588 171776 434594 171788
rect 557534 171776 557540 171788
rect 557592 171776 557598 171828
rect 453574 171028 453580 171080
rect 453632 171068 453638 171080
rect 580166 171068 580172 171080
rect 453632 171040 580172 171068
rect 453632 171028 453638 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 438670 168988 438676 169040
rect 438728 169028 438734 169040
rect 564434 169028 564440 169040
rect 438728 169000 564440 169028
rect 438728 168988 438734 169000
rect 564434 168988 564440 169000
rect 564492 168988 564498 169040
rect 444190 167628 444196 167680
rect 444248 167668 444254 167680
rect 571334 167668 571340 167680
rect 444248 167640 571340 167668
rect 444248 167628 444254 167640
rect 571334 167628 571340 167640
rect 571392 167628 571398 167680
rect 354490 166268 354496 166320
rect 354548 166308 354554 166320
rect 442994 166308 443000 166320
rect 354548 166280 443000 166308
rect 354548 166268 354554 166280
rect 442994 166268 443000 166280
rect 443052 166268 443058 166320
rect 446950 166268 446956 166320
rect 447008 166308 447014 166320
rect 575474 166308 575480 166320
rect 447008 166280 575480 166308
rect 447008 166268 447014 166280
rect 575474 166268 575480 166280
rect 575532 166268 575538 166320
rect 448330 164840 448336 164892
rect 448388 164880 448394 164892
rect 578878 164880 578884 164892
rect 448388 164852 578884 164880
rect 448388 164840 448394 164852
rect 578878 164840 578884 164852
rect 578936 164840 578942 164892
rect 143626 164160 143632 164212
rect 143684 164200 143690 164212
rect 143810 164200 143816 164212
rect 143684 164172 143816 164200
rect 143684 164160 143690 164172
rect 143810 164160 143816 164172
rect 143868 164160 143874 164212
rect 364150 163480 364156 163532
rect 364208 163520 364214 163532
rect 458174 163520 458180 163532
rect 364208 163492 458180 163520
rect 364208 163480 364214 163492
rect 458174 163480 458180 163492
rect 458232 163480 458238 163532
rect 366910 162120 366916 162172
rect 366968 162160 366974 162172
rect 460934 162160 460940 162172
rect 366968 162132 460940 162160
rect 366968 162120 366974 162132
rect 460934 162120 460940 162132
rect 460992 162120 460998 162172
rect 376570 160692 376576 160744
rect 376628 160732 376634 160744
rect 476114 160732 476120 160744
rect 376628 160704 476120 160732
rect 376628 160692 376634 160704
rect 476114 160692 476120 160704
rect 476172 160692 476178 160744
rect 381538 159332 381544 159384
rect 381596 159372 381602 159384
rect 478874 159372 478880 159384
rect 381596 159344 478880 159372
rect 381596 159332 381602 159344
rect 478874 159332 478880 159344
rect 478932 159332 478938 159384
rect 471238 158652 471244 158704
rect 471296 158692 471302 158704
rect 579798 158692 579804 158704
rect 471296 158664 579804 158692
rect 471296 158652 471302 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 365622 157972 365628 158024
rect 365680 158012 365686 158024
rect 459646 158012 459652 158024
rect 365680 157984 459652 158012
rect 365680 157972 365686 157984
rect 459646 157972 459652 157984
rect 459704 157972 459710 158024
rect 387058 156612 387064 156664
rect 387116 156652 387122 156664
rect 484394 156652 484400 156664
rect 387116 156624 484400 156652
rect 387116 156612 387122 156624
rect 484394 156612 484400 156624
rect 484452 156612 484458 156664
rect 384942 155184 384948 155236
rect 385000 155224 385006 155236
rect 487154 155224 487160 155236
rect 385000 155196 487160 155224
rect 385000 155184 385006 155196
rect 487154 155184 487160 155196
rect 487212 155184 487218 155236
rect 135346 154544 135352 154556
rect 135307 154516 135352 154544
rect 135346 154504 135352 154516
rect 135404 154504 135410 154556
rect 393130 153824 393136 153876
rect 393188 153864 393194 153876
rect 498194 153864 498200 153876
rect 393188 153836 498200 153864
rect 393188 153824 393194 153836
rect 498194 153824 498200 153836
rect 498252 153824 498258 153876
rect 397362 152464 397368 152516
rect 397420 152504 397426 152516
rect 505094 152504 505100 152516
rect 397420 152476 505100 152504
rect 397420 152464 397426 152476
rect 505094 152464 505100 152476
rect 505152 152464 505158 152516
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 129274 151756 129280 151768
rect 3200 151728 129280 151756
rect 3200 151716 3206 151728
rect 129274 151716 129280 151728
rect 129332 151716 129338 151768
rect 405550 151036 405556 151088
rect 405608 151076 405614 151088
rect 516134 151076 516140 151088
rect 405608 151048 516140 151076
rect 405608 151036 405614 151048
rect 516134 151036 516140 151048
rect 516192 151036 516198 151088
rect 416038 149676 416044 149728
rect 416096 149716 416102 149728
rect 529934 149716 529940 149728
rect 416096 149688 529940 149716
rect 416096 149676 416102 149688
rect 529934 149676 529940 149688
rect 529992 149676 529998 149728
rect 417970 148316 417976 148368
rect 418028 148356 418034 148368
rect 534074 148356 534080 148368
rect 418028 148328 534080 148356
rect 418028 148316 418034 148328
rect 534074 148316 534080 148328
rect 534132 148316 534138 148368
rect 135349 147611 135407 147617
rect 135349 147577 135361 147611
rect 135395 147608 135407 147611
rect 135438 147608 135444 147620
rect 135395 147580 135444 147608
rect 135395 147577 135407 147580
rect 135349 147571 135407 147577
rect 135438 147568 135444 147580
rect 135496 147568 135502 147620
rect 427630 146888 427636 146940
rect 427688 146928 427694 146940
rect 547874 146928 547880 146940
rect 427688 146900 547880 146928
rect 427688 146888 427694 146900
rect 547874 146888 547880 146900
rect 547932 146888 547938 146940
rect 430390 145528 430396 145580
rect 430448 145568 430454 145580
rect 552014 145568 552020 145580
rect 430448 145540 552020 145568
rect 430448 145528 430454 145540
rect 552014 145528 552020 145540
rect 552072 145528 552078 145580
rect 437382 144168 437388 144220
rect 437440 144208 437446 144220
rect 563054 144208 563060 144220
rect 437440 144180 563060 144208
rect 437440 144168 437446 144180
rect 563054 144168 563060 144180
rect 563112 144168 563118 144220
rect 135438 143488 135444 143540
rect 135496 143528 135502 143540
rect 135533 143531 135591 143537
rect 135533 143528 135545 143531
rect 135496 143500 135545 143528
rect 135496 143488 135502 143500
rect 135533 143497 135545 143500
rect 135579 143497 135591 143531
rect 143810 143528 143816 143540
rect 143771 143500 143816 143528
rect 135533 143491 135591 143497
rect 143810 143488 143816 143500
rect 143868 143488 143874 143540
rect 440050 142808 440056 142860
rect 440108 142848 440114 142860
rect 565814 142848 565820 142860
rect 440108 142820 565820 142848
rect 440108 142808 440114 142820
rect 565814 142808 565820 142820
rect 565872 142808 565878 142860
rect 442810 141380 442816 141432
rect 442868 141420 442874 141432
rect 569954 141420 569960 141432
rect 442868 141392 569960 141420
rect 442868 141380 442874 141392
rect 569954 141380 569960 141392
rect 570012 141380 570018 141432
rect 371050 140020 371056 140072
rect 371108 140060 371114 140072
rect 466454 140060 466460 140072
rect 371108 140032 466460 140060
rect 371108 140020 371114 140032
rect 466454 140020 466460 140032
rect 466512 140020 466518 140072
rect 380710 138660 380716 138712
rect 380768 138700 380774 138712
rect 480254 138700 480260 138712
rect 380768 138672 480260 138700
rect 380768 138660 380774 138672
rect 480254 138660 480260 138672
rect 480312 138660 480318 138712
rect 386230 137232 386236 137284
rect 386288 137272 386294 137284
rect 488534 137272 488540 137284
rect 386288 137244 488540 137272
rect 386288 137232 386294 137244
rect 488534 137232 488540 137244
rect 488592 137232 488598 137284
rect 3418 136484 3424 136536
rect 3476 136524 3482 136536
rect 8938 136524 8944 136536
rect 3476 136496 8944 136524
rect 3476 136484 3482 136496
rect 8938 136484 8944 136496
rect 8996 136484 9002 136536
rect 390370 135872 390376 135924
rect 390428 135912 390434 135924
rect 495434 135912 495440 135924
rect 390428 135884 495440 135912
rect 390428 135872 390434 135884
rect 495434 135872 495440 135884
rect 495492 135872 495498 135924
rect 457438 135192 457444 135244
rect 457496 135232 457502 135244
rect 580166 135232 580172 135244
rect 457496 135204 580172 135232
rect 457496 135192 457502 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 398650 133152 398656 133204
rect 398708 133192 398714 133204
rect 506474 133192 506480 133204
rect 398708 133164 506480 133192
rect 398708 133152 398714 133164
rect 506474 133152 506480 133164
rect 506532 133152 506538 133204
rect 401502 131724 401508 131776
rect 401560 131764 401566 131776
rect 510614 131764 510620 131776
rect 401560 131736 510620 131764
rect 401560 131724 401566 131736
rect 510614 131724 510620 131736
rect 510672 131724 510678 131776
rect 135533 131495 135591 131501
rect 135533 131461 135545 131495
rect 135579 131492 135591 131495
rect 135622 131492 135628 131504
rect 135579 131464 135628 131492
rect 135579 131461 135591 131464
rect 135533 131455 135591 131461
rect 135622 131452 135628 131464
rect 135680 131452 135686 131504
rect 402790 130364 402796 130416
rect 402848 130404 402854 130416
rect 513374 130404 513380 130416
rect 402848 130376 513380 130404
rect 402848 130364 402854 130376
rect 513374 130364 513380 130376
rect 513432 130364 513438 130416
rect 415302 129004 415308 129056
rect 415360 129044 415366 129056
rect 531314 129044 531320 129056
rect 415360 129016 531320 129044
rect 415360 129004 415366 129016
rect 531314 129004 531320 129016
rect 531372 129004 531378 129056
rect 143810 128296 143816 128308
rect 143771 128268 143816 128296
rect 143810 128256 143816 128268
rect 143868 128256 143874 128308
rect 423490 127576 423496 127628
rect 423548 127616 423554 127628
rect 542354 127616 542360 127628
rect 423548 127588 542360 127616
rect 423548 127576 423554 127588
rect 542354 127576 542360 127588
rect 542412 127576 542418 127628
rect 433242 126216 433248 126268
rect 433300 126256 433306 126268
rect 556154 126256 556160 126268
rect 433300 126228 556160 126256
rect 433300 126216 433306 126228
rect 556154 126216 556160 126228
rect 556212 126216 556218 126268
rect 435910 124856 435916 124908
rect 435968 124896 435974 124908
rect 560294 124896 560300 124908
rect 435968 124868 560300 124896
rect 435968 124856 435974 124868
rect 560294 124856 560300 124868
rect 560352 124856 560358 124908
rect 135622 124108 135628 124160
rect 135680 124148 135686 124160
rect 135806 124148 135812 124160
rect 135680 124120 135812 124148
rect 135680 124108 135686 124120
rect 135806 124108 135812 124120
rect 135864 124108 135870 124160
rect 453482 124108 453488 124160
rect 453540 124148 453546 124160
rect 580166 124148 580172 124160
rect 453540 124120 580172 124148
rect 453540 124108 453546 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 10318 122788 10324 122800
rect 3476 122760 10324 122788
rect 3476 122748 3482 122760
rect 10318 122748 10324 122760
rect 10376 122748 10382 122800
rect 135625 122791 135683 122797
rect 135625 122757 135637 122791
rect 135671 122788 135683 122791
rect 135806 122788 135812 122800
rect 135671 122760 135812 122788
rect 135671 122757 135683 122760
rect 135625 122751 135683 122757
rect 135806 122748 135812 122760
rect 135864 122748 135870 122800
rect 351730 113772 351736 113824
rect 351788 113812 351794 113824
rect 438854 113812 438860 113824
rect 351788 113784 438860 113812
rect 351788 113772 351794 113784
rect 438854 113772 438860 113784
rect 438912 113772 438918 113824
rect 343542 112412 343548 112464
rect 343600 112452 343606 112464
rect 427814 112452 427820 112464
rect 343600 112424 427820 112452
rect 343600 112412 343606 112424
rect 427814 112412 427820 112424
rect 427872 112412 427878 112464
rect 469858 111732 469864 111784
rect 469916 111772 469922 111784
rect 579798 111772 579804 111784
rect 469916 111744 579804 111772
rect 469916 111732 469922 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 372430 111052 372436 111104
rect 372488 111092 372494 111104
rect 469214 111092 469220 111104
rect 372488 111064 469220 111092
rect 372488 111052 372494 111064
rect 469214 111052 469220 111064
rect 469272 111052 469278 111104
rect 333790 109692 333796 109744
rect 333848 109732 333854 109744
rect 414014 109732 414020 109744
rect 333848 109704 414020 109732
rect 333848 109692 333854 109704
rect 414014 109692 414020 109704
rect 414072 109692 414078 109744
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 129182 108984 129188 108996
rect 3292 108956 129188 108984
rect 3292 108944 3298 108956
rect 129182 108944 129188 108956
rect 129240 108944 129246 108996
rect 331030 108264 331036 108316
rect 331088 108304 331094 108316
rect 409874 108304 409880 108316
rect 331088 108276 409880 108304
rect 331088 108264 331094 108276
rect 409874 108264 409880 108276
rect 409932 108264 409938 108316
rect 342070 106904 342076 106956
rect 342128 106944 342134 106956
rect 425054 106944 425060 106956
rect 342128 106916 425060 106944
rect 342128 106904 342134 106916
rect 425054 106904 425060 106916
rect 425112 106904 425118 106956
rect 135622 106196 135628 106208
rect 135583 106168 135628 106196
rect 135622 106156 135628 106168
rect 135680 106156 135686 106208
rect 349062 105544 349068 105596
rect 349120 105584 349126 105596
rect 434714 105584 434720 105596
rect 349120 105556 434720 105584
rect 349120 105544 349126 105556
rect 434714 105544 434720 105556
rect 434772 105544 434778 105596
rect 135622 104836 135628 104848
rect 135583 104808 135628 104836
rect 135622 104796 135628 104808
rect 135680 104796 135686 104848
rect 331858 104116 331864 104168
rect 331916 104156 331922 104168
rect 408494 104156 408500 104168
rect 331916 104128 408500 104156
rect 331916 104116 331922 104128
rect 408494 104116 408500 104128
rect 408552 104116 408558 104168
rect 339310 102756 339316 102808
rect 339368 102796 339374 102808
rect 420914 102796 420920 102808
rect 339368 102768 420920 102796
rect 339368 102756 339374 102768
rect 420914 102756 420920 102768
rect 420972 102756 420978 102808
rect 336642 101396 336648 101448
rect 336700 101436 336706 101448
rect 416774 101436 416780 101448
rect 336700 101408 416780 101436
rect 336700 101396 336706 101408
rect 416774 101396 416780 101408
rect 416832 101396 416838 101448
rect 329742 99968 329748 100020
rect 329800 100008 329806 100020
rect 407114 100008 407120 100020
rect 329800 99980 407120 100008
rect 329800 99968 329806 99980
rect 407114 99968 407120 99980
rect 407172 99968 407178 100020
rect 326890 98608 326896 98660
rect 326948 98648 326954 98660
rect 402974 98648 402980 98660
rect 326948 98620 402980 98648
rect 326948 98608 326954 98620
rect 402974 98608 402980 98620
rect 403032 98608 403038 98660
rect 324222 97248 324228 97300
rect 324280 97288 324286 97300
rect 400214 97288 400220 97300
rect 324280 97260 400220 97288
rect 324280 97248 324286 97260
rect 400214 97248 400220 97260
rect 400272 97248 400278 97300
rect 321370 95888 321376 95940
rect 321428 95928 321434 95940
rect 396074 95928 396080 95940
rect 321428 95900 396080 95928
rect 321428 95888 321434 95900
rect 396074 95888 396080 95900
rect 396132 95888 396138 95940
rect 318702 94460 318708 94512
rect 318760 94500 318766 94512
rect 391934 94500 391940 94512
rect 318760 94472 391940 94500
rect 318760 94460 318766 94472
rect 391934 94460 391940 94472
rect 391992 94460 391998 94512
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 15838 93820 15844 93832
rect 3476 93792 15844 93820
rect 3476 93780 3482 93792
rect 15838 93780 15844 93792
rect 15896 93780 15902 93832
rect 317230 93100 317236 93152
rect 317288 93140 317294 93152
rect 389174 93140 389180 93152
rect 317288 93112 389180 93140
rect 317288 93100 317294 93112
rect 389174 93100 389180 93112
rect 389232 93100 389238 93152
rect 314470 91740 314476 91792
rect 314528 91780 314534 91792
rect 385034 91780 385040 91792
rect 314528 91752 385040 91780
rect 314528 91740 314534 91752
rect 385034 91740 385040 91752
rect 385092 91740 385098 91792
rect 328362 90312 328368 90364
rect 328420 90352 328426 90364
rect 405734 90352 405740 90364
rect 328420 90324 405740 90352
rect 328420 90312 328426 90324
rect 405734 90312 405740 90324
rect 405792 90312 405798 90364
rect 135530 89632 135536 89684
rect 135588 89672 135594 89684
rect 135625 89675 135683 89681
rect 135625 89672 135637 89675
rect 135588 89644 135637 89672
rect 135588 89632 135594 89644
rect 135625 89641 135637 89644
rect 135671 89641 135683 89675
rect 135625 89635 135683 89641
rect 311802 88952 311808 89004
rect 311860 88992 311866 89004
rect 382274 88992 382280 89004
rect 311860 88964 382280 88992
rect 311860 88952 311866 88964
rect 382274 88952 382280 88964
rect 382332 88952 382338 89004
rect 473998 88272 474004 88324
rect 474056 88312 474062 88324
rect 580166 88312 580172 88324
rect 474056 88284 580172 88312
rect 474056 88272 474062 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 375190 87592 375196 87644
rect 375248 87632 375254 87644
rect 473354 87632 473360 87644
rect 375248 87604 473360 87632
rect 375248 87592 375254 87604
rect 473354 87592 473360 87604
rect 473412 87592 473418 87644
rect 135438 86912 135444 86964
rect 135496 86952 135502 86964
rect 135714 86952 135720 86964
rect 135496 86924 135720 86952
rect 135496 86912 135502 86924
rect 135714 86912 135720 86924
rect 135772 86912 135778 86964
rect 143629 86955 143687 86961
rect 143629 86921 143641 86955
rect 143675 86952 143687 86955
rect 143718 86952 143724 86964
rect 143675 86924 143724 86952
rect 143675 86921 143687 86924
rect 143629 86915 143687 86921
rect 143718 86912 143724 86924
rect 143776 86912 143782 86964
rect 304810 86232 304816 86284
rect 304868 86272 304874 86284
rect 371234 86272 371240 86284
rect 304868 86244 371240 86272
rect 304868 86232 304874 86244
rect 371234 86232 371240 86244
rect 371292 86232 371298 86284
rect 408402 86232 408408 86284
rect 408460 86272 408466 86284
rect 520274 86272 520280 86284
rect 408460 86244 520280 86272
rect 408460 86232 408466 86244
rect 520274 86232 520280 86244
rect 520332 86232 520338 86284
rect 135714 85524 135720 85536
rect 135675 85496 135720 85524
rect 135714 85484 135720 85496
rect 135772 85484 135778 85536
rect 307662 84804 307668 84856
rect 307720 84844 307726 84856
rect 373994 84844 374000 84856
rect 307720 84816 374000 84844
rect 307720 84804 307726 84816
rect 373994 84804 374000 84816
rect 374052 84804 374058 84856
rect 427722 84804 427728 84856
rect 427780 84844 427786 84856
rect 549254 84844 549260 84856
rect 427780 84816 549260 84844
rect 427780 84804 427786 84816
rect 549254 84804 549260 84816
rect 549312 84804 549318 84856
rect 302142 83444 302148 83496
rect 302200 83484 302206 83496
rect 367094 83484 367100 83496
rect 302200 83456 367100 83484
rect 302200 83444 302206 83456
rect 367094 83444 367100 83456
rect 367152 83444 367158 83496
rect 420822 83444 420828 83496
rect 420880 83484 420886 83496
rect 538214 83484 538220 83496
rect 420880 83456 538220 83484
rect 420880 83444 420886 83456
rect 538214 83444 538220 83456
rect 538272 83444 538278 83496
rect 299290 82084 299296 82136
rect 299348 82124 299354 82136
rect 364334 82124 364340 82136
rect 299348 82096 364340 82124
rect 299348 82084 299354 82096
rect 364334 82084 364340 82096
rect 364392 82084 364398 82136
rect 395982 82084 395988 82136
rect 396040 82124 396046 82136
rect 502334 82124 502340 82136
rect 396040 82096 502340 82124
rect 396040 82084 396046 82096
rect 502334 82084 502340 82096
rect 502392 82084 502398 82136
rect 295242 80656 295248 80708
rect 295300 80696 295306 80708
rect 356054 80696 356060 80708
rect 295300 80668 356060 80696
rect 295300 80656 295306 80668
rect 356054 80656 356060 80668
rect 356112 80656 356118 80708
rect 362770 80656 362776 80708
rect 362828 80696 362834 80708
rect 455414 80696 455420 80708
rect 362828 80668 455420 80696
rect 362828 80656 362834 80668
rect 455414 80656 455420 80668
rect 455472 80656 455478 80708
rect 3418 79976 3424 80028
rect 3476 80016 3482 80028
rect 14458 80016 14464 80028
rect 3476 79988 14464 80016
rect 3476 79976 3482 79988
rect 14458 79976 14464 79988
rect 14516 79976 14522 80028
rect 292390 79296 292396 79348
rect 292448 79336 292454 79348
rect 353294 79336 353300 79348
rect 292448 79308 353300 79336
rect 292448 79296 292454 79308
rect 353294 79296 353300 79308
rect 353352 79296 353358 79348
rect 355870 79296 355876 79348
rect 355928 79336 355934 79348
rect 444374 79336 444380 79348
rect 355928 79308 444380 79336
rect 355928 79296 355934 79308
rect 444374 79296 444380 79308
rect 444432 79296 444438 79348
rect 445662 79296 445668 79348
rect 445720 79336 445726 79348
rect 574094 79336 574100 79348
rect 445720 79308 574100 79336
rect 445720 79296 445726 79308
rect 574094 79296 574100 79308
rect 574152 79296 574158 79348
rect 289722 77936 289728 77988
rect 289780 77976 289786 77988
rect 349154 77976 349160 77988
rect 289780 77948 349160 77976
rect 289780 77936 289786 77948
rect 349154 77936 349160 77948
rect 349212 77936 349218 77988
rect 360010 77936 360016 77988
rect 360068 77976 360074 77988
rect 451274 77976 451280 77988
rect 360068 77948 451280 77976
rect 360068 77936 360074 77948
rect 451274 77936 451280 77948
rect 451332 77936 451338 77988
rect 135714 77296 135720 77308
rect 135675 77268 135720 77296
rect 135714 77256 135720 77268
rect 135772 77256 135778 77308
rect 143626 77296 143632 77308
rect 143587 77268 143632 77296
rect 143626 77256 143632 77268
rect 143684 77256 143690 77308
rect 453390 77188 453396 77240
rect 453448 77228 453454 77240
rect 580166 77228 580172 77240
rect 453448 77200 580172 77228
rect 453448 77188 453454 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 286870 76508 286876 76560
rect 286928 76548 286934 76560
rect 346394 76548 346400 76560
rect 286928 76520 346400 76548
rect 286928 76508 286934 76520
rect 346394 76508 346400 76520
rect 346452 76508 346458 76560
rect 353202 76508 353208 76560
rect 353260 76548 353266 76560
rect 441614 76548 441620 76560
rect 353260 76520 441620 76548
rect 353260 76508 353266 76520
rect 441614 76508 441620 76520
rect 441672 76508 441678 76560
rect 284110 75148 284116 75200
rect 284168 75188 284174 75200
rect 342254 75188 342260 75200
rect 284168 75160 342260 75188
rect 284168 75148 284174 75160
rect 342254 75148 342260 75160
rect 342312 75148 342318 75200
rect 347682 75148 347688 75200
rect 347740 75188 347746 75200
rect 433334 75188 433340 75200
rect 347740 75160 433340 75188
rect 347740 75148 347746 75160
rect 433334 75148 433340 75160
rect 433392 75148 433398 75200
rect 279970 73788 279976 73840
rect 280028 73828 280034 73840
rect 335354 73828 335360 73840
rect 280028 73800 335360 73828
rect 280028 73788 280034 73800
rect 335354 73788 335360 73800
rect 335412 73788 335418 73840
rect 346210 73788 346216 73840
rect 346268 73828 346274 73840
rect 430574 73828 430580 73840
rect 346268 73800 430580 73828
rect 346268 73788 346274 73800
rect 430574 73788 430580 73800
rect 430632 73788 430638 73840
rect 282730 72428 282736 72480
rect 282788 72468 282794 72480
rect 339494 72468 339500 72480
rect 282788 72440 339500 72468
rect 282788 72428 282794 72440
rect 339494 72428 339500 72440
rect 339552 72428 339558 72480
rect 344278 72428 344284 72480
rect 344336 72468 344342 72480
rect 426434 72468 426440 72480
rect 344336 72440 426440 72468
rect 344336 72428 344342 72440
rect 426434 72428 426440 72440
rect 426492 72428 426498 72480
rect 442902 72428 442908 72480
rect 442960 72468 442966 72480
rect 571426 72468 571432 72480
rect 442960 72440 571432 72468
rect 442960 72428 442966 72440
rect 571426 72428 571432 72440
rect 571484 72428 571490 72480
rect 277302 71000 277308 71052
rect 277360 71040 277366 71052
rect 331214 71040 331220 71052
rect 277360 71012 331220 71040
rect 277360 71000 277366 71012
rect 331214 71000 331220 71012
rect 331272 71000 331278 71052
rect 340782 71000 340788 71052
rect 340840 71040 340846 71052
rect 423674 71040 423680 71052
rect 340840 71012 423680 71040
rect 340840 71000 340846 71012
rect 423674 71000 423680 71012
rect 423732 71000 423738 71052
rect 440142 71000 440148 71052
rect 440200 71040 440206 71052
rect 567194 71040 567200 71052
rect 440200 71012 567200 71040
rect 440200 71000 440206 71012
rect 567194 71000 567200 71012
rect 567252 71000 567258 71052
rect 274450 69640 274456 69692
rect 274508 69680 274514 69692
rect 328454 69680 328460 69692
rect 274508 69652 328460 69680
rect 274508 69640 274514 69652
rect 328454 69640 328460 69652
rect 328512 69640 328518 69692
rect 337930 69640 337936 69692
rect 337988 69680 337994 69692
rect 419534 69680 419540 69692
rect 337988 69652 419540 69680
rect 337988 69640 337994 69652
rect 419534 69640 419540 69652
rect 419592 69640 419598 69692
rect 438762 69640 438768 69692
rect 438820 69680 438826 69692
rect 563146 69680 563152 69692
rect 438820 69652 563152 69680
rect 438820 69640 438826 69652
rect 563146 69640 563152 69652
rect 563204 69640 563210 69692
rect 271782 68280 271788 68332
rect 271840 68320 271846 68332
rect 324314 68320 324320 68332
rect 271840 68292 324320 68320
rect 271840 68280 271846 68292
rect 324314 68280 324320 68292
rect 324372 68280 324378 68332
rect 335262 68280 335268 68332
rect 335320 68320 335326 68332
rect 416866 68320 416872 68332
rect 335320 68292 416872 68320
rect 335320 68280 335326 68292
rect 416866 68280 416872 68292
rect 416924 68280 416930 68332
rect 418062 68280 418068 68332
rect 418120 68320 418126 68332
rect 535454 68320 535460 68332
rect 418120 68292 535460 68320
rect 418120 68280 418126 68292
rect 535454 68280 535460 68292
rect 535512 68280 535518 68332
rect 270310 66852 270316 66904
rect 270368 66892 270374 66904
rect 321554 66892 321560 66904
rect 270368 66864 321560 66892
rect 270368 66852 270374 66864
rect 321554 66852 321560 66864
rect 321612 66852 321618 66904
rect 333882 66852 333888 66904
rect 333940 66892 333946 66904
rect 412634 66892 412640 66904
rect 333940 66864 412640 66892
rect 333940 66852 333946 66864
rect 412634 66852 412640 66864
rect 412692 66852 412698 66904
rect 430482 66852 430488 66904
rect 430540 66892 430546 66904
rect 553394 66892 553400 66904
rect 430540 66864 553400 66892
rect 430540 66852 430546 66864
rect 553394 66852 553400 66864
rect 553452 66852 553458 66904
rect 135438 66240 135444 66292
rect 135496 66280 135502 66292
rect 135714 66280 135720 66292
rect 135496 66252 135720 66280
rect 135496 66240 135502 66252
rect 135714 66240 135720 66252
rect 135772 66240 135778 66292
rect 267550 65492 267556 65544
rect 267608 65532 267614 65544
rect 317414 65532 317420 65544
rect 267608 65504 317420 65532
rect 267608 65492 267614 65504
rect 317414 65492 317420 65504
rect 317472 65492 317478 65544
rect 322750 65492 322756 65544
rect 322808 65532 322814 65544
rect 398834 65532 398840 65544
rect 322808 65504 398840 65532
rect 322808 65492 322814 65504
rect 398834 65492 398840 65504
rect 398892 65492 398898 65544
rect 426342 65492 426348 65544
rect 426400 65532 426406 65544
rect 546586 65532 546592 65544
rect 426400 65504 546592 65532
rect 426400 65492 426406 65504
rect 546586 65492 546592 65504
rect 546644 65492 546650 65544
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 129090 64852 129096 64864
rect 3384 64824 129096 64852
rect 3384 64812 3390 64824
rect 129090 64812 129096 64824
rect 129148 64812 129154 64864
rect 456058 64812 456064 64864
rect 456116 64852 456122 64864
rect 579798 64852 579804 64864
rect 456116 64824 579804 64852
rect 456116 64812 456122 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 264882 64132 264888 64184
rect 264940 64172 264946 64184
rect 313274 64172 313280 64184
rect 264940 64144 313280 64172
rect 264940 64132 264946 64144
rect 313274 64132 313280 64144
rect 313332 64132 313338 64184
rect 321462 64132 321468 64184
rect 321520 64172 321526 64184
rect 394694 64172 394700 64184
rect 321520 64144 394700 64172
rect 321520 64132 321526 64144
rect 394694 64132 394700 64144
rect 394752 64132 394758 64184
rect 313090 62772 313096 62824
rect 313148 62812 313154 62824
rect 383654 62812 383660 62824
rect 313148 62784 383660 62812
rect 313148 62772 313154 62784
rect 383654 62772 383660 62784
rect 383712 62772 383718 62824
rect 405642 62772 405648 62824
rect 405700 62812 405706 62824
rect 517514 62812 517520 62824
rect 405700 62784 517520 62812
rect 405700 62772 405706 62784
rect 517514 62772 517520 62784
rect 517572 62772 517578 62824
rect 262030 61344 262036 61396
rect 262088 61384 262094 61396
rect 310514 61384 310520 61396
rect 262088 61356 310520 61384
rect 262088 61344 262094 61356
rect 310514 61344 310520 61356
rect 310572 61344 310578 61396
rect 315298 61344 315304 61396
rect 315356 61384 315362 61396
rect 380894 61384 380900 61396
rect 315356 61356 380900 61384
rect 315356 61344 315362 61356
rect 380894 61344 380900 61356
rect 380952 61344 380958 61396
rect 413922 61344 413928 61396
rect 413980 61384 413986 61396
rect 528646 61384 528652 61396
rect 413980 61356 528652 61384
rect 413980 61344 413986 61356
rect 528646 61344 528652 61356
rect 528704 61344 528710 61396
rect 135438 60840 135444 60852
rect 135399 60812 135444 60840
rect 135438 60800 135444 60812
rect 135496 60800 135502 60852
rect 143718 60664 143724 60716
rect 143776 60704 143782 60716
rect 143902 60704 143908 60716
rect 143776 60676 143908 60704
rect 143776 60664 143782 60676
rect 143902 60664 143908 60676
rect 143960 60664 143966 60716
rect 308950 59984 308956 60036
rect 309008 60024 309014 60036
rect 376754 60024 376760 60036
rect 309008 59996 376760 60024
rect 309008 59984 309014 59996
rect 376754 59984 376760 59996
rect 376812 59984 376818 60036
rect 411162 59984 411168 60036
rect 411220 60024 411226 60036
rect 524414 60024 524420 60036
rect 411220 59996 524420 60024
rect 411220 59984 411226 59996
rect 524414 59984 524420 59996
rect 524472 59984 524478 60036
rect 257982 58624 257988 58676
rect 258040 58664 258046 58676
rect 303614 58664 303620 58676
rect 258040 58636 303620 58664
rect 258040 58624 258046 58636
rect 303614 58624 303620 58636
rect 303672 58624 303678 58676
rect 306282 58624 306288 58676
rect 306340 58664 306346 58676
rect 374086 58664 374092 58676
rect 306340 58636 374092 58664
rect 306340 58624 306346 58636
rect 374086 58624 374092 58636
rect 374144 58624 374150 58676
rect 393222 58624 393228 58676
rect 393280 58664 393286 58676
rect 499574 58664 499580 58676
rect 393280 58636 499580 58664
rect 393280 58624 393286 58636
rect 499574 58624 499580 58636
rect 499632 58624 499638 58676
rect 135438 57916 135444 57928
rect 135399 57888 135444 57916
rect 135438 57876 135444 57888
rect 135496 57876 135502 57928
rect 143721 57919 143779 57925
rect 143721 57885 143733 57919
rect 143767 57916 143779 57919
rect 143902 57916 143908 57928
rect 143767 57888 143908 57916
rect 143767 57885 143779 57888
rect 143721 57879 143779 57885
rect 143902 57876 143908 57888
rect 143960 57876 143966 57928
rect 255130 57196 255136 57248
rect 255188 57236 255194 57248
rect 299474 57236 299480 57248
rect 255188 57208 299480 57236
rect 255188 57196 255194 57208
rect 299474 57196 299480 57208
rect 299532 57196 299538 57248
rect 303430 57196 303436 57248
rect 303488 57236 303494 57248
rect 369854 57236 369860 57248
rect 303488 57208 369860 57236
rect 303488 57196 303494 57208
rect 369854 57196 369860 57208
rect 369912 57196 369918 57248
rect 383562 57196 383568 57248
rect 383620 57236 383626 57248
rect 485866 57236 485872 57248
rect 383620 57208 485872 57236
rect 383620 57196 383626 57208
rect 485866 57196 485872 57208
rect 485924 57196 485930 57248
rect 252462 55836 252468 55888
rect 252520 55876 252526 55888
rect 296806 55876 296812 55888
rect 252520 55848 296812 55876
rect 252520 55836 252526 55848
rect 296806 55836 296812 55848
rect 296864 55836 296870 55888
rect 300670 55836 300676 55888
rect 300728 55876 300734 55888
rect 365714 55876 365720 55888
rect 300728 55848 365720 55876
rect 300728 55836 300734 55848
rect 365714 55836 365720 55848
rect 365772 55836 365778 55888
rect 388990 55836 388996 55888
rect 389048 55876 389054 55888
rect 492674 55876 492680 55888
rect 389048 55848 492680 55876
rect 389048 55836 389054 55848
rect 492674 55836 492680 55848
rect 492732 55836 492738 55888
rect 249610 54476 249616 54528
rect 249668 54516 249674 54528
rect 292574 54516 292580 54528
rect 249668 54488 292580 54516
rect 249668 54476 249674 54488
rect 292574 54476 292580 54488
rect 292632 54476 292638 54528
rect 299382 54476 299388 54528
rect 299440 54516 299446 54528
rect 362954 54516 362960 54528
rect 299440 54488 362960 54516
rect 299440 54476 299446 54488
rect 362954 54476 362960 54488
rect 363012 54476 363018 54528
rect 378042 54476 378048 54528
rect 378100 54516 378106 54528
rect 477586 54516 477592 54528
rect 378100 54488 477592 54516
rect 378100 54476 378106 54488
rect 477586 54476 477592 54488
rect 477644 54476 477650 54528
rect 246850 53048 246856 53100
rect 246908 53088 246914 53100
rect 288434 53088 288440 53100
rect 246908 53060 288440 53088
rect 246908 53048 246914 53060
rect 288434 53048 288440 53060
rect 288492 53048 288498 53100
rect 293862 53048 293868 53100
rect 293920 53088 293926 53100
rect 356146 53088 356152 53100
rect 293920 53060 356152 53088
rect 293920 53048 293926 53060
rect 356146 53048 356152 53060
rect 356204 53048 356210 53100
rect 358630 53048 358636 53100
rect 358688 53088 358694 53100
rect 448514 53088 448520 53100
rect 358688 53060 448520 53088
rect 358688 53048 358694 53060
rect 448514 53048 448520 53060
rect 448572 53048 448578 53100
rect 291010 51756 291016 51808
rect 291068 51796 291074 51808
rect 351914 51796 351920 51808
rect 291068 51768 351920 51796
rect 291068 51756 291074 51768
rect 351914 51756 351920 51768
rect 351972 51756 351978 51808
rect 245470 51688 245476 51740
rect 245528 51728 245534 51740
rect 285674 51728 285680 51740
rect 245528 51700 285680 51728
rect 245528 51688 245534 51700
rect 285674 51688 285680 51700
rect 285732 51688 285738 51740
rect 350442 51688 350448 51740
rect 350500 51728 350506 51740
rect 437474 51728 437480 51740
rect 350500 51700 437480 51728
rect 350500 51688 350506 51700
rect 437474 51688 437480 51700
rect 437532 51688 437538 51740
rect 444282 51688 444288 51740
rect 444340 51728 444346 51740
rect 572714 51728 572720 51740
rect 444340 51700 572720 51728
rect 444340 51688 444346 51700
rect 572714 51688 572720 51700
rect 572772 51688 572778 51740
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 11698 51048 11704 51060
rect 3476 51020 11704 51048
rect 3476 51008 3482 51020
rect 11698 51008 11704 51020
rect 11756 51008 11762 51060
rect 288250 50396 288256 50448
rect 288308 50436 288314 50448
rect 347774 50436 347780 50448
rect 288308 50408 347780 50436
rect 288308 50396 288314 50408
rect 347774 50396 347780 50408
rect 347832 50396 347838 50448
rect 242802 50328 242808 50380
rect 242860 50368 242866 50380
rect 281534 50368 281540 50380
rect 242860 50340 281540 50368
rect 242860 50328 242866 50340
rect 281534 50328 281540 50340
rect 281592 50328 281598 50380
rect 346302 50328 346308 50380
rect 346360 50368 346366 50380
rect 431954 50368 431960 50380
rect 346360 50340 431960 50368
rect 346360 50328 346366 50340
rect 431954 50328 431960 50340
rect 432012 50328 432018 50380
rect 434622 50328 434628 50380
rect 434680 50368 434686 50380
rect 558914 50368 558920 50380
rect 434680 50340 558920 50368
rect 434680 50328 434686 50340
rect 558914 50328 558920 50340
rect 558972 50328 558978 50380
rect 239950 48968 239956 49020
rect 240008 49008 240014 49020
rect 278774 49008 278780 49020
rect 240008 48980 278780 49008
rect 240008 48968 240014 48980
rect 278774 48968 278780 48980
rect 278832 48968 278838 49020
rect 284202 48968 284208 49020
rect 284260 49008 284266 49020
rect 340874 49008 340880 49020
rect 284260 48980 340880 49008
rect 284260 48968 284266 48980
rect 340874 48968 340880 48980
rect 340932 48968 340938 49020
rect 409782 48968 409788 49020
rect 409840 49008 409846 49020
rect 523034 49008 523040 49020
rect 409840 48980 523040 49008
rect 409840 48968 409846 48980
rect 523034 48968 523040 48980
rect 523092 48968 523098 49020
rect 143718 48328 143724 48340
rect 143679 48300 143724 48328
rect 143718 48288 143724 48300
rect 143776 48288 143782 48340
rect 331122 47608 331128 47660
rect 331180 47648 331186 47660
rect 408586 47648 408592 47660
rect 331180 47620 408592 47648
rect 331180 47608 331186 47620
rect 408586 47608 408592 47620
rect 408644 47608 408650 47660
rect 237190 47540 237196 47592
rect 237248 47580 237254 47592
rect 274634 47580 274640 47592
rect 237248 47552 274640 47580
rect 237248 47540 237254 47552
rect 274634 47540 274640 47552
rect 274692 47540 274698 47592
rect 275922 47540 275928 47592
rect 275980 47580 275986 47592
rect 331306 47580 331312 47592
rect 275980 47552 331312 47580
rect 275980 47540 275986 47552
rect 331306 47540 331312 47552
rect 331364 47540 331370 47592
rect 407022 47540 407028 47592
rect 407080 47580 407086 47592
rect 520366 47580 520372 47592
rect 407080 47552 520372 47580
rect 407080 47540 407086 47552
rect 520366 47540 520372 47552
rect 520424 47540 520430 47592
rect 235902 46180 235908 46232
rect 235960 46220 235966 46232
rect 270494 46220 270500 46232
rect 235960 46192 270500 46220
rect 235960 46180 235966 46192
rect 270494 46180 270500 46192
rect 270552 46180 270558 46232
rect 278590 46180 278596 46232
rect 278648 46220 278654 46232
rect 333974 46220 333980 46232
rect 278648 46192 333980 46220
rect 278648 46180 278654 46192
rect 333974 46180 333980 46192
rect 334032 46180 334038 46232
rect 375282 46180 375288 46232
rect 375340 46220 375346 46232
rect 471974 46220 471980 46232
rect 375340 46192 471980 46220
rect 375340 46180 375346 46192
rect 471974 46180 471980 46192
rect 472032 46180 472038 46232
rect 274542 44888 274548 44940
rect 274600 44928 274606 44940
rect 327074 44928 327080 44940
rect 274600 44900 327080 44928
rect 274600 44888 274606 44900
rect 327074 44888 327080 44900
rect 327132 44888 327138 44940
rect 233050 44820 233056 44872
rect 233108 44860 233114 44872
rect 267734 44860 267740 44872
rect 233108 44832 267740 44860
rect 233108 44820 233114 44832
rect 267734 44820 267740 44832
rect 267792 44820 267798 44872
rect 325602 44820 325608 44872
rect 325660 44860 325666 44872
rect 401594 44860 401600 44872
rect 325660 44832 401600 44860
rect 325660 44820 325666 44832
rect 401594 44820 401600 44832
rect 401652 44820 401658 44872
rect 424962 44820 424968 44872
rect 425020 44860 425026 44872
rect 545114 44860 545120 44872
rect 425020 44832 545120 44860
rect 425020 44820 425026 44832
rect 545114 44820 545120 44832
rect 545172 44820 545178 44872
rect 269022 43392 269028 43444
rect 269080 43432 269086 43444
rect 320174 43432 320180 43444
rect 269080 43404 320180 43432
rect 269080 43392 269086 43404
rect 320174 43392 320180 43404
rect 320232 43392 320238 43444
rect 360102 43392 360108 43444
rect 360160 43432 360166 43444
rect 451366 43432 451372 43444
rect 360160 43404 451372 43432
rect 360160 43392 360166 43404
rect 451366 43392 451372 43404
rect 451424 43392 451430 43444
rect 266170 42100 266176 42152
rect 266228 42140 266234 42152
rect 316034 42140 316040 42152
rect 266228 42112 316040 42140
rect 266228 42100 266234 42112
rect 316034 42100 316040 42112
rect 316092 42100 316098 42152
rect 230382 42032 230388 42084
rect 230440 42072 230446 42084
rect 263594 42072 263600 42084
rect 230440 42044 263600 42072
rect 230440 42032 230446 42044
rect 263594 42032 263600 42044
rect 263652 42032 263658 42084
rect 315942 42032 315948 42084
rect 316000 42072 316006 42084
rect 387794 42072 387800 42084
rect 316000 42044 387800 42072
rect 316000 42032 316006 42044
rect 387794 42032 387800 42044
rect 387852 42032 387858 42084
rect 402882 42032 402888 42084
rect 402940 42072 402946 42084
rect 512086 42072 512092 42084
rect 402940 42044 512092 42072
rect 402940 42032 402946 42044
rect 512086 42032 512092 42044
rect 512144 42032 512150 42084
rect 478138 41352 478144 41404
rect 478196 41392 478202 41404
rect 580166 41392 580172 41404
rect 478196 41364 580172 41392
rect 478196 41352 478202 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 227622 40672 227628 40724
rect 227680 40712 227686 40724
rect 260834 40712 260840 40724
rect 227680 40684 260840 40712
rect 227680 40672 227686 40684
rect 260834 40672 260840 40684
rect 260892 40672 260898 40724
rect 263410 40672 263416 40724
rect 263468 40712 263474 40724
rect 313366 40712 313372 40724
rect 263468 40684 313372 40712
rect 263468 40672 263474 40684
rect 313366 40672 313372 40684
rect 313424 40672 313430 40724
rect 354582 40672 354588 40724
rect 354640 40712 354646 40724
rect 443086 40712 443092 40724
rect 354640 40684 443092 40712
rect 354640 40672 354646 40684
rect 443086 40672 443092 40684
rect 443144 40672 443150 40724
rect 262122 39380 262128 39432
rect 262180 39420 262186 39432
rect 309134 39420 309140 39432
rect 262180 39392 309140 39420
rect 262180 39380 262186 39392
rect 309134 39380 309140 39392
rect 309192 39380 309198 39432
rect 224770 39312 224776 39364
rect 224828 39352 224834 39364
rect 256694 39352 256700 39364
rect 224828 39324 256700 39352
rect 224828 39312 224834 39324
rect 256694 39312 256700 39324
rect 256752 39312 256758 39364
rect 296530 39312 296536 39364
rect 296588 39352 296594 39364
rect 360194 39352 360200 39364
rect 296588 39324 360200 39352
rect 296588 39312 296594 39324
rect 360194 39312 360200 39324
rect 360252 39312 360258 39364
rect 362862 39312 362868 39364
rect 362920 39352 362926 39364
rect 454034 39352 454040 39364
rect 362920 39324 454040 39352
rect 362920 39312 362926 39324
rect 454034 39312 454040 39324
rect 454092 39312 454098 39364
rect 143718 38632 143724 38684
rect 143776 38672 143782 38684
rect 143902 38672 143908 38684
rect 143776 38644 143908 38672
rect 143776 38632 143782 38644
rect 143902 38632 143908 38644
rect 143960 38632 143966 38684
rect 256602 37884 256608 37936
rect 256660 37924 256666 37936
rect 302234 37924 302240 37936
rect 256660 37896 302240 37924
rect 256660 37884 256666 37896
rect 302234 37884 302240 37896
rect 302292 37884 302298 37936
rect 342162 37884 342168 37936
rect 342220 37924 342226 37936
rect 425146 37924 425152 37936
rect 342220 37896 425152 37924
rect 342220 37884 342226 37896
rect 425146 37884 425152 37896
rect 425204 37884 425210 37936
rect 431862 37884 431868 37936
rect 431920 37924 431926 37936
rect 554866 37924 554872 37936
rect 431920 37896 554872 37924
rect 431920 37884 431926 37896
rect 554866 37884 554872 37896
rect 554924 37884 554930 37936
rect 296622 36592 296628 36644
rect 296680 36632 296686 36644
rect 358814 36632 358820 36644
rect 296680 36604 358820 36632
rect 296680 36592 296686 36604
rect 358814 36592 358820 36604
rect 358872 36592 358878 36644
rect 220630 36524 220636 36576
rect 220688 36564 220694 36576
rect 249794 36564 249800 36576
rect 220688 36536 249800 36564
rect 220688 36524 220694 36536
rect 249794 36524 249800 36536
rect 249852 36524 249858 36576
rect 250990 36524 250996 36576
rect 251048 36564 251054 36576
rect 295334 36564 295340 36576
rect 251048 36536 295340 36564
rect 251048 36524 251054 36536
rect 295334 36524 295340 36536
rect 295392 36524 295398 36576
rect 357342 36524 357348 36576
rect 357400 36564 357406 36576
rect 447134 36564 447140 36576
rect 357400 36536 447140 36564
rect 357400 36524 357406 36536
rect 447134 36524 447140 36536
rect 447192 36524 447198 36576
rect 449802 36524 449808 36576
rect 449860 36564 449866 36576
rect 578970 36564 578976 36576
rect 449860 36536 578976 36564
rect 449860 36524 449866 36536
rect 578970 36524 578976 36536
rect 579028 36524 579034 36576
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 7558 35884 7564 35896
rect 3476 35856 7564 35884
rect 3476 35844 3482 35856
rect 7558 35844 7564 35856
rect 7616 35844 7622 35896
rect 249702 35164 249708 35216
rect 249760 35204 249766 35216
rect 291194 35204 291200 35216
rect 249760 35176 291200 35204
rect 249760 35164 249766 35176
rect 291194 35164 291200 35176
rect 291252 35164 291258 35216
rect 317322 35164 317328 35216
rect 317380 35204 317386 35216
rect 390646 35204 390652 35216
rect 317380 35176 390652 35204
rect 317380 35164 317386 35176
rect 390646 35164 390652 35176
rect 390704 35164 390710 35216
rect 394602 35164 394608 35216
rect 394660 35204 394666 35216
rect 502426 35204 502432 35216
rect 394660 35176 502432 35204
rect 394660 35164 394666 35176
rect 502426 35164 502432 35176
rect 502484 35164 502490 35216
rect 246942 33804 246948 33856
rect 247000 33844 247006 33856
rect 287054 33844 287060 33856
rect 247000 33816 287060 33844
rect 247000 33804 247006 33816
rect 287054 33804 287060 33816
rect 287112 33804 287118 33856
rect 217962 33736 217968 33788
rect 218020 33776 218026 33788
rect 245654 33776 245660 33788
rect 218020 33748 245660 33776
rect 218020 33736 218026 33748
rect 245654 33736 245660 33748
rect 245712 33736 245718 33788
rect 286962 33736 286968 33788
rect 287020 33776 287026 33788
rect 345014 33776 345020 33788
rect 287020 33748 345020 33776
rect 287020 33736 287026 33748
rect 345014 33736 345020 33748
rect 345072 33736 345078 33788
rect 351822 33736 351828 33788
rect 351880 33776 351886 33788
rect 440234 33776 440240 33788
rect 351880 33748 440240 33776
rect 351880 33736 351886 33748
rect 440234 33736 440240 33748
rect 440292 33736 440298 33788
rect 447042 33736 447048 33788
rect 447100 33776 447106 33788
rect 576854 33776 576860 33788
rect 447100 33748 576860 33776
rect 447100 33736 447106 33748
rect 576854 33736 576860 33748
rect 576912 33736 576918 33788
rect 215110 32376 215116 32428
rect 215168 32416 215174 32428
rect 242894 32416 242900 32428
rect 215168 32388 242900 32416
rect 215168 32376 215174 32388
rect 242894 32376 242900 32388
rect 242952 32376 242958 32428
rect 244090 32376 244096 32428
rect 244148 32416 244154 32428
rect 284294 32416 284300 32428
rect 244148 32388 284300 32416
rect 244148 32376 244154 32388
rect 284294 32376 284300 32388
rect 284352 32376 284358 32428
rect 314562 32376 314568 32428
rect 314620 32416 314626 32428
rect 386414 32416 386420 32428
rect 314620 32388 386420 32416
rect 314620 32376 314626 32388
rect 386414 32376 386420 32388
rect 386472 32376 386478 32428
rect 387702 32376 387708 32428
rect 387760 32416 387766 32428
rect 491294 32416 491300 32428
rect 387760 32388 491300 32416
rect 387760 32376 387766 32388
rect 491294 32376 491300 32388
rect 491352 32376 491358 32428
rect 241422 31016 241428 31068
rect 241480 31056 241486 31068
rect 280154 31056 280160 31068
rect 241480 31028 280160 31056
rect 241480 31016 241486 31028
rect 280154 31016 280160 31028
rect 280212 31016 280218 31068
rect 281442 31016 281448 31068
rect 281500 31056 281506 31068
rect 338114 31056 338120 31068
rect 281500 31028 338120 31056
rect 281500 31016 281506 31028
rect 338114 31016 338120 31028
rect 338172 31016 338178 31068
rect 348418 31016 348424 31068
rect 348476 31056 348482 31068
rect 433426 31056 433432 31068
rect 348476 31028 433432 31056
rect 348476 31016 348482 31028
rect 433426 31016 433432 31028
rect 433484 31016 433490 31068
rect 441522 31016 441528 31068
rect 441580 31056 441586 31068
rect 568574 31056 568580 31068
rect 441580 31028 568580 31056
rect 441580 31016 441586 31028
rect 568574 31016 568580 31028
rect 568632 31016 568638 31068
rect 453298 30268 453304 30320
rect 453356 30308 453362 30320
rect 580166 30308 580172 30320
rect 453356 30280 580172 30308
rect 453356 30268 453362 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 240042 29588 240048 29640
rect 240100 29628 240106 29640
rect 277394 29628 277400 29640
rect 240100 29600 277400 29628
rect 240100 29588 240106 29600
rect 277394 29588 277400 29600
rect 277452 29588 277458 29640
rect 304902 29588 304908 29640
rect 304960 29628 304966 29640
rect 372614 29628 372620 29640
rect 304960 29600 372620 29628
rect 304960 29588 304966 29600
rect 372614 29588 372620 29600
rect 372672 29588 372678 29640
rect 259362 28296 259368 28348
rect 259420 28336 259426 28348
rect 306374 28336 306380 28348
rect 259420 28308 306380 28336
rect 259420 28296 259426 28308
rect 306374 28296 306380 28308
rect 306432 28296 306438 28348
rect 234522 28228 234528 28280
rect 234580 28268 234586 28280
rect 270586 28268 270592 28280
rect 234580 28240 270592 28268
rect 234580 28228 234586 28240
rect 270586 28228 270592 28240
rect 270644 28228 270650 28280
rect 303522 28228 303528 28280
rect 303580 28268 303586 28280
rect 368474 28268 368480 28280
rect 303580 28240 368480 28268
rect 303580 28228 303586 28240
rect 368474 28228 368480 28240
rect 368532 28228 368538 28280
rect 369762 28228 369768 28280
rect 369820 28268 369826 28280
rect 465074 28268 465080 28280
rect 369820 28240 465080 28268
rect 369820 28228 369826 28240
rect 465074 28228 465080 28240
rect 465132 28228 465138 28280
rect 135438 27548 135444 27600
rect 135496 27588 135502 27600
rect 135533 27591 135591 27597
rect 135533 27588 135545 27591
rect 135496 27560 135545 27588
rect 135496 27548 135502 27560
rect 135533 27557 135545 27560
rect 135579 27557 135591 27591
rect 135533 27551 135591 27557
rect 143718 27548 143724 27600
rect 143776 27588 143782 27600
rect 143994 27588 144000 27600
rect 143776 27560 144000 27588
rect 143776 27548 143782 27560
rect 143994 27548 144000 27560
rect 144052 27548 144058 27600
rect 224862 26868 224868 26920
rect 224920 26908 224926 26920
rect 255314 26908 255320 26920
rect 224920 26880 255320 26908
rect 224920 26868 224926 26880
rect 255314 26868 255320 26880
rect 255372 26868 255378 26920
rect 257338 26868 257344 26920
rect 257396 26908 257402 26920
rect 298094 26908 298100 26920
rect 257396 26880 298100 26908
rect 257396 26868 257402 26880
rect 298094 26868 298100 26880
rect 298152 26868 298158 26920
rect 300762 26868 300768 26920
rect 300820 26908 300826 26920
rect 365806 26908 365812 26920
rect 300820 26880 365812 26908
rect 300820 26868 300826 26880
rect 365806 26868 365812 26880
rect 365864 26868 365870 26920
rect 372522 26868 372528 26920
rect 372580 26908 372586 26920
rect 467926 26908 467932 26920
rect 372580 26880 467932 26908
rect 372580 26868 372586 26880
rect 467926 26868 467932 26880
rect 467984 26868 467990 26920
rect 212350 25576 212356 25628
rect 212408 25616 212414 25628
rect 237374 25616 237380 25628
rect 212408 25588 237380 25616
rect 212408 25576 212414 25588
rect 237374 25576 237380 25588
rect 237432 25576 237438 25628
rect 237282 25508 237288 25560
rect 237340 25548 237346 25560
rect 273254 25548 273260 25560
rect 237340 25520 273260 25548
rect 237340 25508 237346 25520
rect 273254 25508 273260 25520
rect 273312 25508 273318 25560
rect 298002 25508 298008 25560
rect 298060 25548 298066 25560
rect 361574 25548 361580 25560
rect 298060 25520 361580 25548
rect 298060 25508 298066 25520
rect 361574 25508 361580 25520
rect 361632 25508 361638 25560
rect 429102 25508 429108 25560
rect 429160 25548 429166 25560
rect 550634 25548 550640 25560
rect 429160 25520 550640 25548
rect 429160 25508 429166 25520
rect 550634 25508 550640 25520
rect 550692 25508 550698 25560
rect 339402 24148 339408 24200
rect 339460 24188 339466 24200
rect 422294 24188 422300 24200
rect 339460 24160 422300 24188
rect 339460 24148 339466 24160
rect 422294 24148 422300 24160
rect 422352 24148 422358 24200
rect 206830 24080 206836 24132
rect 206888 24120 206894 24132
rect 230474 24120 230480 24132
rect 206888 24092 230480 24120
rect 206888 24080 206894 24092
rect 230474 24080 230480 24092
rect 230532 24080 230538 24132
rect 231670 24080 231676 24132
rect 231728 24120 231734 24132
rect 266354 24120 266360 24132
rect 231728 24092 266360 24120
rect 231728 24080 231734 24092
rect 266354 24080 266360 24092
rect 266412 24080 266418 24132
rect 282822 24080 282828 24132
rect 282880 24120 282886 24132
rect 339586 24120 339592 24132
rect 282880 24092 339592 24120
rect 282880 24080 282886 24092
rect 339586 24080 339592 24092
rect 339644 24080 339650 24132
rect 422202 24080 422208 24132
rect 422260 24120 422266 24132
rect 540974 24120 540980 24132
rect 422260 24092 540980 24120
rect 422260 24080 422266 24092
rect 540974 24080 540980 24092
rect 541032 24080 541038 24132
rect 204070 22720 204076 22772
rect 204128 22760 204134 22772
rect 227806 22760 227812 22772
rect 204128 22732 227812 22760
rect 204128 22720 204134 22732
rect 227806 22720 227812 22732
rect 227864 22720 227870 22772
rect 228910 22720 228916 22772
rect 228968 22760 228974 22772
rect 262214 22760 262220 22772
rect 228968 22732 262220 22760
rect 228968 22720 228974 22732
rect 262214 22720 262220 22732
rect 262272 22720 262278 22772
rect 280062 22720 280068 22772
rect 280120 22760 280126 22772
rect 336734 22760 336740 22772
rect 280120 22732 336740 22760
rect 280120 22720 280126 22732
rect 336734 22720 336740 22732
rect 336792 22720 336798 22772
rect 338022 22720 338028 22772
rect 338080 22760 338086 22772
rect 418154 22760 418160 22772
rect 338080 22732 418160 22760
rect 338080 22720 338086 22732
rect 418154 22720 418160 22732
rect 418212 22720 418218 22772
rect 419442 22720 419448 22772
rect 419500 22760 419506 22772
rect 536926 22760 536932 22772
rect 419500 22732 536932 22760
rect 419500 22720 419506 22732
rect 536926 22720 536932 22732
rect 536984 22720 536990 22772
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 128998 22080 129004 22092
rect 3200 22052 129004 22080
rect 3200 22040 3206 22052
rect 128998 22040 129004 22052
rect 129056 22040 129062 22092
rect 204898 21428 204904 21480
rect 204956 21468 204962 21480
rect 223574 21468 223580 21480
rect 204956 21440 223580 21468
rect 204956 21428 204962 21440
rect 223574 21428 223580 21440
rect 223632 21428 223638 21480
rect 278682 21428 278688 21480
rect 278740 21468 278746 21480
rect 332594 21468 332600 21480
rect 278740 21440 332600 21468
rect 278740 21428 278746 21440
rect 332594 21428 332600 21440
rect 332652 21428 332658 21480
rect 222838 21360 222844 21412
rect 222896 21400 222902 21412
rect 252646 21400 252652 21412
rect 222896 21372 252652 21400
rect 222896 21360 222902 21372
rect 252646 21360 252652 21372
rect 252704 21360 252710 21412
rect 332502 21360 332508 21412
rect 332560 21400 332566 21412
rect 411254 21400 411260 21412
rect 332560 21372 411260 21400
rect 332560 21360 332566 21372
rect 411254 21360 411260 21372
rect 411312 21360 411318 21412
rect 412542 21360 412548 21412
rect 412600 21400 412606 21412
rect 527174 21400 527180 21412
rect 412600 21372 527180 21400
rect 412600 21360 412606 21372
rect 527174 21360 527180 21372
rect 527232 21360 527238 21412
rect 200758 20000 200764 20052
rect 200816 20040 200822 20052
rect 219434 20040 219440 20052
rect 200816 20012 219440 20040
rect 200816 20000 200822 20012
rect 219434 20000 219440 20012
rect 219492 20000 219498 20052
rect 219250 19932 219256 19984
rect 219308 19972 219314 19984
rect 248414 19972 248420 19984
rect 219308 19944 248420 19972
rect 219308 19932 219314 19944
rect 248414 19932 248420 19944
rect 248472 19932 248478 19984
rect 266262 19932 266268 19984
rect 266320 19972 266326 19984
rect 314654 19972 314660 19984
rect 266320 19944 314660 19972
rect 266320 19932 266326 19944
rect 314654 19932 314660 19944
rect 314712 19932 314718 19984
rect 326982 19932 326988 19984
rect 327040 19972 327046 19984
rect 404354 19972 404360 19984
rect 327040 19944 404360 19972
rect 327040 19932 327046 19944
rect 404354 19932 404360 19944
rect 404412 19932 404418 19984
rect 416682 19932 416688 19984
rect 416740 19972 416746 19984
rect 532694 19972 532700 19984
rect 416740 19944 532700 19972
rect 416740 19932 416746 19944
rect 532694 19932 532700 19944
rect 532752 19932 532758 19984
rect 301498 19252 301504 19304
rect 301556 19292 301562 19304
rect 305086 19292 305092 19304
rect 301556 19264 305092 19292
rect 301556 19252 301562 19264
rect 305086 19252 305092 19264
rect 305144 19252 305150 19304
rect 197262 18640 197268 18692
rect 197320 18680 197326 18692
rect 216674 18680 216680 18692
rect 197320 18652 216680 18680
rect 197320 18640 197326 18652
rect 216674 18640 216680 18652
rect 216732 18640 216738 18692
rect 216490 18572 216496 18624
rect 216548 18612 216554 18624
rect 244274 18612 244280 18624
rect 216548 18584 244280 18612
rect 216548 18572 216554 18584
rect 244274 18572 244280 18584
rect 244332 18572 244338 18624
rect 255222 18572 255228 18624
rect 255280 18612 255286 18624
rect 300854 18612 300860 18624
rect 255280 18584 300860 18612
rect 255280 18572 255286 18584
rect 300854 18572 300860 18584
rect 300912 18572 300918 18624
rect 310422 18572 310428 18624
rect 310480 18612 310486 18624
rect 379514 18612 379520 18624
rect 310480 18584 379520 18612
rect 310480 18572 310486 18584
rect 379514 18572 379520 18584
rect 379572 18572 379578 18624
rect 390462 18572 390468 18624
rect 390520 18612 390526 18624
rect 494146 18612 494152 18624
rect 390520 18584 494152 18612
rect 390520 18572 390526 18584
rect 494146 18572 494152 18584
rect 494204 18572 494210 18624
rect 483658 17892 483664 17944
rect 483716 17932 483722 17944
rect 579798 17932 579804 17944
rect 483716 17904 579804 17932
rect 483716 17892 483722 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 251082 17280 251088 17332
rect 251140 17320 251146 17332
rect 293954 17320 293960 17332
rect 251140 17292 293960 17320
rect 251140 17280 251146 17292
rect 293954 17280 293960 17292
rect 294012 17280 294018 17332
rect 194410 17212 194416 17264
rect 194468 17252 194474 17264
rect 212534 17252 212540 17264
rect 194468 17224 212540 17252
rect 194468 17212 194474 17224
rect 212534 17212 212540 17224
rect 212592 17212 212598 17264
rect 215202 17212 215208 17264
rect 215260 17252 215266 17264
rect 241514 17252 241520 17264
rect 215260 17224 241520 17252
rect 215260 17212 215266 17224
rect 241514 17212 241520 17224
rect 241572 17212 241578 17264
rect 292482 17212 292488 17264
rect 292540 17252 292546 17264
rect 354674 17252 354680 17264
rect 292540 17224 354680 17252
rect 292540 17212 292546 17224
rect 354674 17212 354680 17224
rect 354732 17212 354738 17264
rect 384298 17212 384304 17264
rect 384356 17252 384362 17264
rect 436094 17252 436100 17264
rect 384356 17224 436100 17252
rect 384356 17212 384362 17224
rect 436094 17212 436100 17224
rect 436152 17212 436158 17264
rect 209682 15920 209688 15972
rect 209740 15960 209746 15972
rect 234614 15960 234620 15972
rect 209740 15932 234620 15960
rect 209740 15920 209746 15932
rect 234614 15920 234620 15932
rect 234672 15920 234678 15972
rect 191650 15852 191656 15904
rect 191708 15892 191714 15904
rect 209866 15892 209872 15904
rect 191708 15864 209872 15892
rect 191708 15852 191714 15864
rect 209866 15852 209872 15864
rect 209924 15852 209930 15904
rect 233142 15852 233148 15904
rect 233200 15892 233206 15904
rect 269114 15892 269120 15904
rect 233200 15864 269120 15892
rect 233200 15852 233206 15864
rect 269114 15852 269120 15864
rect 269172 15852 269178 15904
rect 270402 15852 270408 15904
rect 270460 15892 270466 15904
rect 321646 15892 321652 15904
rect 270460 15864 321652 15892
rect 270460 15852 270466 15864
rect 321646 15852 321652 15864
rect 321704 15852 321710 15904
rect 322842 15852 322848 15904
rect 322900 15892 322906 15904
rect 397454 15892 397460 15904
rect 322900 15864 397460 15892
rect 322900 15852 322906 15864
rect 397454 15852 397460 15864
rect 397512 15852 397518 15904
rect 400122 15852 400128 15904
rect 400180 15892 400186 15904
rect 509234 15892 509240 15904
rect 400180 15864 509240 15892
rect 400180 15852 400186 15864
rect 509234 15852 509240 15864
rect 509292 15852 509298 15904
rect 288342 14492 288348 14544
rect 288400 14532 288406 14544
rect 347866 14532 347872 14544
rect 288400 14504 347872 14532
rect 288400 14492 288406 14504
rect 347866 14492 347872 14504
rect 347924 14492 347930 14544
rect 190270 14424 190276 14476
rect 190328 14464 190334 14476
rect 205634 14464 205640 14476
rect 190328 14436 205640 14464
rect 190328 14424 190334 14436
rect 205634 14424 205640 14436
rect 205692 14424 205698 14476
rect 216582 14424 216588 14476
rect 216640 14464 216646 14476
rect 244366 14464 244372 14476
rect 216640 14436 244372 14464
rect 216640 14424 216646 14436
rect 244366 14424 244372 14436
rect 244424 14424 244430 14476
rect 245562 14424 245568 14476
rect 245620 14464 245626 14476
rect 287146 14464 287152 14476
rect 245620 14436 287152 14464
rect 245620 14424 245626 14436
rect 287146 14424 287152 14436
rect 287204 14424 287210 14476
rect 344922 14424 344928 14476
rect 344980 14464 344986 14476
rect 429194 14464 429200 14476
rect 344980 14436 429200 14464
rect 344980 14424 344986 14436
rect 429194 14424 429200 14436
rect 429252 14424 429258 14476
rect 436002 14424 436008 14476
rect 436060 14464 436066 14476
rect 561674 14464 561680 14476
rect 436060 14436 561680 14464
rect 436060 14424 436066 14436
rect 561674 14424 561680 14436
rect 561732 14424 561738 14476
rect 187510 13064 187516 13116
rect 187568 13104 187574 13116
rect 201494 13104 201500 13116
rect 187568 13076 201500 13104
rect 187568 13064 187574 13076
rect 201494 13064 201500 13076
rect 201552 13064 201558 13116
rect 208210 13064 208216 13116
rect 208268 13104 208274 13116
rect 233234 13104 233240 13116
rect 208268 13076 233240 13104
rect 208268 13064 208274 13076
rect 233234 13064 233240 13076
rect 233292 13064 233298 13116
rect 244182 13064 244188 13116
rect 244240 13104 244246 13116
rect 282914 13104 282920 13116
rect 244240 13076 282920 13104
rect 244240 13064 244246 13076
rect 282914 13064 282920 13076
rect 282972 13064 282978 13116
rect 285582 13064 285588 13116
rect 285640 13104 285646 13116
rect 343634 13104 343640 13116
rect 285640 13076 343640 13104
rect 285640 13064 285646 13076
rect 343634 13064 343640 13076
rect 343692 13064 343698 13116
rect 404262 13064 404268 13116
rect 404320 13104 404326 13116
rect 514754 13104 514760 13116
rect 404320 13076 514760 13104
rect 404320 13064 404326 13076
rect 514754 13064 514760 13076
rect 514812 13064 514818 13116
rect 135530 11744 135536 11756
rect 135491 11716 135536 11744
rect 135530 11704 135536 11716
rect 135588 11704 135594 11756
rect 184842 11704 184848 11756
rect 184900 11744 184906 11756
rect 198734 11744 198740 11756
rect 184900 11716 198740 11744
rect 184900 11704 184906 11716
rect 198734 11704 198740 11716
rect 198792 11704 198798 11756
rect 204162 11704 204168 11756
rect 204220 11744 204226 11756
rect 226334 11744 226340 11756
rect 204220 11716 226340 11744
rect 204220 11704 204226 11716
rect 226334 11704 226340 11716
rect 226392 11704 226398 11756
rect 229002 11704 229008 11756
rect 229060 11744 229066 11756
rect 262306 11744 262312 11756
rect 229060 11716 262312 11744
rect 229060 11704 229066 11716
rect 262306 11704 262312 11716
rect 262364 11704 262370 11756
rect 263502 11704 263508 11756
rect 263560 11744 263566 11756
rect 311894 11744 311900 11756
rect 263560 11716 311900 11744
rect 263560 11704 263566 11716
rect 311894 11704 311900 11716
rect 311952 11704 311958 11756
rect 313182 11704 313188 11756
rect 313240 11744 313246 11756
rect 382366 11744 382372 11756
rect 313240 11716 382372 11744
rect 313240 11704 313246 11716
rect 382366 11704 382372 11716
rect 382424 11704 382430 11756
rect 391842 11704 391848 11756
rect 391900 11744 391906 11756
rect 496814 11744 496820 11756
rect 391900 11716 496820 11744
rect 391900 11704 391906 11716
rect 496814 11704 496820 11716
rect 496872 11704 496878 11756
rect 188982 10276 188988 10328
rect 189040 10316 189046 10328
rect 204254 10316 204260 10328
rect 189040 10288 204260 10316
rect 189040 10276 189046 10288
rect 204254 10276 204260 10288
rect 204312 10276 204318 10328
rect 206922 10276 206928 10328
rect 206980 10316 206986 10328
rect 229094 10316 229100 10328
rect 206980 10288 229100 10316
rect 206980 10276 206986 10288
rect 229094 10276 229100 10288
rect 229152 10276 229158 10328
rect 231762 10276 231768 10328
rect 231820 10316 231826 10328
rect 264974 10316 264980 10328
rect 231820 10288 264980 10316
rect 231820 10276 231826 10288
rect 264974 10276 264980 10288
rect 265032 10276 265038 10328
rect 267642 10276 267648 10328
rect 267700 10316 267706 10328
rect 318794 10316 318800 10328
rect 267700 10288 318800 10316
rect 267700 10276 267706 10288
rect 318794 10276 318800 10288
rect 318852 10276 318858 10328
rect 320082 10276 320088 10328
rect 320140 10316 320146 10328
rect 393314 10316 393320 10328
rect 320140 10288 393320 10316
rect 320140 10276 320146 10288
rect 393314 10276 393320 10288
rect 393372 10276 393378 10328
rect 423582 10276 423588 10328
rect 423640 10316 423646 10328
rect 543734 10316 543740 10328
rect 423640 10288 543740 10316
rect 423640 10276 423646 10288
rect 543734 10276 543740 10288
rect 543792 10276 543798 10328
rect 238662 8984 238668 9036
rect 238720 9024 238726 9036
rect 276474 9024 276480 9036
rect 238720 8996 276480 9024
rect 238720 8984 238726 8996
rect 276474 8984 276480 8996
rect 276532 8984 276538 9036
rect 191742 8916 191748 8968
rect 191800 8956 191806 8968
rect 208670 8956 208676 8968
rect 191800 8928 208676 8956
rect 191800 8916 191806 8928
rect 208670 8916 208676 8928
rect 208728 8916 208734 8968
rect 210970 8916 210976 8968
rect 211028 8956 211034 8968
rect 237190 8956 237196 8968
rect 211028 8928 237196 8956
rect 211028 8916 211034 8928
rect 237190 8916 237196 8928
rect 237248 8916 237254 8968
rect 273162 8916 273168 8968
rect 273220 8956 273226 8968
rect 326430 8956 326436 8968
rect 273220 8928 326436 8956
rect 273220 8916 273226 8928
rect 326430 8916 326436 8928
rect 326488 8916 326494 8968
rect 327718 8916 327724 8968
rect 327776 8956 327782 8968
rect 401318 8956 401324 8968
rect 327776 8928 401324 8956
rect 327776 8916 327782 8928
rect 401318 8916 401324 8928
rect 401376 8916 401382 8968
rect 451918 8916 451924 8968
rect 451976 8956 451982 8968
rect 526254 8956 526260 8968
rect 451976 8928 526260 8956
rect 451976 8916 451982 8928
rect 526254 8916 526260 8928
rect 526312 8916 526318 8968
rect 2774 8100 2780 8152
rect 2832 8140 2838 8152
rect 6178 8140 6184 8152
rect 2832 8112 6184 8140
rect 2832 8100 2838 8112
rect 6178 8100 6184 8112
rect 6236 8100 6242 8152
rect 183370 7556 183376 7608
rect 183428 7596 183434 7608
rect 197998 7596 198004 7608
rect 183428 7568 198004 7596
rect 183428 7556 183434 7568
rect 197998 7556 198004 7568
rect 198056 7556 198062 7608
rect 198550 7556 198556 7608
rect 198608 7596 198614 7608
rect 198608 7568 209820 7596
rect 198608 7556 198614 7568
rect 209792 7528 209820 7568
rect 219342 7556 219348 7608
rect 219400 7596 219406 7608
rect 247954 7596 247960 7608
rect 219400 7568 247960 7596
rect 219400 7556 219406 7568
rect 247954 7556 247960 7568
rect 248012 7556 248018 7608
rect 248322 7556 248328 7608
rect 248380 7596 248386 7608
rect 290734 7596 290740 7608
rect 248380 7568 290740 7596
rect 248380 7556 248386 7568
rect 290734 7556 290740 7568
rect 290792 7556 290798 7608
rect 291102 7556 291108 7608
rect 291160 7596 291166 7608
rect 351362 7596 351368 7608
rect 291160 7568 351368 7596
rect 291160 7556 291166 7568
rect 351362 7556 351368 7568
rect 351420 7556 351426 7608
rect 398742 7556 398748 7608
rect 398800 7596 398806 7608
rect 508406 7596 508412 7608
rect 398800 7568 508412 7596
rect 398800 7556 398806 7568
rect 508406 7556 508412 7568
rect 508464 7556 508470 7608
rect 209792 7500 219480 7528
rect 219342 7352 219348 7404
rect 219400 7392 219406 7404
rect 219452 7392 219480 7500
rect 219400 7364 219480 7392
rect 219400 7352 219406 7364
rect 186130 6196 186136 6248
rect 186188 6236 186194 6248
rect 201586 6236 201592 6248
rect 186188 6208 201592 6236
rect 186188 6196 186194 6208
rect 201586 6196 201592 6208
rect 201644 6196 201650 6248
rect 176470 6128 176476 6180
rect 176528 6168 176534 6180
rect 187234 6168 187240 6180
rect 176528 6140 187240 6168
rect 176528 6128 176534 6140
rect 187234 6128 187240 6140
rect 187292 6128 187298 6180
rect 201402 6128 201408 6180
rect 201460 6168 201466 6180
rect 222930 6168 222936 6180
rect 201460 6140 222936 6168
rect 201460 6128 201466 6140
rect 222930 6128 222936 6140
rect 222988 6128 222994 6180
rect 226242 6128 226248 6180
rect 226300 6168 226306 6180
rect 258626 6168 258632 6180
rect 226300 6140 258632 6168
rect 226300 6128 226306 6140
rect 258626 6128 258632 6140
rect 258684 6128 258690 6180
rect 260742 6128 260748 6180
rect 260800 6168 260806 6180
rect 308582 6168 308588 6180
rect 260800 6140 308588 6168
rect 260800 6128 260806 6140
rect 308582 6128 308588 6140
rect 308640 6128 308646 6180
rect 309778 6128 309784 6180
rect 309836 6168 309842 6180
rect 376386 6168 376392 6180
rect 309836 6140 376392 6168
rect 309836 6128 309842 6140
rect 376386 6128 376392 6140
rect 376444 6128 376450 6180
rect 386322 6128 386328 6180
rect 386380 6168 386386 6180
rect 490558 6168 490564 6180
rect 386380 6140 490564 6168
rect 386380 6128 386386 6140
rect 490558 6128 490564 6140
rect 490616 6128 490622 6180
rect 280798 4904 280804 4956
rect 280856 4944 280862 4956
rect 280856 4916 291884 4944
rect 280856 4904 280862 4916
rect 188338 4836 188344 4888
rect 188396 4876 188402 4888
rect 190822 4876 190828 4888
rect 188396 4848 190828 4876
rect 188396 4836 188402 4848
rect 190822 4836 190828 4848
rect 190880 4836 190886 4888
rect 291856 4876 291884 4916
rect 330018 4876 330024 4888
rect 291856 4848 330024 4876
rect 330018 4836 330024 4848
rect 330076 4836 330082 4888
rect 352558 4836 352564 4888
rect 352616 4876 352622 4888
rect 358538 4876 358544 4888
rect 352616 4848 358544 4876
rect 352616 4836 352622 4848
rect 358538 4836 358544 4848
rect 358596 4836 358602 4888
rect 173710 4768 173716 4820
rect 173768 4808 173774 4820
rect 183738 4808 183744 4820
rect 173768 4780 183744 4808
rect 173768 4768 173774 4780
rect 183738 4768 183744 4780
rect 183796 4768 183802 4820
rect 194502 4768 194508 4820
rect 194560 4808 194566 4820
rect 212258 4808 212264 4820
rect 194560 4780 212264 4808
rect 194560 4768 194566 4780
rect 212258 4768 212264 4780
rect 212316 4768 212322 4820
rect 221458 4768 221464 4820
rect 221516 4808 221522 4820
rect 240778 4808 240784 4820
rect 221516 4780 240784 4808
rect 221516 4768 221522 4780
rect 240778 4768 240784 4780
rect 240836 4768 240842 4820
rect 242158 4768 242164 4820
rect 242216 4808 242222 4820
rect 255038 4808 255044 4820
rect 242216 4780 255044 4808
rect 242216 4768 242222 4780
rect 255038 4768 255044 4780
rect 255096 4768 255102 4820
rect 255958 4768 255964 4820
rect 256016 4808 256022 4820
rect 280062 4808 280068 4820
rect 256016 4780 280068 4808
rect 256016 4768 256022 4780
rect 280062 4768 280068 4780
rect 280120 4768 280126 4820
rect 309042 4768 309048 4820
rect 309100 4808 309106 4820
rect 378778 4808 378784 4820
rect 309100 4780 378784 4808
rect 309100 4768 309106 4780
rect 378778 4768 378784 4780
rect 378836 4768 378842 4820
rect 382182 4768 382188 4820
rect 382240 4808 382246 4820
rect 483474 4808 483480 4820
rect 382240 4780 483480 4808
rect 382240 4768 382246 4780
rect 483474 4768 483480 4780
rect 483532 4768 483538 4820
rect 192478 4156 192484 4208
rect 192536 4196 192542 4208
rect 194410 4196 194416 4208
rect 192536 4168 194416 4196
rect 192536 4156 192542 4168
rect 194410 4156 194416 4168
rect 194468 4156 194474 4208
rect 213178 4156 213184 4208
rect 213236 4196 213242 4208
rect 215846 4196 215852 4208
rect 213236 4168 215852 4196
rect 213236 4156 213242 4168
rect 215846 4156 215852 4168
rect 215904 4156 215910 4208
rect 425146 4156 425152 4208
rect 425204 4196 425210 4208
rect 426342 4196 426348 4208
rect 425204 4168 426348 4196
rect 425204 4156 425210 4168
rect 426342 4156 426348 4168
rect 426400 4156 426406 4208
rect 451274 4156 451280 4208
rect 451332 4196 451338 4208
rect 452470 4196 452476 4208
rect 451332 4168 452476 4196
rect 451332 4156 451338 4168
rect 452470 4156 452476 4168
rect 452528 4156 452534 4208
rect 127802 4088 127808 4140
rect 127860 4128 127866 4140
rect 134150 4128 134156 4140
rect 127860 4100 134156 4128
rect 127860 4088 127866 4100
rect 134150 4088 134156 4100
rect 134208 4088 134214 4140
rect 144454 4088 144460 4140
rect 144512 4128 144518 4140
rect 146386 4128 146392 4140
rect 144512 4100 146392 4128
rect 144512 4088 144518 4100
rect 146386 4088 146392 4100
rect 146444 4088 146450 4140
rect 160002 4088 160008 4140
rect 160060 4128 160066 4140
rect 163498 4128 163504 4140
rect 160060 4100 163504 4128
rect 160060 4088 160066 4100
rect 163498 4088 163504 4100
rect 163556 4088 163562 4140
rect 166902 4088 166908 4140
rect 166960 4128 166966 4140
rect 172974 4128 172980 4140
rect 166960 4100 172980 4128
rect 166960 4088 166966 4100
rect 172974 4088 172980 4100
rect 173032 4088 173038 4140
rect 361482 4088 361488 4140
rect 361540 4128 361546 4140
rect 453666 4128 453672 4140
rect 361540 4100 453672 4128
rect 361540 4088 361546 4100
rect 453666 4088 453672 4100
rect 453724 4088 453730 4140
rect 130194 4020 130200 4072
rect 130252 4060 130258 4072
rect 135530 4060 135536 4072
rect 130252 4032 135536 4060
rect 130252 4020 130258 4032
rect 135530 4020 135536 4032
rect 135588 4020 135594 4072
rect 140866 4020 140872 4072
rect 140924 4060 140930 4072
rect 143534 4060 143540 4072
rect 140924 4032 143540 4060
rect 140924 4020 140930 4032
rect 143534 4020 143540 4032
rect 143592 4020 143598 4072
rect 159910 4020 159916 4072
rect 159968 4060 159974 4072
rect 162302 4060 162308 4072
rect 159968 4032 162308 4060
rect 159968 4020 159974 4032
rect 162302 4020 162308 4032
rect 162360 4020 162366 4072
rect 364242 4020 364248 4072
rect 364300 4060 364306 4072
rect 457254 4060 457260 4072
rect 364300 4032 457260 4060
rect 364300 4020 364306 4032
rect 457254 4020 457260 4032
rect 457312 4020 457318 4072
rect 128998 3952 129004 4004
rect 129056 3992 129062 4004
rect 135254 3992 135260 4004
rect 129056 3964 135260 3992
rect 129056 3952 129062 3964
rect 135254 3952 135260 3964
rect 135312 3952 135318 4004
rect 176562 3952 176568 4004
rect 176620 3992 176626 4004
rect 186038 3992 186044 4004
rect 176620 3964 186044 3992
rect 176620 3952 176626 3964
rect 186038 3952 186044 3964
rect 186096 3952 186102 4004
rect 367002 3952 367008 4004
rect 367060 3992 367066 4004
rect 460842 3992 460848 4004
rect 367060 3964 460848 3992
rect 367060 3952 367066 3964
rect 460842 3952 460848 3964
rect 460900 3952 460906 4004
rect 139670 3884 139676 3936
rect 139728 3924 139734 3936
rect 142154 3924 142160 3936
rect 139728 3896 142160 3924
rect 139728 3884 139734 3896
rect 142154 3884 142160 3896
rect 142212 3884 142218 3936
rect 169570 3884 169576 3936
rect 169628 3924 169634 3936
rect 176470 3924 176476 3936
rect 169628 3896 176476 3924
rect 169628 3884 169634 3896
rect 176470 3884 176476 3896
rect 176528 3884 176534 3936
rect 177850 3884 177856 3936
rect 177908 3924 177914 3936
rect 188430 3924 188436 3936
rect 177908 3896 188436 3924
rect 177908 3884 177914 3896
rect 188430 3884 188436 3896
rect 188488 3884 188494 3936
rect 195882 3884 195888 3936
rect 195940 3924 195946 3936
rect 214650 3924 214656 3936
rect 195940 3896 214656 3924
rect 195940 3884 195946 3896
rect 214650 3884 214656 3896
rect 214708 3884 214714 3936
rect 368382 3884 368388 3936
rect 368440 3924 368446 3936
rect 464430 3924 464436 3936
rect 368440 3896 464436 3924
rect 368440 3884 368446 3896
rect 464430 3884 464436 3896
rect 464488 3884 464494 3936
rect 142062 3816 142068 3868
rect 142120 3856 142126 3868
rect 143902 3856 143908 3868
rect 142120 3828 143908 3856
rect 142120 3816 142126 3828
rect 143902 3816 143908 3828
rect 143960 3816 143966 3868
rect 169662 3816 169668 3868
rect 169720 3856 169726 3868
rect 177758 3856 177764 3868
rect 169720 3828 177764 3856
rect 169720 3816 169726 3828
rect 177758 3816 177764 3828
rect 177816 3816 177822 3868
rect 182082 3816 182088 3868
rect 182140 3856 182146 3868
rect 195606 3856 195612 3868
rect 182140 3828 195612 3856
rect 182140 3816 182146 3828
rect 195606 3816 195612 3828
rect 195664 3816 195670 3868
rect 198642 3816 198648 3868
rect 198700 3856 198706 3868
rect 218146 3856 218152 3868
rect 198700 3828 218152 3856
rect 198700 3816 198706 3828
rect 218146 3816 218152 3828
rect 218204 3816 218210 3868
rect 373902 3816 373908 3868
rect 373960 3856 373966 3868
rect 471514 3856 471520 3868
rect 373960 3828 471520 3856
rect 373960 3816 373966 3828
rect 471514 3816 471520 3828
rect 471572 3816 471578 3868
rect 143258 3748 143264 3800
rect 143316 3788 143322 3800
rect 144914 3788 144920 3800
rect 143316 3760 144920 3788
rect 143316 3748 143322 3760
rect 144914 3748 144920 3760
rect 144972 3748 144978 3800
rect 182542 3788 182548 3800
rect 177868 3760 182548 3788
rect 173802 3680 173808 3732
rect 173860 3720 173866 3732
rect 177868 3720 177896 3760
rect 182542 3748 182548 3760
rect 182600 3748 182606 3800
rect 183462 3748 183468 3800
rect 183520 3788 183526 3800
rect 196802 3788 196808 3800
rect 183520 3760 196808 3788
rect 183520 3748 183526 3760
rect 196802 3748 196808 3760
rect 196860 3748 196866 3800
rect 200022 3748 200028 3800
rect 200080 3788 200086 3800
rect 221734 3788 221740 3800
rect 200080 3760 221740 3788
rect 200080 3748 200086 3760
rect 221734 3748 221740 3760
rect 221792 3748 221798 3800
rect 371142 3748 371148 3800
rect 371200 3788 371206 3800
rect 467834 3788 467840 3800
rect 371200 3760 467840 3788
rect 371200 3748 371206 3760
rect 467834 3748 467840 3760
rect 467892 3748 467898 3800
rect 173860 3692 177896 3720
rect 173860 3680 173866 3692
rect 180702 3680 180708 3732
rect 180760 3720 180766 3732
rect 193214 3720 193220 3732
rect 180760 3692 193220 3720
rect 180760 3680 180766 3692
rect 193214 3680 193220 3692
rect 193272 3680 193278 3732
rect 205542 3680 205548 3732
rect 205600 3720 205606 3732
rect 228910 3720 228916 3732
rect 205600 3692 228916 3720
rect 205600 3680 205606 3692
rect 228910 3680 228916 3692
rect 228968 3680 228974 3732
rect 379422 3680 379428 3732
rect 379480 3720 379486 3732
rect 478690 3720 478696 3732
rect 379480 3692 478696 3720
rect 379480 3680 379486 3692
rect 478690 3680 478696 3692
rect 478748 3680 478754 3732
rect 168190 3612 168196 3664
rect 168248 3652 168254 3664
rect 174170 3652 174176 3664
rect 168248 3624 174176 3652
rect 168248 3612 168254 3624
rect 174170 3612 174176 3624
rect 174228 3612 174234 3664
rect 175182 3612 175188 3664
rect 175240 3652 175246 3664
rect 184842 3652 184848 3664
rect 175240 3624 184848 3652
rect 175240 3612 175246 3624
rect 184842 3612 184848 3624
rect 184900 3612 184906 3664
rect 186222 3612 186228 3664
rect 186280 3652 186286 3664
rect 200390 3652 200396 3664
rect 186280 3624 200396 3652
rect 186280 3612 186286 3624
rect 200390 3612 200396 3624
rect 200448 3612 200454 3664
rect 202782 3612 202788 3664
rect 202840 3652 202846 3664
rect 225322 3652 225328 3664
rect 202840 3624 225328 3652
rect 202840 3612 202846 3624
rect 225322 3612 225328 3624
rect 225380 3612 225386 3664
rect 376662 3612 376668 3664
rect 376720 3652 376726 3664
rect 475102 3652 475108 3664
rect 376720 3624 475108 3652
rect 376720 3612 376726 3624
rect 475102 3612 475108 3624
rect 475160 3612 475166 3664
rect 132586 3544 132592 3596
rect 132644 3584 132650 3596
rect 138014 3584 138020 3596
rect 132644 3556 138020 3584
rect 132644 3544 132650 3556
rect 138014 3544 138020 3556
rect 138072 3544 138078 3596
rect 138474 3544 138480 3596
rect 138532 3584 138538 3596
rect 142246 3584 142252 3596
rect 138532 3556 142252 3584
rect 138532 3544 138538 3556
rect 142246 3544 142252 3556
rect 142304 3544 142310 3596
rect 146846 3544 146852 3596
rect 146904 3584 146910 3596
rect 147766 3584 147772 3596
rect 146904 3556 147772 3584
rect 146904 3544 146910 3556
rect 147766 3544 147772 3556
rect 147824 3544 147830 3596
rect 150434 3544 150440 3596
rect 150492 3584 150498 3596
rect 151538 3584 151544 3596
rect 150492 3556 151544 3584
rect 150492 3544 150498 3556
rect 151538 3544 151544 3556
rect 151596 3544 151602 3596
rect 161382 3544 161388 3596
rect 161440 3584 161446 3596
rect 164694 3584 164700 3596
rect 161440 3556 164700 3584
rect 161440 3544 161446 3556
rect 164694 3544 164700 3556
rect 164752 3544 164758 3596
rect 165430 3544 165436 3596
rect 165488 3584 165494 3596
rect 170582 3584 170588 3596
rect 165488 3556 170588 3584
rect 165488 3544 165494 3556
rect 170582 3544 170588 3556
rect 170640 3544 170646 3596
rect 172330 3544 172336 3596
rect 172388 3584 172394 3596
rect 181346 3584 181352 3596
rect 172388 3556 181352 3584
rect 172388 3544 172394 3556
rect 181346 3544 181352 3556
rect 181404 3544 181410 3596
rect 187602 3544 187608 3596
rect 187660 3584 187666 3596
rect 203886 3584 203892 3596
rect 187660 3556 203892 3584
rect 187660 3544 187666 3556
rect 203886 3544 203892 3556
rect 203944 3544 203950 3596
rect 208302 3544 208308 3596
rect 208360 3584 208366 3596
rect 232498 3584 232504 3596
rect 208360 3556 232504 3584
rect 208360 3544 208366 3556
rect 232498 3544 232504 3556
rect 232556 3544 232562 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 263410 3584 263416 3596
rect 262272 3556 263416 3584
rect 262272 3544 262278 3556
rect 263410 3544 263416 3556
rect 263468 3544 263474 3596
rect 270494 3544 270500 3596
rect 270552 3584 270558 3596
rect 271690 3584 271696 3596
rect 270552 3556 271696 3584
rect 270552 3544 270558 3556
rect 271690 3544 271696 3556
rect 271748 3544 271754 3596
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 331214 3544 331220 3596
rect 331272 3584 331278 3596
rect 332410 3584 332416 3596
rect 331272 3556 332416 3584
rect 331272 3544 331278 3556
rect 332410 3544 332416 3556
rect 332468 3544 332474 3596
rect 365714 3544 365720 3596
rect 365772 3584 365778 3596
rect 366910 3584 366916 3596
rect 365772 3556 366916 3584
rect 365772 3544 365778 3556
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 373994 3544 374000 3596
rect 374052 3584 374058 3596
rect 375190 3584 375196 3596
rect 374052 3556 375196 3584
rect 374052 3544 374058 3556
rect 375190 3544 375196 3556
rect 375248 3544 375254 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 482278 3584 482284 3596
rect 380860 3556 482284 3584
rect 380860 3544 380866 3556
rect 482278 3544 482284 3556
rect 482336 3544 482342 3596
rect 485774 3544 485780 3596
rect 485832 3584 485838 3596
rect 486970 3584 486976 3596
rect 485832 3556 486976 3584
rect 485832 3544 485838 3556
rect 486970 3544 486976 3556
rect 487028 3544 487034 3596
rect 494146 3544 494152 3596
rect 494204 3584 494210 3596
rect 495342 3584 495348 3596
rect 494204 3556 495348 3584
rect 494204 3544 494210 3556
rect 495342 3544 495348 3556
rect 495400 3544 495406 3596
rect 520274 3544 520280 3596
rect 520332 3584 520338 3596
rect 521470 3584 521476 3596
rect 520332 3556 521476 3584
rect 520332 3544 520338 3556
rect 521470 3544 521476 3556
rect 521528 3544 521534 3596
rect 528554 3544 528560 3596
rect 528612 3584 528618 3596
rect 529842 3584 529848 3596
rect 528612 3556 529848 3584
rect 528612 3544 528618 3556
rect 529842 3544 529848 3556
rect 529900 3544 529906 3596
rect 536926 3544 536932 3596
rect 536984 3584 536990 3596
rect 538122 3584 538128 3596
rect 536984 3556 538128 3584
rect 536984 3544 536990 3556
rect 538122 3544 538128 3556
rect 538180 3544 538186 3596
rect 546494 3544 546500 3596
rect 546552 3584 546558 3596
rect 547690 3584 547696 3596
rect 546552 3556 547696 3584
rect 546552 3544 546558 3556
rect 547690 3544 547696 3556
rect 547748 3544 547754 3596
rect 563146 3544 563152 3596
rect 563204 3584 563210 3596
rect 564342 3584 564348 3596
rect 563204 3556 564348 3584
rect 563204 3544 563210 3556
rect 564342 3544 564348 3556
rect 564400 3544 564406 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 132494 3516 132500 3528
rect 1728 3488 132500 3516
rect 1728 3476 1734 3488
rect 132494 3476 132500 3488
rect 132552 3476 132558 3528
rect 137278 3476 137284 3528
rect 137336 3516 137342 3528
rect 140774 3516 140780 3528
rect 137336 3488 140780 3516
rect 137336 3476 137342 3488
rect 140774 3476 140780 3488
rect 140832 3476 140838 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 152734 3516 152740 3528
rect 151872 3488 152740 3516
rect 151872 3476 151878 3488
rect 152734 3476 152740 3488
rect 152792 3476 152798 3528
rect 153102 3476 153108 3528
rect 153160 3516 153166 3528
rect 153930 3516 153936 3528
rect 153160 3488 153936 3516
rect 153160 3476 153166 3488
rect 153930 3476 153936 3488
rect 153988 3476 153994 3528
rect 155770 3476 155776 3528
rect 155828 3516 155834 3528
rect 156322 3516 156328 3528
rect 155828 3488 156328 3516
rect 155828 3476 155834 3488
rect 156322 3476 156328 3488
rect 156380 3476 156386 3528
rect 157242 3476 157248 3528
rect 157300 3516 157306 3528
rect 158714 3516 158720 3528
rect 157300 3488 158720 3516
rect 157300 3476 157306 3488
rect 158714 3476 158720 3488
rect 158772 3476 158778 3528
rect 162762 3476 162768 3528
rect 162820 3516 162826 3528
rect 167086 3516 167092 3528
rect 162820 3488 167092 3516
rect 162820 3476 162826 3488
rect 167086 3476 167092 3488
rect 167144 3476 167150 3528
rect 168282 3476 168288 3528
rect 168340 3516 168346 3528
rect 175366 3516 175372 3528
rect 168340 3488 175372 3516
rect 168340 3476 168346 3488
rect 175366 3476 175372 3488
rect 175424 3476 175430 3528
rect 177942 3476 177948 3528
rect 178000 3516 178006 3528
rect 189626 3516 189632 3528
rect 178000 3488 189632 3516
rect 178000 3476 178006 3488
rect 189626 3476 189632 3488
rect 189684 3476 189690 3528
rect 190362 3476 190368 3528
rect 190420 3516 190426 3528
rect 201405 3519 201463 3525
rect 201405 3516 201417 3519
rect 190420 3488 201417 3516
rect 190420 3476 190426 3488
rect 201405 3485 201417 3488
rect 201451 3485 201463 3519
rect 201405 3479 201463 3485
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202690 3516 202696 3528
rect 201552 3488 202696 3516
rect 201552 3476 201558 3488
rect 202690 3476 202696 3488
rect 202748 3476 202754 3528
rect 211154 3476 211160 3528
rect 211212 3516 211218 3528
rect 235994 3516 236000 3528
rect 211212 3488 236000 3516
rect 211212 3476 211218 3488
rect 235994 3476 236000 3488
rect 236052 3476 236058 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 252554 3476 252560 3528
rect 252612 3516 252618 3528
rect 253842 3516 253848 3528
rect 252612 3488 253848 3516
rect 252612 3476 252618 3488
rect 253842 3476 253848 3488
rect 253900 3476 253906 3528
rect 287054 3476 287060 3528
rect 287112 3516 287118 3528
rect 288342 3516 288348 3528
rect 287112 3488 288348 3516
rect 287112 3476 287118 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 296714 3476 296720 3528
rect 296772 3516 296778 3528
rect 297910 3516 297916 3528
rect 296772 3488 297916 3516
rect 296772 3476 296778 3488
rect 297910 3476 297916 3488
rect 297968 3476 297974 3528
rect 304994 3476 305000 3528
rect 305052 3516 305058 3528
rect 306190 3516 306196 3528
rect 305052 3488 306196 3516
rect 305052 3476 305058 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 313274 3476 313280 3528
rect 313332 3516 313338 3528
rect 314562 3516 314568 3528
rect 313332 3488 314568 3516
rect 313332 3476 313338 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 347774 3476 347780 3528
rect 347832 3516 347838 3528
rect 349062 3516 349068 3528
rect 347832 3488 349068 3516
rect 347832 3476 347838 3488
rect 349062 3476 349068 3488
rect 349120 3476 349126 3528
rect 356054 3476 356060 3528
rect 356112 3516 356118 3528
rect 357342 3516 357348 3528
rect 356112 3488 357348 3516
rect 356112 3476 356118 3488
rect 357342 3476 357348 3488
rect 357400 3476 357406 3528
rect 446582 3516 446588 3528
rect 357544 3488 446588 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 131114 3448 131120 3460
rect 624 3420 131120 3448
rect 624 3408 630 3420
rect 131114 3408 131120 3420
rect 131172 3408 131178 3460
rect 134886 3408 134892 3460
rect 134944 3448 134950 3460
rect 139394 3448 139400 3460
rect 134944 3420 139400 3448
rect 134944 3408 134950 3420
rect 139394 3408 139400 3420
rect 139452 3408 139458 3460
rect 154482 3408 154488 3460
rect 154540 3448 154546 3460
rect 155126 3448 155132 3460
rect 154540 3420 155132 3448
rect 154540 3408 154546 3420
rect 155126 3408 155132 3420
rect 155184 3408 155190 3460
rect 158622 3408 158628 3460
rect 158680 3448 158686 3460
rect 161106 3448 161112 3460
rect 158680 3420 161112 3448
rect 158680 3408 158686 3420
rect 161106 3408 161112 3420
rect 161164 3408 161170 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 165890 3448 165896 3460
rect 161348 3420 165896 3448
rect 161348 3408 161354 3420
rect 165890 3408 165896 3420
rect 165948 3408 165954 3460
rect 171042 3408 171048 3460
rect 171100 3448 171106 3460
rect 178954 3448 178960 3460
rect 171100 3420 178960 3448
rect 171100 3408 171106 3420
rect 178954 3408 178960 3420
rect 179012 3408 179018 3460
rect 179322 3408 179328 3460
rect 179380 3448 179386 3460
rect 192018 3448 192024 3460
rect 179380 3420 192024 3448
rect 179380 3408 179386 3420
rect 192018 3408 192024 3420
rect 192076 3408 192082 3460
rect 193122 3408 193128 3460
rect 193180 3448 193186 3460
rect 211062 3448 211068 3460
rect 193180 3420 211068 3448
rect 193180 3408 193186 3420
rect 211062 3408 211068 3420
rect 211120 3408 211126 3460
rect 212442 3408 212448 3460
rect 212500 3448 212506 3460
rect 239582 3448 239588 3460
rect 212500 3420 239588 3448
rect 212500 3408 212506 3420
rect 239582 3408 239588 3420
rect 239640 3408 239646 3460
rect 355962 3408 355968 3460
rect 356020 3448 356026 3460
rect 357544 3448 357572 3488
rect 446582 3476 446588 3488
rect 446640 3476 446646 3528
rect 448422 3476 448428 3528
rect 448480 3516 448486 3528
rect 578602 3516 578608 3528
rect 448480 3488 578608 3516
rect 448480 3476 448486 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 578970 3476 578976 3528
rect 579028 3516 579034 3528
rect 580994 3516 581000 3528
rect 579028 3488 581000 3516
rect 579028 3476 579034 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 356020 3420 357572 3448
rect 356020 3408 356026 3420
rect 358722 3408 358728 3460
rect 358780 3448 358786 3460
rect 450170 3448 450176 3460
rect 358780 3420 450176 3448
rect 358780 3408 358786 3420
rect 450170 3408 450176 3420
rect 450228 3408 450234 3460
rect 451182 3408 451188 3460
rect 451240 3448 451246 3460
rect 582190 3448 582196 3460
rect 451240 3420 582196 3448
rect 451240 3408 451246 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 136082 3340 136088 3392
rect 136140 3380 136146 3392
rect 139486 3380 139492 3392
rect 136140 3352 139492 3380
rect 136140 3340 136146 3352
rect 139486 3340 139492 3352
rect 139544 3340 139550 3392
rect 201405 3383 201463 3389
rect 201405 3349 201417 3383
rect 201451 3380 201463 3383
rect 207474 3380 207480 3392
rect 201451 3352 207480 3380
rect 201451 3349 201463 3352
rect 201405 3343 201463 3349
rect 207474 3340 207480 3352
rect 207532 3340 207538 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 416774 3340 416780 3392
rect 416832 3380 416838 3392
rect 417970 3380 417976 3392
rect 416832 3352 417976 3380
rect 416832 3340 416838 3352
rect 417970 3340 417976 3352
rect 418028 3340 418034 3392
rect 433334 3340 433340 3392
rect 433392 3380 433398 3392
rect 434622 3380 434628 3392
rect 433392 3352 434628 3380
rect 433392 3340 433398 3352
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 145650 3272 145656 3324
rect 145708 3312 145714 3324
rect 146294 3312 146300 3324
rect 145708 3284 146300 3312
rect 145708 3272 145714 3284
rect 146294 3272 146300 3284
rect 146352 3272 146358 3324
rect 155862 3272 155868 3324
rect 155920 3312 155926 3324
rect 157518 3312 157524 3324
rect 155920 3284 157524 3312
rect 155920 3272 155926 3284
rect 157518 3272 157524 3284
rect 157576 3272 157582 3324
rect 164050 3272 164056 3324
rect 164108 3312 164114 3324
rect 168190 3312 168196 3324
rect 164108 3284 168196 3312
rect 164108 3272 164114 3284
rect 168190 3272 168196 3284
rect 168248 3272 168254 3324
rect 571334 3272 571340 3324
rect 571392 3312 571398 3324
rect 572622 3312 572628 3324
rect 571392 3284 572628 3312
rect 571392 3272 571398 3284
rect 572622 3272 572628 3284
rect 572680 3272 572686 3324
rect 578878 3272 578884 3324
rect 578936 3312 578942 3324
rect 579798 3312 579804 3324
rect 578936 3284 579804 3312
rect 578936 3272 578942 3284
rect 579798 3272 579804 3284
rect 579856 3272 579862 3324
rect 133782 3204 133788 3256
rect 133840 3244 133846 3256
rect 138290 3244 138296 3256
rect 133840 3216 138296 3244
rect 133840 3204 133846 3216
rect 138290 3204 138296 3216
rect 138348 3204 138354 3256
rect 164142 3136 164148 3188
rect 164200 3176 164206 3188
rect 169386 3176 169392 3188
rect 164200 3148 169392 3176
rect 164200 3136 164206 3148
rect 169386 3136 169392 3148
rect 169444 3136 169450 3188
rect 126606 3068 126612 3120
rect 126664 3108 126670 3120
rect 133874 3108 133880 3120
rect 126664 3080 133880 3108
rect 126664 3068 126670 3080
rect 133874 3068 133880 3080
rect 133932 3068 133938 3120
rect 131390 3000 131396 3052
rect 131448 3040 131454 3052
rect 136634 3040 136640 3052
rect 131448 3012 136640 3040
rect 131448 3000 131454 3012
rect 136634 3000 136640 3012
rect 136692 3000 136698 3052
rect 157150 3000 157156 3052
rect 157208 3040 157214 3052
rect 159910 3040 159916 3052
rect 157208 3012 159916 3040
rect 157208 3000 157214 3012
rect 159910 3000 159916 3012
rect 159968 3000 159974 3052
rect 165522 3000 165528 3052
rect 165580 3040 165586 3052
rect 171778 3040 171784 3052
rect 165580 3012 171784 3040
rect 165580 3000 165586 3012
rect 171778 3000 171784 3012
rect 171836 3000 171842 3052
rect 172422 2932 172428 2984
rect 172480 2972 172486 2984
rect 180150 2972 180156 2984
rect 172480 2944 180156 2972
rect 172480 2932 172486 2944
rect 180150 2932 180156 2944
rect 180208 2932 180214 2984
rect 502334 2728 502340 2780
rect 502392 2768 502398 2780
rect 503622 2768 503628 2780
rect 502392 2740 503628 2768
rect 502392 2728 502398 2740
rect 503622 2728 503628 2740
rect 503680 2728 503686 2780
rect 364334 552 364340 604
rect 364392 592 364398 604
rect 364518 592 364524 604
rect 364392 564 364524 592
rect 364392 552 364398 564
rect 364518 552 364524 564
rect 364576 552 364582 604
rect 367094 552 367100 604
rect 367152 592 367158 604
rect 368014 592 368020 604
rect 367152 564 368020 592
rect 367152 552 367158 564
rect 368014 552 368020 564
rect 368072 552 368078 604
rect 368474 552 368480 604
rect 368532 592 368538 604
rect 369210 592 369216 604
rect 368532 564 369216 592
rect 368532 552 368538 564
rect 369210 552 369216 564
rect 369268 552 369274 604
rect 369854 552 369860 604
rect 369912 592 369918 604
rect 370406 592 370412 604
rect 369912 564 370412 592
rect 369912 552 369918 564
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 372614 552 372620 604
rect 372672 592 372678 604
rect 372798 592 372804 604
rect 372672 564 372804 592
rect 372672 552 372678 564
rect 372798 552 372804 564
rect 372856 552 372862 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 379514 552 379520 604
rect 379572 592 379578 604
rect 379974 592 379980 604
rect 379572 564 379980 592
rect 379572 552 379578 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 500954 552 500960 604
rect 501012 592 501018 604
rect 501230 592 501236 604
rect 501012 564 501236 592
rect 501012 552 501018 564
rect 501230 552 501236 564
rect 501288 552 501294 604
rect 503714 552 503720 604
rect 503772 592 503778 604
rect 504818 592 504824 604
rect 503772 564 504824 592
rect 503772 552 503778 564
rect 504818 552 504824 564
rect 504876 552 504882 604
rect 505094 552 505100 604
rect 505152 592 505158 604
rect 506014 592 506020 604
rect 505152 564 506020 592
rect 505152 552 505158 564
rect 506014 552 506020 564
rect 506072 552 506078 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 576854 552 576860 604
rect 576912 592 576918 604
rect 577406 592 577412 604
rect 576912 564 577412 592
rect 576912 552 576918 564
rect 577406 552 577412 564
rect 577464 552 577470 604
<< via1 >>
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 331220 697552 331272 697604
rect 332508 697552 332560 697604
rect 476764 696940 476816 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 694084 72752 694136
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 347780 692792 347832 692844
rect 348884 692792 348936 692844
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 412824 692724 412876 692776
rect 542544 692724 542596 692776
rect 542728 692724 542780 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 494244 685856 494296 685908
rect 494888 685856 494940 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 429200 684428 429252 684480
rect 429844 684428 429896 684480
rect 558920 684428 558972 684480
rect 559656 684428 559708 684480
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 412640 683068 412692 683120
rect 429200 683068 429252 683120
rect 542360 683068 542412 683120
rect 558920 683068 558972 683120
rect 3332 681708 3384 681760
rect 6184 681708 6236 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 347780 673480 347832 673532
rect 347964 673480 348016 673532
rect 364340 673480 364392 673532
rect 364524 673480 364576 673532
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 483664 673480 483716 673532
rect 580172 673480 580224 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 219072 666544 219124 666596
rect 413100 666544 413152 666596
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 73068 656820 73120 656872
rect 219348 656820 219400 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 284024 654100 284076 654152
rect 284208 654100 284260 654152
rect 347780 654100 347832 654152
rect 347964 654100 348016 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 9036 652740 9088 652792
rect 475384 650020 475436 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 72976 640364 73028 640416
rect 219256 640364 219308 640416
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 72792 640228 72844 640280
rect 219072 640228 219124 640280
rect 72792 637508 72844 637560
rect 72884 637508 72936 637560
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 284024 634788 284076 634840
rect 284208 634788 284260 634840
rect 347780 634788 347832 634840
rect 347964 634788 348016 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 479524 626560 479576 626612
rect 580172 626560 580224 626612
rect 73068 626535 73120 626544
rect 73068 626501 73077 626535
rect 73077 626501 73111 626535
rect 73111 626501 73120 626535
rect 73068 626492 73120 626501
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 9036 624384 9088 624436
rect 129004 624384 129056 624436
rect 3240 623772 3292 623824
rect 8944 623772 8996 623824
rect 73068 616879 73120 616888
rect 73068 616845 73077 616879
rect 73077 616845 73111 616879
rect 73111 616845 73120 616879
rect 73068 616836 73120 616845
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 284024 615476 284076 615528
rect 284208 615476 284260 615528
rect 347780 615476 347832 615528
rect 347964 615476 348016 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 477500 615476 477552 615528
rect 477684 615476 477736 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 73068 611396 73120 611448
rect 219348 611396 219400 611448
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 72884 611260 72936 611312
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 412824 608583 412876 608592
rect 412824 608549 412833 608583
rect 412833 608549 412867 608583
rect 412867 608549 412876 608583
rect 412824 608540 412876 608549
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 542544 608583 542596 608592
rect 542544 608549 542553 608583
rect 542553 608549 542587 608583
rect 542587 608549 542596 608583
rect 542544 608540 542596 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 471244 603100 471296 603152
rect 580172 603100 580224 603152
rect 413008 601672 413060 601724
rect 429568 601672 429620 601724
rect 542728 601672 542780 601724
rect 559288 601672 559340 601724
rect 72976 601536 73028 601588
rect 73160 601536 73212 601588
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 72976 598884 73028 598936
rect 219256 598884 219308 598936
rect 413008 598927 413060 598936
rect 413008 598893 413017 598927
rect 413017 598893 413051 598927
rect 413051 598893 413060 598927
rect 413008 598884 413060 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 542728 598927 542780 598936
rect 542728 598893 542737 598927
rect 542737 598893 542771 598927
rect 542771 598893 542780 598927
rect 542728 598884 542780 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 137744 596164 137796 596216
rect 137928 596164 137980 596216
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 284024 596164 284076 596216
rect 284208 596164 284260 596216
rect 347780 596164 347832 596216
rect 347964 596164 348016 596216
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 477500 596164 477552 596216
rect 477684 596164 477736 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3332 594804 3384 594856
rect 11704 594804 11756 594856
rect 482284 592016 482336 592068
rect 579896 592016 579948 592068
rect 72884 589339 72936 589348
rect 72884 589305 72893 589339
rect 72893 589305 72927 589339
rect 72927 589305 72936 589339
rect 72884 589296 72936 589305
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 413100 589296 413152 589348
rect 429660 589296 429712 589348
rect 542820 589296 542872 589348
rect 559380 589296 559432 589348
rect 8024 589271 8076 589280
rect 8024 589237 8033 589271
rect 8033 589237 8067 589271
rect 8067 589237 8076 589271
rect 8024 589228 8076 589237
rect 137744 589271 137796 589280
rect 137744 589237 137753 589271
rect 137753 589237 137787 589271
rect 137787 589237 137796 589271
rect 137744 589228 137796 589237
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 284024 589271 284076 589280
rect 284024 589237 284033 589271
rect 284033 589237 284067 589271
rect 284067 589237 284076 589271
rect 284024 589228 284076 589237
rect 347872 589228 347924 589280
rect 364432 589228 364484 589280
rect 477592 589228 477644 589280
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 72700 582360 72752 582412
rect 72884 582360 72936 582412
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 413100 582428 413152 582480
rect 429660 582428 429712 582480
rect 542820 582428 542872 582480
rect 559380 582428 559432 582480
rect 413008 582292 413060 582344
rect 429568 582292 429620 582344
rect 542728 582292 542780 582344
rect 559288 582292 559340 582344
rect 8024 579751 8076 579760
rect 8024 579717 8033 579751
rect 8033 579717 8067 579751
rect 8067 579717 8076 579751
rect 8024 579708 8076 579717
rect 137744 579751 137796 579760
rect 137744 579717 137753 579751
rect 137753 579717 137787 579751
rect 137787 579717 137796 579751
rect 137744 579708 137796 579717
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 284024 579751 284076 579760
rect 284024 579717 284033 579751
rect 284033 579717 284067 579751
rect 284067 579717 284076 579751
rect 284024 579708 284076 579717
rect 347780 579683 347832 579692
rect 347780 579649 347789 579683
rect 347789 579649 347823 579683
rect 347823 579649 347832 579683
rect 364340 579683 364392 579692
rect 347780 579640 347832 579649
rect 364340 579649 364349 579683
rect 364349 579649 364383 579683
rect 364383 579649 364392 579683
rect 364340 579640 364392 579649
rect 477500 579683 477552 579692
rect 477500 579649 477509 579683
rect 477509 579649 477543 579683
rect 477543 579649 477552 579683
rect 477500 579640 477552 579649
rect 489184 579640 489236 579692
rect 580172 579640 580224 579692
rect 7932 579572 7984 579624
rect 8116 579572 8168 579624
rect 72700 579572 72752 579624
rect 137652 579572 137704 579624
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 283932 579572 283984 579624
rect 284116 579572 284168 579624
rect 72608 569959 72660 569968
rect 72608 569925 72617 569959
rect 72617 569925 72651 569959
rect 72651 569925 72660 569959
rect 72608 569916 72660 569925
rect 137560 569959 137612 569968
rect 137560 569925 137569 569959
rect 137569 569925 137603 569959
rect 137603 569925 137612 569959
rect 137560 569916 137612 569925
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 347872 569891 347924 569900
rect 347872 569857 347881 569891
rect 347881 569857 347915 569891
rect 347915 569857 347924 569891
rect 347872 569848 347924 569857
rect 364432 569891 364484 569900
rect 364432 569857 364441 569891
rect 364441 569857 364475 569891
rect 364475 569857 364484 569891
rect 364432 569848 364484 569857
rect 477592 569891 477644 569900
rect 477592 569857 477601 569891
rect 477601 569857 477635 569891
rect 477635 569857 477644 569891
rect 477592 569848 477644 569857
rect 494152 569891 494204 569900
rect 494152 569857 494161 569891
rect 494161 569857 494195 569891
rect 494195 569857 494204 569891
rect 494152 569848 494204 569857
rect 4068 567264 4120 567316
rect 10324 567264 10376 567316
rect 412732 563116 412784 563168
rect 429292 563116 429344 563168
rect 542452 563116 542504 563168
rect 559012 563116 559064 563168
rect 72608 563048 72660 563100
rect 137560 563048 137612 563100
rect 218888 563048 218940 563100
rect 348056 563048 348108 563100
rect 364616 563048 364668 563100
rect 7932 562912 7984 562964
rect 8116 562912 8168 562964
rect 72700 562912 72752 562964
rect 137652 562912 137704 562964
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 477776 563048 477828 563100
rect 494336 563048 494388 563100
rect 412732 562980 412784 563032
rect 429292 562980 429344 563032
rect 542452 562980 542504 563032
rect 559012 562980 559064 563032
rect 218980 562912 219032 562964
rect 283932 562912 283984 562964
rect 284116 562912 284168 562964
rect 72700 560235 72752 560244
rect 72700 560201 72709 560235
rect 72709 560201 72743 560235
rect 72743 560201 72752 560235
rect 72700 560192 72752 560201
rect 137652 560235 137704 560244
rect 137652 560201 137661 560235
rect 137661 560201 137695 560235
rect 137695 560201 137704 560235
rect 137652 560192 137704 560201
rect 218980 560235 219032 560244
rect 218980 560201 218989 560235
rect 218989 560201 219023 560235
rect 219023 560201 219032 560235
rect 218980 560192 219032 560201
rect 412732 560235 412784 560244
rect 412732 560201 412741 560235
rect 412741 560201 412775 560235
rect 412775 560201 412784 560235
rect 412732 560192 412784 560201
rect 429292 560235 429344 560244
rect 429292 560201 429301 560235
rect 429301 560201 429335 560235
rect 429335 560201 429344 560235
rect 429292 560192 429344 560201
rect 542452 560235 542504 560244
rect 542452 560201 542461 560235
rect 542461 560201 542495 560235
rect 542495 560201 542504 560235
rect 542452 560192 542504 560201
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 467104 556180 467156 556232
rect 580172 556180 580224 556232
rect 72884 550604 72936 550656
rect 137836 550604 137888 550656
rect 219164 550604 219216 550656
rect 347872 550604 347924 550656
rect 348148 550604 348200 550656
rect 364432 550604 364484 550656
rect 364708 550604 364760 550656
rect 412916 550604 412968 550656
rect 429476 550604 429528 550656
rect 477592 550604 477644 550656
rect 477868 550604 477920 550656
rect 494152 550604 494204 550656
rect 494428 550604 494480 550656
rect 542636 550604 542688 550656
rect 559196 550604 559248 550656
rect 8024 550579 8076 550588
rect 8024 550545 8033 550579
rect 8033 550545 8067 550579
rect 8067 550545 8076 550579
rect 8024 550536 8076 550545
rect 154304 550579 154356 550588
rect 154304 550545 154313 550579
rect 154313 550545 154347 550579
rect 154347 550545 154356 550579
rect 154304 550536 154356 550545
rect 284024 550579 284076 550588
rect 284024 550545 284033 550579
rect 284033 550545 284067 550579
rect 284067 550545 284076 550579
rect 284024 550536 284076 550545
rect 480904 545096 480956 545148
rect 579896 545096 579948 545148
rect 8208 543736 8260 543788
rect 154488 543736 154540 543788
rect 284208 543736 284260 543788
rect 348148 543804 348200 543856
rect 364708 543804 364760 543856
rect 477868 543804 477920 543856
rect 494428 543804 494480 543856
rect 348056 543668 348108 543720
rect 364616 543668 364668 543720
rect 477776 543668 477828 543720
rect 494336 543668 494388 543720
rect 72700 543600 72752 543652
rect 72884 543600 72936 543652
rect 137652 543600 137704 543652
rect 137836 543600 137888 543652
rect 218980 543600 219032 543652
rect 219164 543600 219216 543652
rect 412732 543600 412784 543652
rect 412916 543600 412968 543652
rect 429292 543600 429344 543652
rect 429476 543600 429528 543652
rect 542452 543600 542504 543652
rect 542636 543600 542688 543652
rect 559012 543600 559064 543652
rect 559196 543600 559248 543652
rect 72700 534012 72752 534064
rect 72884 534012 72936 534064
rect 137652 534012 137704 534064
rect 137836 534012 137888 534064
rect 218980 534012 219032 534064
rect 219164 534012 219216 534064
rect 485044 532720 485096 532772
rect 580172 532720 580224 532772
rect 154212 531292 154264 531344
rect 154304 531292 154356 531344
rect 347872 531292 347924 531344
rect 348148 531292 348200 531344
rect 364432 531292 364484 531344
rect 364708 531292 364760 531344
rect 477592 531292 477644 531344
rect 477868 531292 477920 531344
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 72792 524467 72844 524476
rect 72792 524433 72801 524467
rect 72801 524433 72835 524467
rect 72835 524433 72844 524467
rect 72792 524424 72844 524433
rect 137744 524467 137796 524476
rect 137744 524433 137753 524467
rect 137753 524433 137787 524467
rect 137787 524433 137796 524467
rect 137744 524424 137796 524433
rect 154304 524424 154356 524476
rect 219072 524467 219124 524476
rect 219072 524433 219081 524467
rect 219081 524433 219115 524467
rect 219115 524433 219124 524467
rect 219072 524424 219124 524433
rect 8116 524288 8168 524340
rect 8300 524288 8352 524340
rect 154396 524288 154448 524340
rect 284116 524288 284168 524340
rect 284300 524288 284352 524340
rect 72792 521679 72844 521688
rect 72792 521645 72801 521679
rect 72801 521645 72835 521679
rect 72835 521645 72844 521679
rect 72792 521636 72844 521645
rect 137744 521679 137796 521688
rect 137744 521645 137753 521679
rect 137753 521645 137787 521679
rect 137787 521645 137796 521679
rect 137744 521636 137796 521645
rect 219072 521679 219124 521688
rect 219072 521645 219081 521679
rect 219081 521645 219115 521679
rect 219115 521645 219124 521679
rect 219072 521636 219124 521645
rect 347964 521636 348016 521688
rect 348148 521636 348200 521688
rect 364524 521636 364576 521688
rect 364708 521636 364760 521688
rect 477684 521636 477736 521688
rect 477868 521636 477920 521688
rect 494244 521636 494296 521688
rect 494428 521636 494480 521688
rect 284116 516060 284168 516112
rect 291108 516060 291160 516112
rect 106188 515720 106240 515772
rect 196808 515720 196860 515772
rect 385500 515720 385552 515772
rect 462320 515720 462372 515772
rect 89628 515652 89680 515704
rect 185032 515652 185084 515704
rect 397276 515652 397328 515704
rect 477684 515652 477736 515704
rect 72792 515584 72844 515636
rect 173256 515584 173308 515636
rect 202788 515584 202840 515636
rect 244004 515584 244056 515636
rect 409052 515584 409104 515636
rect 494244 515584 494296 515636
rect 41328 515516 41380 515568
rect 161480 515516 161532 515568
rect 171048 515516 171100 515568
rect 232228 515516 232280 515568
rect 350080 515516 350132 515568
rect 397460 515516 397512 515568
rect 420828 515516 420880 515568
rect 527180 515516 527232 515568
rect 24768 515448 24820 515500
rect 149704 515448 149756 515500
rect 154396 515448 154448 515500
rect 220452 515448 220504 515500
rect 235908 515448 235960 515500
rect 267556 515448 267608 515500
rect 326528 515448 326580 515500
rect 347964 515448 348016 515500
rect 361856 515448 361908 515500
rect 412916 515448 412968 515500
rect 432604 515448 432656 515500
rect 542636 515448 542688 515500
rect 8116 515380 8168 515432
rect 137928 515380 137980 515432
rect 138020 515380 138072 515432
rect 208584 515380 208636 515432
rect 219072 515380 219124 515432
rect 255780 515380 255832 515432
rect 267648 515380 267700 515432
rect 279332 515380 279384 515432
rect 314752 515380 314804 515432
rect 331220 515380 331272 515432
rect 338304 515380 338356 515432
rect 364524 515380 364576 515432
rect 373632 515380 373684 515432
rect 429476 515380 429528 515432
rect 444380 515380 444432 515432
rect 559196 515380 559248 515432
rect 300768 514836 300820 514888
rect 302976 514836 303028 514888
rect 3240 509260 3292 509312
rect 7564 509260 7616 509312
rect 462964 509260 463016 509312
rect 580172 509260 580224 509312
rect 6184 509192 6236 509244
rect 128360 509192 128412 509244
rect 453212 509192 453264 509244
rect 476764 509192 476816 509244
rect 3424 502256 3476 502308
rect 128360 502256 128412 502308
rect 453396 502256 453448 502308
rect 580264 502256 580316 502308
rect 460204 498176 460256 498228
rect 580172 498176 580224 498228
rect 453948 495388 454000 495440
rect 483664 495388 483716 495440
rect 453764 488452 453816 488504
rect 475384 488452 475436 488504
rect 456064 485800 456116 485852
rect 580172 485800 580224 485852
rect 8944 485732 8996 485784
rect 128360 485732 128412 485784
rect 453764 481584 453816 481636
rect 580356 481584 580408 481636
rect 3516 478796 3568 478848
rect 128360 478796 128412 478848
rect 453948 473288 454000 473340
rect 479524 473288 479576 473340
rect 11704 470500 11756 470552
rect 128360 470500 128412 470552
rect 452752 466352 452804 466404
rect 471244 466352 471296 466404
rect 10324 463632 10376 463684
rect 128360 463632 128412 463684
rect 543004 462340 543056 462392
rect 580172 462340 580224 462392
rect 453396 459484 453448 459536
rect 482284 459484 482336 459536
rect 3608 455336 3660 455388
rect 128360 455336 128412 455388
rect 453948 452548 454000 452600
rect 489184 452548 489236 452600
rect 3700 448468 3752 448520
rect 128360 448468 128412 448520
rect 453672 445680 453724 445732
rect 467104 445680 467156 445732
rect 7564 440172 7616 440224
rect 128360 440172 128412 440224
rect 453304 438880 453356 438932
rect 579896 438880 579948 438932
rect 453764 438812 453816 438864
rect 480904 438812 480956 438864
rect 3424 433236 3476 433288
rect 128360 433236 128412 433288
rect 453948 430516 454000 430568
rect 485044 430516 485096 430568
rect 3792 425008 3844 425060
rect 128360 425008 128412 425060
rect 453948 423580 454000 423632
rect 462964 423580 463016 423632
rect 3516 418072 3568 418124
rect 128360 418072 128412 418124
rect 453948 416372 454000 416424
rect 460204 416372 460256 416424
rect 3608 409776 3660 409828
rect 128360 409776 128412 409828
rect 453396 409368 453448 409420
rect 456064 409368 456116 409420
rect 3424 402908 3476 402960
rect 128360 402908 128412 402960
rect 453948 402908 454000 402960
rect 543004 402908 543056 402960
rect 453764 395972 453816 396024
rect 580264 395972 580316 396024
rect 3424 394612 3476 394664
rect 128360 394612 128412 394664
rect 460204 391960 460256 392012
rect 580172 391960 580224 392012
rect 3240 380808 3292 380860
rect 129004 380808 129056 380860
rect 453948 380808 454000 380860
rect 578884 380808 578936 380860
rect 453396 373940 453448 373992
rect 580356 373940 580408 373992
rect 3148 367004 3200 367056
rect 129004 367004 129056 367056
rect 453948 366664 454000 366716
rect 460204 366664 460256 366716
rect 453948 360136 454000 360188
rect 580264 360136 580316 360188
rect 453764 353200 453816 353252
rect 580264 353200 580316 353252
rect 3424 347760 3476 347812
rect 128360 347760 128412 347812
rect 453948 345652 454000 345704
rect 580172 345652 580224 345704
rect 3516 338036 3568 338088
rect 129280 338036 129332 338088
rect 8944 332596 8996 332648
rect 128360 332596 128412 332648
rect 7564 324300 7616 324352
rect 128360 324300 128412 324352
rect 3516 324232 3568 324284
rect 129004 324232 129056 324284
rect 453488 322872 453540 322924
rect 580172 322872 580224 322924
rect 453396 311788 453448 311840
rect 580172 311788 580224 311840
rect 11704 309136 11756 309188
rect 128360 309136 128412 309188
rect 3332 309068 3384 309120
rect 129188 309068 129240 309120
rect 453672 302336 453724 302388
rect 456064 302336 456116 302388
rect 6184 302200 6236 302252
rect 128360 302200 128412 302252
rect 453304 299412 453356 299464
rect 579804 299412 579856 299464
rect 13084 287036 13136 287088
rect 128360 287036 128412 287088
rect 453948 280168 454000 280220
rect 461584 280168 461636 280220
rect 3424 280100 3476 280152
rect 129096 280100 129148 280152
rect 3424 277992 3476 278044
rect 128268 277992 128320 278044
rect 453580 275952 453632 276004
rect 580172 275952 580224 276004
rect 3516 266024 3568 266076
rect 8944 266024 8996 266076
rect 453488 264868 453540 264920
rect 580172 264868 580224 264920
rect 8944 263576 8996 263628
rect 128360 263576 128412 263628
rect 453948 259428 454000 259480
rect 471244 259428 471296 259480
rect 10324 256708 10376 256760
rect 128360 256708 128412 256760
rect 456064 252492 456116 252544
rect 579804 252492 579856 252544
rect 3516 251608 3568 251660
rect 7564 251608 7616 251660
rect 453028 251200 453080 251252
rect 457444 251200 457496 251252
rect 15844 241476 15896 241528
rect 128360 241476 128412 241528
rect 453948 237396 454000 237448
rect 469864 237396 469916 237448
rect 3516 237328 3568 237380
rect 129004 237328 129056 237380
rect 14464 233248 14516 233300
rect 128360 233248 128412 233300
rect 453120 230460 453172 230512
rect 474004 230460 474056 230512
rect 453396 229032 453448 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 11704 223524 11756 223576
rect 11704 218016 11756 218068
rect 128360 218016 128412 218068
rect 453304 217948 453356 218000
rect 580172 217948 580224 218000
rect 453764 216792 453816 216844
rect 456064 216792 456116 216844
rect 7564 211148 7616 211200
rect 128360 211148 128412 211200
rect 453948 209788 454000 209840
rect 478144 209788 478196 209840
rect 3148 208156 3200 208208
rect 6184 208156 6236 208208
rect 461584 205572 461636 205624
rect 579804 205572 579856 205624
rect 6184 194556 6236 194608
rect 128636 194556 128688 194608
rect 453948 194556 454000 194608
rect 483664 194556 483716 194608
rect 2872 194488 2924 194540
rect 129372 194488 129424 194540
rect 303896 190340 303948 190392
rect 304816 190340 304868 190392
rect 168656 190272 168708 190324
rect 169576 190272 169628 190324
rect 201592 190204 201644 190256
rect 204904 190204 204956 190256
rect 332784 190204 332836 190256
rect 333888 190204 333940 190256
rect 375656 190204 375708 190256
rect 376668 190204 376720 190256
rect 392124 190204 392176 190256
rect 393136 190204 393188 190256
rect 416872 190204 416924 190256
rect 417976 190204 418028 190256
rect 434996 190204 435048 190256
rect 435916 190204 435968 190256
rect 281632 190136 281684 190188
rect 282736 190136 282788 190188
rect 408592 190136 408644 190188
rect 409696 190136 409748 190188
rect 441620 190136 441672 190188
rect 442816 190136 442868 190188
rect 154672 190068 154724 190120
rect 155776 190068 155828 190120
rect 164516 190068 164568 190120
rect 165436 190068 165488 190120
rect 244556 190068 244608 190120
rect 245476 190068 245528 190120
rect 253572 190068 253624 190120
rect 257344 190068 257396 190120
rect 316224 190068 316276 190120
rect 317236 190068 317288 190120
rect 345112 190068 345164 190120
rect 346216 190068 346268 190120
rect 353392 190068 353444 190120
rect 354496 190068 354548 190120
rect 433340 190068 433392 190120
rect 434536 190068 434588 190120
rect 226340 190000 226392 190052
rect 227536 190000 227588 190052
rect 369860 190000 369912 190052
rect 371056 190000 371108 190052
rect 162860 189932 162912 189984
rect 164056 189932 164108 189984
rect 237932 189932 237984 189984
rect 238668 189932 238720 189984
rect 269212 189932 269264 189984
rect 270316 189932 270368 189984
rect 329472 189932 329524 189984
rect 331864 189932 331916 189984
rect 340972 189932 341024 189984
rect 342076 189932 342128 189984
rect 357532 189932 357584 189984
rect 358636 189932 358688 189984
rect 373172 189932 373224 189984
rect 373908 189932 373960 189984
rect 429200 189932 429252 189984
rect 430396 189932 430448 189984
rect 445760 189932 445812 189984
rect 446956 189932 447008 189984
rect 310520 189864 310572 189916
rect 315304 189864 315356 189916
rect 382280 189864 382332 189916
rect 387064 189864 387116 189916
rect 158720 189796 158772 189848
rect 159916 189796 159968 189848
rect 178500 189796 178552 189848
rect 188344 189796 188396 189848
rect 240416 189796 240468 189848
rect 255964 189796 256016 189848
rect 257712 189796 257764 189848
rect 301504 189796 301556 189848
rect 349252 189796 349304 189848
rect 384304 189796 384356 189848
rect 411076 189796 411128 189848
rect 451924 189796 451976 189848
rect 180984 189728 181036 189780
rect 192484 189728 192536 189780
rect 195888 189728 195940 189780
rect 213184 189728 213236 189780
rect 223120 189728 223172 189780
rect 242164 189728 242216 189780
rect 275008 189728 275060 189780
rect 280804 189728 280856 189780
rect 294788 189728 294840 189780
rect 352564 189728 352616 189780
rect 383844 189728 383896 189780
rect 485780 189728 485832 189780
rect 229652 189660 229704 189712
rect 230388 189660 230440 189712
rect 309692 189660 309744 189712
rect 310428 189660 310480 189712
rect 222292 189456 222344 189508
rect 223488 189456 223540 189508
rect 250260 189456 250312 189508
rect 251088 189456 251140 189508
rect 285772 189456 285824 189508
rect 286968 189456 287020 189508
rect 322020 189456 322072 189508
rect 322848 189456 322900 189508
rect 330300 189456 330352 189508
rect 331128 189456 331180 189508
rect 182640 189388 182692 189440
rect 183468 189388 183520 189440
rect 203248 189388 203300 189440
rect 204168 189388 204220 189440
rect 219808 189388 219860 189440
rect 220636 189388 220688 189440
rect 283288 189388 283340 189440
rect 284208 189388 284260 189440
rect 293960 189388 294012 189440
rect 295248 189388 295300 189440
rect 328644 189388 328696 189440
rect 329748 189388 329800 189440
rect 389640 189388 389692 189440
rect 390468 189388 390520 189440
rect 156236 189320 156288 189372
rect 157248 189320 157300 189372
rect 172796 189320 172848 189372
rect 173808 189320 173860 189372
rect 197544 189320 197596 189372
rect 198648 189320 198700 189372
rect 214012 189320 214064 189372
rect 215208 189320 215260 189372
rect 236276 189320 236328 189372
rect 237288 189320 237340 189372
rect 261024 189320 261076 189372
rect 262128 189320 262180 189372
rect 277492 189320 277544 189372
rect 278688 189320 278740 189372
rect 299756 189320 299808 189372
rect 300768 189320 300820 189372
rect 371516 189320 371568 189372
rect 372528 189320 372580 189372
rect 412732 189320 412784 189372
rect 413928 189320 413980 189372
rect 175280 189252 175332 189304
rect 176568 189252 176620 189304
rect 185124 189252 185176 189304
rect 186228 189252 186280 189304
rect 193404 189252 193456 189304
rect 194508 189252 194560 189304
rect 205732 189252 205784 189304
rect 206928 189252 206980 189304
rect 209872 189252 209924 189304
rect 211068 189252 211120 189304
rect 221464 189252 221516 189304
rect 222844 189252 222896 189304
rect 223856 189252 223908 189304
rect 224868 189252 224920 189304
rect 230480 189252 230532 189304
rect 231768 189252 231820 189304
rect 234620 189252 234672 189304
rect 235908 189252 235960 189304
rect 238760 189252 238812 189304
rect 240048 189252 240100 189304
rect 248604 189252 248656 189304
rect 249708 189252 249760 189304
rect 265164 189252 265216 189304
rect 266268 189252 266320 189304
rect 270868 189252 270920 189304
rect 271972 189252 272024 189304
rect 302240 189252 302292 189304
rect 303528 189252 303580 189304
rect 306380 189252 306432 189304
rect 307668 189252 307720 189304
rect 312176 189252 312228 189304
rect 313188 189252 313240 189304
rect 320364 189252 320416 189304
rect 321468 189252 321520 189304
rect 336924 189252 336976 189304
rect 338028 189252 338080 189304
rect 365720 189252 365772 189304
rect 367008 189252 367060 189304
rect 374000 189252 374052 189304
rect 375288 189252 375340 189304
rect 378140 189252 378192 189304
rect 379428 189252 379480 189304
rect 425152 189252 425204 189304
rect 426348 189252 426400 189304
rect 437480 189252 437532 189304
rect 438768 189252 438820 189304
rect 439136 189252 439188 189304
rect 440056 189252 440108 189304
rect 160376 189116 160428 189168
rect 161388 189116 161440 189168
rect 213552 189116 213604 189168
rect 221464 189116 221516 189168
rect 307208 189116 307260 189168
rect 309784 189116 309836 189168
rect 378968 189116 379020 189168
rect 381544 189116 381596 189168
rect 157892 189048 157944 189100
rect 158628 189048 158680 189100
rect 166172 189048 166224 189100
rect 166908 189048 166960 189100
rect 167000 189048 167052 189100
rect 168196 189048 168248 189100
rect 171140 189048 171192 189100
rect 172428 189048 172480 189100
rect 174452 189048 174504 189100
rect 175188 189048 175240 189100
rect 176936 189048 176988 189100
rect 177856 189048 177908 189100
rect 186780 189048 186832 189100
rect 187516 189048 187568 189100
rect 189264 189048 189316 189100
rect 190276 189048 190328 189100
rect 190920 189048 190972 189100
rect 191748 189048 191800 189100
rect 195060 189048 195112 189100
rect 195888 189048 195940 189100
rect 199200 189048 199252 189100
rect 200764 189048 200816 189100
rect 207388 189048 207440 189100
rect 208308 189048 208360 189100
rect 211528 189048 211580 189100
rect 212356 189048 212408 189100
rect 215668 189048 215720 189100
rect 216588 189048 216640 189100
rect 218152 189048 218204 189100
rect 219348 189048 219400 189100
rect 227996 189048 228048 189100
rect 229008 189048 229060 189100
rect 232136 189048 232188 189100
rect 233056 189048 233108 189100
rect 242900 189048 242952 189100
rect 244188 189048 244240 189100
rect 246120 189048 246172 189100
rect 246948 189048 247000 189100
rect 256884 189048 256936 189100
rect 257988 189048 258040 189100
rect 258540 189048 258592 189100
rect 259276 189048 259328 189100
rect 262680 189048 262732 189100
rect 263508 189048 263560 189100
rect 266820 189048 266872 189100
rect 267556 189048 267608 189100
rect 273352 189048 273404 189100
rect 274548 189048 274600 189100
rect 279148 189048 279200 189100
rect 279976 189048 280028 189100
rect 287428 189048 287480 189100
rect 288348 189048 288400 189100
rect 289912 189048 289964 189100
rect 291108 189048 291160 189100
rect 291568 189048 291620 189100
rect 292396 189048 292448 189100
rect 293132 189048 293184 189100
rect 293868 189048 293920 189100
rect 295616 189048 295668 189100
rect 296628 189048 296680 189100
rect 298100 189048 298152 189100
rect 299388 189048 299440 189100
rect 301412 189048 301464 189100
rect 302148 189048 302200 189100
rect 308036 189048 308088 189100
rect 308956 189048 309008 189100
rect 324504 189048 324556 189100
rect 327724 189048 327776 189100
rect 338488 189048 338540 189100
rect 339316 189048 339368 189100
rect 342628 189048 342680 189100
rect 344284 189048 344336 189100
rect 346768 189048 346820 189100
rect 348424 189048 348476 189100
rect 350908 189048 350960 189100
rect 351736 189048 351788 189100
rect 355048 189048 355100 189100
rect 355876 189048 355928 189100
rect 359188 189048 359240 189100
rect 360108 189048 360160 189100
rect 361580 189048 361632 189100
rect 362868 189048 362920 189100
rect 363236 189048 363288 189100
rect 364248 189048 364300 189100
rect 364892 189048 364944 189100
rect 365628 189048 365680 189100
rect 379796 189048 379848 189100
rect 380716 189048 380768 189100
rect 381452 189048 381504 189100
rect 382188 189048 382240 189100
rect 385500 189048 385552 189100
rect 386236 189048 386288 189100
rect 387984 189048 388036 189100
rect 388996 189048 389048 189100
rect 400404 189048 400456 189100
rect 401508 189048 401560 189100
rect 402060 189048 402112 189100
rect 402888 189048 402940 189100
rect 404544 189048 404596 189100
rect 405556 189048 405608 189100
rect 410248 189048 410300 189100
rect 411168 189048 411220 189100
rect 414388 189048 414440 189100
rect 416044 189048 416096 189100
rect 418528 189048 418580 189100
rect 420184 189048 420236 189100
rect 421012 189048 421064 189100
rect 422116 189048 422168 189100
rect 422668 189048 422720 189100
rect 423496 189048 423548 189100
rect 426808 189048 426860 189100
rect 427636 189048 427688 189100
rect 428372 189048 428424 189100
rect 429108 189048 429160 189100
rect 430856 189048 430908 189100
rect 431776 189048 431828 189100
rect 436652 189048 436704 189100
rect 437388 189048 437440 189100
rect 443276 189048 443328 189100
rect 444196 189048 444248 189100
rect 444932 189048 444984 189100
rect 445668 189048 445720 189100
rect 447416 189048 447468 189100
rect 448428 189048 448480 189100
rect 449900 189048 449952 189100
rect 451188 189048 451240 189100
rect 220728 188300 220780 188352
rect 251180 188300 251232 188352
rect 252744 188300 252796 188352
rect 296720 188300 296772 188352
rect 388812 188300 388864 188352
rect 494060 188300 494112 188352
rect 235448 186940 235500 186992
rect 271880 186940 271932 186992
rect 271972 186940 272024 186992
rect 322940 186940 322992 186992
rect 393780 186940 393832 186992
rect 500960 186940 501012 186992
rect 147680 185580 147732 185632
rect 148508 185580 148560 185632
rect 150440 185580 150492 185632
rect 151084 185580 151136 185632
rect 396264 185580 396316 185632
rect 503720 185580 503772 185632
rect 401232 184152 401284 184204
rect 512000 184152 512052 184204
rect 135536 183472 135588 183524
rect 135628 183472 135680 183524
rect 406108 182792 406160 182844
rect 518900 182792 518952 182844
rect 453672 182112 453724 182164
rect 580172 182112 580224 182164
rect 142160 181432 142212 181484
rect 142804 181432 142856 181484
rect 367376 181432 367428 181484
rect 462320 181432 462372 181484
rect 146300 180888 146352 180940
rect 146852 180888 146904 180940
rect 3240 180752 3292 180804
rect 13084 180752 13136 180804
rect 409696 180072 409748 180124
rect 521660 180072 521712 180124
rect 223488 178644 223540 178696
rect 252560 178644 252612 178696
rect 259276 178644 259328 178696
rect 305000 178644 305052 178696
rect 318616 178644 318668 178696
rect 390560 178644 390612 178696
rect 413836 178644 413888 178696
rect 528560 178644 528612 178696
rect 227536 177284 227588 177336
rect 259460 177284 259512 177336
rect 335176 177284 335228 177336
rect 415400 177284 415452 177336
rect 420184 177284 420236 177336
rect 536840 177284 536892 177336
rect 422116 175924 422168 175976
rect 539600 175924 539652 175976
rect 426256 174496 426308 174548
rect 546500 174496 546552 174548
rect 143908 173884 143960 173936
rect 144184 173884 144236 173936
rect 431776 173136 431828 173188
rect 554780 173136 554832 173188
rect 434536 171776 434588 171828
rect 557540 171776 557592 171828
rect 453580 171028 453632 171080
rect 580172 171028 580224 171080
rect 438676 168988 438728 169040
rect 564440 168988 564492 169040
rect 444196 167628 444248 167680
rect 571340 167628 571392 167680
rect 354496 166268 354548 166320
rect 443000 166268 443052 166320
rect 446956 166268 447008 166320
rect 575480 166268 575532 166320
rect 448336 164840 448388 164892
rect 578884 164840 578936 164892
rect 143632 164160 143684 164212
rect 143816 164160 143868 164212
rect 364156 163480 364208 163532
rect 458180 163480 458232 163532
rect 366916 162120 366968 162172
rect 460940 162120 460992 162172
rect 376576 160692 376628 160744
rect 476120 160692 476172 160744
rect 381544 159332 381596 159384
rect 478880 159332 478932 159384
rect 471244 158652 471296 158704
rect 579804 158652 579856 158704
rect 365628 157972 365680 158024
rect 459652 157972 459704 158024
rect 387064 156612 387116 156664
rect 484400 156612 484452 156664
rect 384948 155184 385000 155236
rect 487160 155184 487212 155236
rect 135352 154547 135404 154556
rect 135352 154513 135361 154547
rect 135361 154513 135395 154547
rect 135395 154513 135404 154547
rect 135352 154504 135404 154513
rect 393136 153824 393188 153876
rect 498200 153824 498252 153876
rect 397368 152464 397420 152516
rect 505100 152464 505152 152516
rect 3148 151716 3200 151768
rect 129280 151716 129332 151768
rect 405556 151036 405608 151088
rect 516140 151036 516192 151088
rect 416044 149676 416096 149728
rect 529940 149676 529992 149728
rect 417976 148316 418028 148368
rect 534080 148316 534132 148368
rect 135444 147568 135496 147620
rect 427636 146888 427688 146940
rect 547880 146888 547932 146940
rect 430396 145528 430448 145580
rect 552020 145528 552072 145580
rect 437388 144168 437440 144220
rect 563060 144168 563112 144220
rect 135444 143488 135496 143540
rect 143816 143531 143868 143540
rect 143816 143497 143825 143531
rect 143825 143497 143859 143531
rect 143859 143497 143868 143531
rect 143816 143488 143868 143497
rect 440056 142808 440108 142860
rect 565820 142808 565872 142860
rect 442816 141380 442868 141432
rect 569960 141380 570012 141432
rect 371056 140020 371108 140072
rect 466460 140020 466512 140072
rect 380716 138660 380768 138712
rect 480260 138660 480312 138712
rect 386236 137232 386288 137284
rect 488540 137232 488592 137284
rect 3424 136484 3476 136536
rect 8944 136484 8996 136536
rect 390376 135872 390428 135924
rect 495440 135872 495492 135924
rect 457444 135192 457496 135244
rect 580172 135192 580224 135244
rect 398656 133152 398708 133204
rect 506480 133152 506532 133204
rect 401508 131724 401560 131776
rect 510620 131724 510672 131776
rect 135628 131452 135680 131504
rect 402796 130364 402848 130416
rect 513380 130364 513432 130416
rect 415308 129004 415360 129056
rect 531320 129004 531372 129056
rect 143816 128299 143868 128308
rect 143816 128265 143825 128299
rect 143825 128265 143859 128299
rect 143859 128265 143868 128299
rect 143816 128256 143868 128265
rect 423496 127576 423548 127628
rect 542360 127576 542412 127628
rect 433248 126216 433300 126268
rect 556160 126216 556212 126268
rect 435916 124856 435968 124908
rect 560300 124856 560352 124908
rect 135628 124108 135680 124160
rect 135812 124108 135864 124160
rect 453488 124108 453540 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 10324 122748 10376 122800
rect 135812 122748 135864 122800
rect 351736 113772 351788 113824
rect 438860 113772 438912 113824
rect 343548 112412 343600 112464
rect 427820 112412 427872 112464
rect 469864 111732 469916 111784
rect 579804 111732 579856 111784
rect 372436 111052 372488 111104
rect 469220 111052 469272 111104
rect 333796 109692 333848 109744
rect 414020 109692 414072 109744
rect 3240 108944 3292 108996
rect 129188 108944 129240 108996
rect 331036 108264 331088 108316
rect 409880 108264 409932 108316
rect 342076 106904 342128 106956
rect 425060 106904 425112 106956
rect 135628 106199 135680 106208
rect 135628 106165 135637 106199
rect 135637 106165 135671 106199
rect 135671 106165 135680 106199
rect 135628 106156 135680 106165
rect 349068 105544 349120 105596
rect 434720 105544 434772 105596
rect 135628 104839 135680 104848
rect 135628 104805 135637 104839
rect 135637 104805 135671 104839
rect 135671 104805 135680 104839
rect 135628 104796 135680 104805
rect 331864 104116 331916 104168
rect 408500 104116 408552 104168
rect 339316 102756 339368 102808
rect 420920 102756 420972 102808
rect 336648 101396 336700 101448
rect 416780 101396 416832 101448
rect 329748 99968 329800 100020
rect 407120 99968 407172 100020
rect 326896 98608 326948 98660
rect 402980 98608 403032 98660
rect 324228 97248 324280 97300
rect 400220 97248 400272 97300
rect 321376 95888 321428 95940
rect 396080 95888 396132 95940
rect 318708 94460 318760 94512
rect 391940 94460 391992 94512
rect 3424 93780 3476 93832
rect 15844 93780 15896 93832
rect 317236 93100 317288 93152
rect 389180 93100 389232 93152
rect 314476 91740 314528 91792
rect 385040 91740 385092 91792
rect 328368 90312 328420 90364
rect 405740 90312 405792 90364
rect 135536 89632 135588 89684
rect 311808 88952 311860 89004
rect 382280 88952 382332 89004
rect 474004 88272 474056 88324
rect 580172 88272 580224 88324
rect 375196 87592 375248 87644
rect 473360 87592 473412 87644
rect 135444 86912 135496 86964
rect 135720 86912 135772 86964
rect 143724 86912 143776 86964
rect 304816 86232 304868 86284
rect 371240 86232 371292 86284
rect 408408 86232 408460 86284
rect 520280 86232 520332 86284
rect 135720 85527 135772 85536
rect 135720 85493 135729 85527
rect 135729 85493 135763 85527
rect 135763 85493 135772 85527
rect 135720 85484 135772 85493
rect 307668 84804 307720 84856
rect 374000 84804 374052 84856
rect 427728 84804 427780 84856
rect 549260 84804 549312 84856
rect 302148 83444 302200 83496
rect 367100 83444 367152 83496
rect 420828 83444 420880 83496
rect 538220 83444 538272 83496
rect 299296 82084 299348 82136
rect 364340 82084 364392 82136
rect 395988 82084 396040 82136
rect 502340 82084 502392 82136
rect 295248 80656 295300 80708
rect 356060 80656 356112 80708
rect 362776 80656 362828 80708
rect 455420 80656 455472 80708
rect 3424 79976 3476 80028
rect 14464 79976 14516 80028
rect 292396 79296 292448 79348
rect 353300 79296 353352 79348
rect 355876 79296 355928 79348
rect 444380 79296 444432 79348
rect 445668 79296 445720 79348
rect 574100 79296 574152 79348
rect 289728 77936 289780 77988
rect 349160 77936 349212 77988
rect 360016 77936 360068 77988
rect 451280 77936 451332 77988
rect 135720 77299 135772 77308
rect 135720 77265 135729 77299
rect 135729 77265 135763 77299
rect 135763 77265 135772 77299
rect 135720 77256 135772 77265
rect 143632 77299 143684 77308
rect 143632 77265 143641 77299
rect 143641 77265 143675 77299
rect 143675 77265 143684 77299
rect 143632 77256 143684 77265
rect 453396 77188 453448 77240
rect 580172 77188 580224 77240
rect 286876 76508 286928 76560
rect 346400 76508 346452 76560
rect 353208 76508 353260 76560
rect 441620 76508 441672 76560
rect 284116 75148 284168 75200
rect 342260 75148 342312 75200
rect 347688 75148 347740 75200
rect 433340 75148 433392 75200
rect 279976 73788 280028 73840
rect 335360 73788 335412 73840
rect 346216 73788 346268 73840
rect 430580 73788 430632 73840
rect 282736 72428 282788 72480
rect 339500 72428 339552 72480
rect 344284 72428 344336 72480
rect 426440 72428 426492 72480
rect 442908 72428 442960 72480
rect 571432 72428 571484 72480
rect 277308 71000 277360 71052
rect 331220 71000 331272 71052
rect 340788 71000 340840 71052
rect 423680 71000 423732 71052
rect 440148 71000 440200 71052
rect 567200 71000 567252 71052
rect 274456 69640 274508 69692
rect 328460 69640 328512 69692
rect 337936 69640 337988 69692
rect 419540 69640 419592 69692
rect 438768 69640 438820 69692
rect 563152 69640 563204 69692
rect 271788 68280 271840 68332
rect 324320 68280 324372 68332
rect 335268 68280 335320 68332
rect 416872 68280 416924 68332
rect 418068 68280 418120 68332
rect 535460 68280 535512 68332
rect 270316 66852 270368 66904
rect 321560 66852 321612 66904
rect 333888 66852 333940 66904
rect 412640 66852 412692 66904
rect 430488 66852 430540 66904
rect 553400 66852 553452 66904
rect 135444 66240 135496 66292
rect 135720 66240 135772 66292
rect 267556 65492 267608 65544
rect 317420 65492 317472 65544
rect 322756 65492 322808 65544
rect 398840 65492 398892 65544
rect 426348 65492 426400 65544
rect 546592 65492 546644 65544
rect 3332 64812 3384 64864
rect 129096 64812 129148 64864
rect 456064 64812 456116 64864
rect 579804 64812 579856 64864
rect 264888 64132 264940 64184
rect 313280 64132 313332 64184
rect 321468 64132 321520 64184
rect 394700 64132 394752 64184
rect 313096 62772 313148 62824
rect 383660 62772 383712 62824
rect 405648 62772 405700 62824
rect 517520 62772 517572 62824
rect 262036 61344 262088 61396
rect 310520 61344 310572 61396
rect 315304 61344 315356 61396
rect 380900 61344 380952 61396
rect 413928 61344 413980 61396
rect 528652 61344 528704 61396
rect 135444 60843 135496 60852
rect 135444 60809 135453 60843
rect 135453 60809 135487 60843
rect 135487 60809 135496 60843
rect 135444 60800 135496 60809
rect 143724 60664 143776 60716
rect 143908 60664 143960 60716
rect 308956 59984 309008 60036
rect 376760 59984 376812 60036
rect 411168 59984 411220 60036
rect 524420 59984 524472 60036
rect 257988 58624 258040 58676
rect 303620 58624 303672 58676
rect 306288 58624 306340 58676
rect 374092 58624 374144 58676
rect 393228 58624 393280 58676
rect 499580 58624 499632 58676
rect 135444 57919 135496 57928
rect 135444 57885 135453 57919
rect 135453 57885 135487 57919
rect 135487 57885 135496 57919
rect 135444 57876 135496 57885
rect 143908 57876 143960 57928
rect 255136 57196 255188 57248
rect 299480 57196 299532 57248
rect 303436 57196 303488 57248
rect 369860 57196 369912 57248
rect 383568 57196 383620 57248
rect 485872 57196 485924 57248
rect 252468 55836 252520 55888
rect 296812 55836 296864 55888
rect 300676 55836 300728 55888
rect 365720 55836 365772 55888
rect 388996 55836 389048 55888
rect 492680 55836 492732 55888
rect 249616 54476 249668 54528
rect 292580 54476 292632 54528
rect 299388 54476 299440 54528
rect 362960 54476 363012 54528
rect 378048 54476 378100 54528
rect 477592 54476 477644 54528
rect 246856 53048 246908 53100
rect 288440 53048 288492 53100
rect 293868 53048 293920 53100
rect 356152 53048 356204 53100
rect 358636 53048 358688 53100
rect 448520 53048 448572 53100
rect 291016 51756 291068 51808
rect 351920 51756 351972 51808
rect 245476 51688 245528 51740
rect 285680 51688 285732 51740
rect 350448 51688 350500 51740
rect 437480 51688 437532 51740
rect 444288 51688 444340 51740
rect 572720 51688 572772 51740
rect 3424 51008 3476 51060
rect 11704 51008 11756 51060
rect 288256 50396 288308 50448
rect 347780 50396 347832 50448
rect 242808 50328 242860 50380
rect 281540 50328 281592 50380
rect 346308 50328 346360 50380
rect 431960 50328 432012 50380
rect 434628 50328 434680 50380
rect 558920 50328 558972 50380
rect 239956 48968 240008 49020
rect 278780 48968 278832 49020
rect 284208 48968 284260 49020
rect 340880 48968 340932 49020
rect 409788 48968 409840 49020
rect 523040 48968 523092 49020
rect 143724 48331 143776 48340
rect 143724 48297 143733 48331
rect 143733 48297 143767 48331
rect 143767 48297 143776 48331
rect 143724 48288 143776 48297
rect 331128 47608 331180 47660
rect 408592 47608 408644 47660
rect 237196 47540 237248 47592
rect 274640 47540 274692 47592
rect 275928 47540 275980 47592
rect 331312 47540 331364 47592
rect 407028 47540 407080 47592
rect 520372 47540 520424 47592
rect 235908 46180 235960 46232
rect 270500 46180 270552 46232
rect 278596 46180 278648 46232
rect 333980 46180 334032 46232
rect 375288 46180 375340 46232
rect 471980 46180 472032 46232
rect 274548 44888 274600 44940
rect 327080 44888 327132 44940
rect 233056 44820 233108 44872
rect 267740 44820 267792 44872
rect 325608 44820 325660 44872
rect 401600 44820 401652 44872
rect 424968 44820 425020 44872
rect 545120 44820 545172 44872
rect 269028 43392 269080 43444
rect 320180 43392 320232 43444
rect 360108 43392 360160 43444
rect 451372 43392 451424 43444
rect 266176 42100 266228 42152
rect 316040 42100 316092 42152
rect 230388 42032 230440 42084
rect 263600 42032 263652 42084
rect 315948 42032 316000 42084
rect 387800 42032 387852 42084
rect 402888 42032 402940 42084
rect 512092 42032 512144 42084
rect 478144 41352 478196 41404
rect 580172 41352 580224 41404
rect 227628 40672 227680 40724
rect 260840 40672 260892 40724
rect 263416 40672 263468 40724
rect 313372 40672 313424 40724
rect 354588 40672 354640 40724
rect 443092 40672 443144 40724
rect 262128 39380 262180 39432
rect 309140 39380 309192 39432
rect 224776 39312 224828 39364
rect 256700 39312 256752 39364
rect 296536 39312 296588 39364
rect 360200 39312 360252 39364
rect 362868 39312 362920 39364
rect 454040 39312 454092 39364
rect 143724 38632 143776 38684
rect 143908 38632 143960 38684
rect 256608 37884 256660 37936
rect 302240 37884 302292 37936
rect 342168 37884 342220 37936
rect 425152 37884 425204 37936
rect 431868 37884 431920 37936
rect 554872 37884 554924 37936
rect 296628 36592 296680 36644
rect 358820 36592 358872 36644
rect 220636 36524 220688 36576
rect 249800 36524 249852 36576
rect 250996 36524 251048 36576
rect 295340 36524 295392 36576
rect 357348 36524 357400 36576
rect 447140 36524 447192 36576
rect 449808 36524 449860 36576
rect 578976 36524 579028 36576
rect 3424 35844 3476 35896
rect 7564 35844 7616 35896
rect 249708 35164 249760 35216
rect 291200 35164 291252 35216
rect 317328 35164 317380 35216
rect 390652 35164 390704 35216
rect 394608 35164 394660 35216
rect 502432 35164 502484 35216
rect 246948 33804 247000 33856
rect 287060 33804 287112 33856
rect 217968 33736 218020 33788
rect 245660 33736 245712 33788
rect 286968 33736 287020 33788
rect 345020 33736 345072 33788
rect 351828 33736 351880 33788
rect 440240 33736 440292 33788
rect 447048 33736 447100 33788
rect 576860 33736 576912 33788
rect 215116 32376 215168 32428
rect 242900 32376 242952 32428
rect 244096 32376 244148 32428
rect 284300 32376 284352 32428
rect 314568 32376 314620 32428
rect 386420 32376 386472 32428
rect 387708 32376 387760 32428
rect 491300 32376 491352 32428
rect 241428 31016 241480 31068
rect 280160 31016 280212 31068
rect 281448 31016 281500 31068
rect 338120 31016 338172 31068
rect 348424 31016 348476 31068
rect 433432 31016 433484 31068
rect 441528 31016 441580 31068
rect 568580 31016 568632 31068
rect 453304 30268 453356 30320
rect 580172 30268 580224 30320
rect 240048 29588 240100 29640
rect 277400 29588 277452 29640
rect 304908 29588 304960 29640
rect 372620 29588 372672 29640
rect 259368 28296 259420 28348
rect 306380 28296 306432 28348
rect 234528 28228 234580 28280
rect 270592 28228 270644 28280
rect 303528 28228 303580 28280
rect 368480 28228 368532 28280
rect 369768 28228 369820 28280
rect 465080 28228 465132 28280
rect 135444 27548 135496 27600
rect 143724 27548 143776 27600
rect 144000 27548 144052 27600
rect 224868 26868 224920 26920
rect 255320 26868 255372 26920
rect 257344 26868 257396 26920
rect 298100 26868 298152 26920
rect 300768 26868 300820 26920
rect 365812 26868 365864 26920
rect 372528 26868 372580 26920
rect 467932 26868 467984 26920
rect 212356 25576 212408 25628
rect 237380 25576 237432 25628
rect 237288 25508 237340 25560
rect 273260 25508 273312 25560
rect 298008 25508 298060 25560
rect 361580 25508 361632 25560
rect 429108 25508 429160 25560
rect 550640 25508 550692 25560
rect 339408 24148 339460 24200
rect 422300 24148 422352 24200
rect 206836 24080 206888 24132
rect 230480 24080 230532 24132
rect 231676 24080 231728 24132
rect 266360 24080 266412 24132
rect 282828 24080 282880 24132
rect 339592 24080 339644 24132
rect 422208 24080 422260 24132
rect 540980 24080 541032 24132
rect 204076 22720 204128 22772
rect 227812 22720 227864 22772
rect 228916 22720 228968 22772
rect 262220 22720 262272 22772
rect 280068 22720 280120 22772
rect 336740 22720 336792 22772
rect 338028 22720 338080 22772
rect 418160 22720 418212 22772
rect 419448 22720 419500 22772
rect 536932 22720 536984 22772
rect 3148 22040 3200 22092
rect 129004 22040 129056 22092
rect 204904 21428 204956 21480
rect 223580 21428 223632 21480
rect 278688 21428 278740 21480
rect 332600 21428 332652 21480
rect 222844 21360 222896 21412
rect 252652 21360 252704 21412
rect 332508 21360 332560 21412
rect 411260 21360 411312 21412
rect 412548 21360 412600 21412
rect 527180 21360 527232 21412
rect 200764 20000 200816 20052
rect 219440 20000 219492 20052
rect 219256 19932 219308 19984
rect 248420 19932 248472 19984
rect 266268 19932 266320 19984
rect 314660 19932 314712 19984
rect 326988 19932 327040 19984
rect 404360 19932 404412 19984
rect 416688 19932 416740 19984
rect 532700 19932 532752 19984
rect 301504 19252 301556 19304
rect 305092 19252 305144 19304
rect 197268 18640 197320 18692
rect 216680 18640 216732 18692
rect 216496 18572 216548 18624
rect 244280 18572 244332 18624
rect 255228 18572 255280 18624
rect 300860 18572 300912 18624
rect 310428 18572 310480 18624
rect 379520 18572 379572 18624
rect 390468 18572 390520 18624
rect 494152 18572 494204 18624
rect 483664 17892 483716 17944
rect 579804 17892 579856 17944
rect 251088 17280 251140 17332
rect 293960 17280 294012 17332
rect 194416 17212 194468 17264
rect 212540 17212 212592 17264
rect 215208 17212 215260 17264
rect 241520 17212 241572 17264
rect 292488 17212 292540 17264
rect 354680 17212 354732 17264
rect 384304 17212 384356 17264
rect 436100 17212 436152 17264
rect 209688 15920 209740 15972
rect 234620 15920 234672 15972
rect 191656 15852 191708 15904
rect 209872 15852 209924 15904
rect 233148 15852 233200 15904
rect 269120 15852 269172 15904
rect 270408 15852 270460 15904
rect 321652 15852 321704 15904
rect 322848 15852 322900 15904
rect 397460 15852 397512 15904
rect 400128 15852 400180 15904
rect 509240 15852 509292 15904
rect 288348 14492 288400 14544
rect 347872 14492 347924 14544
rect 190276 14424 190328 14476
rect 205640 14424 205692 14476
rect 216588 14424 216640 14476
rect 244372 14424 244424 14476
rect 245568 14424 245620 14476
rect 287152 14424 287204 14476
rect 344928 14424 344980 14476
rect 429200 14424 429252 14476
rect 436008 14424 436060 14476
rect 561680 14424 561732 14476
rect 187516 13064 187568 13116
rect 201500 13064 201552 13116
rect 208216 13064 208268 13116
rect 233240 13064 233292 13116
rect 244188 13064 244240 13116
rect 282920 13064 282972 13116
rect 285588 13064 285640 13116
rect 343640 13064 343692 13116
rect 404268 13064 404320 13116
rect 514760 13064 514812 13116
rect 135536 11747 135588 11756
rect 135536 11713 135545 11747
rect 135545 11713 135579 11747
rect 135579 11713 135588 11747
rect 135536 11704 135588 11713
rect 184848 11704 184900 11756
rect 198740 11704 198792 11756
rect 204168 11704 204220 11756
rect 226340 11704 226392 11756
rect 229008 11704 229060 11756
rect 262312 11704 262364 11756
rect 263508 11704 263560 11756
rect 311900 11704 311952 11756
rect 313188 11704 313240 11756
rect 382372 11704 382424 11756
rect 391848 11704 391900 11756
rect 496820 11704 496872 11756
rect 188988 10276 189040 10328
rect 204260 10276 204312 10328
rect 206928 10276 206980 10328
rect 229100 10276 229152 10328
rect 231768 10276 231820 10328
rect 264980 10276 265032 10328
rect 267648 10276 267700 10328
rect 318800 10276 318852 10328
rect 320088 10276 320140 10328
rect 393320 10276 393372 10328
rect 423588 10276 423640 10328
rect 543740 10276 543792 10328
rect 238668 8984 238720 9036
rect 276480 8984 276532 9036
rect 191748 8916 191800 8968
rect 208676 8916 208728 8968
rect 210976 8916 211028 8968
rect 237196 8916 237248 8968
rect 273168 8916 273220 8968
rect 326436 8916 326488 8968
rect 327724 8916 327776 8968
rect 401324 8916 401376 8968
rect 451924 8916 451976 8968
rect 526260 8916 526312 8968
rect 2780 8100 2832 8152
rect 6184 8100 6236 8152
rect 183376 7556 183428 7608
rect 198004 7556 198056 7608
rect 198556 7556 198608 7608
rect 219348 7556 219400 7608
rect 247960 7556 248012 7608
rect 248328 7556 248380 7608
rect 290740 7556 290792 7608
rect 291108 7556 291160 7608
rect 351368 7556 351420 7608
rect 398748 7556 398800 7608
rect 508412 7556 508464 7608
rect 219348 7352 219400 7404
rect 186136 6196 186188 6248
rect 201592 6196 201644 6248
rect 176476 6128 176528 6180
rect 187240 6128 187292 6180
rect 201408 6128 201460 6180
rect 222936 6128 222988 6180
rect 226248 6128 226300 6180
rect 258632 6128 258684 6180
rect 260748 6128 260800 6180
rect 308588 6128 308640 6180
rect 309784 6128 309836 6180
rect 376392 6128 376444 6180
rect 386328 6128 386380 6180
rect 490564 6128 490616 6180
rect 280804 4904 280856 4956
rect 188344 4836 188396 4888
rect 190828 4836 190880 4888
rect 330024 4836 330076 4888
rect 352564 4836 352616 4888
rect 358544 4836 358596 4888
rect 173716 4768 173768 4820
rect 183744 4768 183796 4820
rect 194508 4768 194560 4820
rect 212264 4768 212316 4820
rect 221464 4768 221516 4820
rect 240784 4768 240836 4820
rect 242164 4768 242216 4820
rect 255044 4768 255096 4820
rect 255964 4768 256016 4820
rect 280068 4768 280120 4820
rect 309048 4768 309100 4820
rect 378784 4768 378836 4820
rect 382188 4768 382240 4820
rect 483480 4768 483532 4820
rect 192484 4156 192536 4208
rect 194416 4156 194468 4208
rect 213184 4156 213236 4208
rect 215852 4156 215904 4208
rect 425152 4156 425204 4208
rect 426348 4156 426400 4208
rect 451280 4156 451332 4208
rect 452476 4156 452528 4208
rect 127808 4088 127860 4140
rect 134156 4088 134208 4140
rect 144460 4088 144512 4140
rect 146392 4088 146444 4140
rect 160008 4088 160060 4140
rect 163504 4088 163556 4140
rect 166908 4088 166960 4140
rect 172980 4088 173032 4140
rect 361488 4088 361540 4140
rect 453672 4088 453724 4140
rect 130200 4020 130252 4072
rect 135536 4020 135588 4072
rect 140872 4020 140924 4072
rect 143540 4020 143592 4072
rect 159916 4020 159968 4072
rect 162308 4020 162360 4072
rect 364248 4020 364300 4072
rect 457260 4020 457312 4072
rect 129004 3952 129056 4004
rect 135260 3952 135312 4004
rect 176568 3952 176620 4004
rect 186044 3952 186096 4004
rect 367008 3952 367060 4004
rect 460848 3952 460900 4004
rect 139676 3884 139728 3936
rect 142160 3884 142212 3936
rect 169576 3884 169628 3936
rect 176476 3884 176528 3936
rect 177856 3884 177908 3936
rect 188436 3884 188488 3936
rect 195888 3884 195940 3936
rect 214656 3884 214708 3936
rect 368388 3884 368440 3936
rect 464436 3884 464488 3936
rect 142068 3816 142120 3868
rect 143908 3816 143960 3868
rect 169668 3816 169720 3868
rect 177764 3816 177816 3868
rect 182088 3816 182140 3868
rect 195612 3816 195664 3868
rect 198648 3816 198700 3868
rect 218152 3816 218204 3868
rect 373908 3816 373960 3868
rect 471520 3816 471572 3868
rect 143264 3748 143316 3800
rect 144920 3748 144972 3800
rect 173808 3680 173860 3732
rect 182548 3748 182600 3800
rect 183468 3748 183520 3800
rect 196808 3748 196860 3800
rect 200028 3748 200080 3800
rect 221740 3748 221792 3800
rect 371148 3748 371200 3800
rect 467840 3748 467892 3800
rect 180708 3680 180760 3732
rect 193220 3680 193272 3732
rect 205548 3680 205600 3732
rect 228916 3680 228968 3732
rect 379428 3680 379480 3732
rect 478696 3680 478748 3732
rect 168196 3612 168248 3664
rect 174176 3612 174228 3664
rect 175188 3612 175240 3664
rect 184848 3612 184900 3664
rect 186228 3612 186280 3664
rect 200396 3612 200448 3664
rect 202788 3612 202840 3664
rect 225328 3612 225380 3664
rect 376668 3612 376720 3664
rect 475108 3612 475160 3664
rect 132592 3544 132644 3596
rect 138020 3544 138072 3596
rect 138480 3544 138532 3596
rect 142252 3544 142304 3596
rect 146852 3544 146904 3596
rect 147772 3544 147824 3596
rect 150440 3544 150492 3596
rect 151544 3544 151596 3596
rect 161388 3544 161440 3596
rect 164700 3544 164752 3596
rect 165436 3544 165488 3596
rect 170588 3544 170640 3596
rect 172336 3544 172388 3596
rect 181352 3544 181404 3596
rect 187608 3544 187660 3596
rect 203892 3544 203944 3596
rect 208308 3544 208360 3596
rect 232504 3544 232556 3596
rect 262220 3544 262272 3596
rect 263416 3544 263468 3596
rect 270500 3544 270552 3596
rect 271696 3544 271748 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 331220 3544 331272 3596
rect 332416 3544 332468 3596
rect 365720 3544 365772 3596
rect 366916 3544 366968 3596
rect 374000 3544 374052 3596
rect 375196 3544 375248 3596
rect 380808 3544 380860 3596
rect 482284 3544 482336 3596
rect 485780 3544 485832 3596
rect 486976 3544 487028 3596
rect 494152 3544 494204 3596
rect 495348 3544 495400 3596
rect 520280 3544 520332 3596
rect 521476 3544 521528 3596
rect 528560 3544 528612 3596
rect 529848 3544 529900 3596
rect 536932 3544 536984 3596
rect 538128 3544 538180 3596
rect 546500 3544 546552 3596
rect 547696 3544 547748 3596
rect 563152 3544 563204 3596
rect 564348 3544 564400 3596
rect 1676 3476 1728 3528
rect 132500 3476 132552 3528
rect 137284 3476 137336 3528
rect 140780 3476 140832 3528
rect 151820 3476 151872 3528
rect 152740 3476 152792 3528
rect 153108 3476 153160 3528
rect 153936 3476 153988 3528
rect 155776 3476 155828 3528
rect 156328 3476 156380 3528
rect 157248 3476 157300 3528
rect 158720 3476 158772 3528
rect 162768 3476 162820 3528
rect 167092 3476 167144 3528
rect 168288 3476 168340 3528
rect 175372 3476 175424 3528
rect 177948 3476 178000 3528
rect 189632 3476 189684 3528
rect 190368 3476 190420 3528
rect 201500 3476 201552 3528
rect 202696 3476 202748 3528
rect 211160 3476 211212 3528
rect 236000 3476 236052 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 252560 3476 252612 3528
rect 253848 3476 253900 3528
rect 287060 3476 287112 3528
rect 288348 3476 288400 3528
rect 296720 3476 296772 3528
rect 297916 3476 297968 3528
rect 305000 3476 305052 3528
rect 306196 3476 306248 3528
rect 313280 3476 313332 3528
rect 314568 3476 314620 3528
rect 347780 3476 347832 3528
rect 349068 3476 349120 3528
rect 356060 3476 356112 3528
rect 357348 3476 357400 3528
rect 572 3408 624 3460
rect 131120 3408 131172 3460
rect 134892 3408 134944 3460
rect 139400 3408 139452 3460
rect 154488 3408 154540 3460
rect 155132 3408 155184 3460
rect 158628 3408 158680 3460
rect 161112 3408 161164 3460
rect 161296 3408 161348 3460
rect 165896 3408 165948 3460
rect 171048 3408 171100 3460
rect 178960 3408 179012 3460
rect 179328 3408 179380 3460
rect 192024 3408 192076 3460
rect 193128 3408 193180 3460
rect 211068 3408 211120 3460
rect 212448 3408 212500 3460
rect 239588 3408 239640 3460
rect 355968 3408 356020 3460
rect 446588 3476 446640 3528
rect 448428 3476 448480 3528
rect 578608 3476 578660 3528
rect 578976 3476 579028 3528
rect 581000 3476 581052 3528
rect 358728 3408 358780 3460
rect 450176 3408 450228 3460
rect 451188 3408 451240 3460
rect 582196 3408 582248 3460
rect 136088 3340 136140 3392
rect 139492 3340 139544 3392
rect 207480 3340 207532 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 416780 3340 416832 3392
rect 417976 3340 418028 3392
rect 433340 3340 433392 3392
rect 434628 3340 434680 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 145656 3272 145708 3324
rect 146300 3272 146352 3324
rect 155868 3272 155920 3324
rect 157524 3272 157576 3324
rect 164056 3272 164108 3324
rect 168196 3272 168248 3324
rect 571340 3272 571392 3324
rect 572628 3272 572680 3324
rect 578884 3272 578936 3324
rect 579804 3272 579856 3324
rect 133788 3204 133840 3256
rect 138296 3204 138348 3256
rect 164148 3136 164200 3188
rect 169392 3136 169444 3188
rect 126612 3068 126664 3120
rect 133880 3068 133932 3120
rect 131396 3000 131448 3052
rect 136640 3000 136692 3052
rect 157156 3000 157208 3052
rect 159916 3000 159968 3052
rect 165528 3000 165580 3052
rect 171784 3000 171836 3052
rect 172428 2932 172480 2984
rect 180156 2932 180208 2984
rect 502340 2728 502392 2780
rect 503628 2728 503680 2780
rect 364340 552 364392 604
rect 364524 552 364576 604
rect 367100 552 367152 604
rect 368020 552 368072 604
rect 368480 552 368532 604
rect 369216 552 369268 604
rect 369860 552 369912 604
rect 370412 552 370464 604
rect 372620 552 372672 604
rect 372804 552 372856 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 379520 552 379572 604
rect 379980 552 380032 604
rect 499580 552 499632 604
rect 500132 552 500184 604
rect 500960 552 501012 604
rect 501236 552 501288 604
rect 503720 552 503772 604
rect 504824 552 504876 604
rect 505100 552 505152 604
rect 506020 552 506072 604
rect 506480 552 506532 604
rect 507216 552 507268 604
rect 576860 552 576912 604
rect 577412 552 577464 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3330 682272 3386 682281
rect 3330 682207 3386 682216
rect 3344 681766 3372 682207
rect 3332 681760 3384 681766
rect 3332 681702 3384 681708
rect 6184 681760 6236 681766
rect 6184 681702 6236 681708
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3238 624880 3294 624889
rect 3238 624815 3294 624824
rect 3252 623830 3280 624815
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 3238 509960 3294 509969
rect 3238 509895 3294 509904
rect 3252 509318 3280 509895
rect 3240 509312 3292 509318
rect 3240 509254 3292 509260
rect 3436 502314 3464 667927
rect 3514 610464 3570 610473
rect 3514 610399 3570 610408
rect 3424 502308 3476 502314
rect 3424 502250 3476 502256
rect 3422 495544 3478 495553
rect 3422 495479 3478 495488
rect 3436 433294 3464 495479
rect 3528 478854 3556 610399
rect 4066 567352 4122 567361
rect 4066 567287 4068 567296
rect 4120 567287 4122 567296
rect 4068 567258 4120 567264
rect 3606 553072 3662 553081
rect 3606 553007 3662 553016
rect 3516 478848 3568 478854
rect 3516 478790 3568 478796
rect 3620 455394 3648 553007
rect 3698 538656 3754 538665
rect 3698 538591 3754 538600
rect 3608 455388 3660 455394
rect 3608 455330 3660 455336
rect 3514 452432 3570 452441
rect 3514 452367 3570 452376
rect 3424 433288 3476 433294
rect 3424 433230 3476 433236
rect 3422 423736 3478 423745
rect 3422 423671 3478 423680
rect 3436 402966 3464 423671
rect 3528 418130 3556 452367
rect 3712 448526 3740 538591
rect 6196 509250 6224 681702
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 9036 652792 9088 652798
rect 9036 652734 9088 652740
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 9048 624442 9076 652734
rect 9036 624436 9088 624442
rect 9036 624378 9088 624384
rect 8944 623824 8996 623830
rect 8944 623766 8996 623772
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 589286 8064 591926
rect 8024 589280 8076 589286
rect 8024 589222 8076 589228
rect 8024 579760 8076 579766
rect 7944 579708 8024 579714
rect 7944 579702 8076 579708
rect 7944 579686 8064 579702
rect 7944 579630 7972 579686
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 8116 579624 8168 579630
rect 8116 579566 8168 579572
rect 8128 562970 8156 579566
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 8116 562964 8168 562970
rect 8116 562906 8168 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8208 543788 8260 543794
rect 8208 543730 8260 543736
rect 8220 540977 8248 543730
rect 8206 540968 8262 540977
rect 8206 540903 8262 540912
rect 8390 540968 8446 540977
rect 8390 540903 8446 540912
rect 8404 533882 8432 540903
rect 8128 533854 8432 533882
rect 8128 531321 8156 533854
rect 8114 531312 8170 531321
rect 8114 531247 8170 531256
rect 8298 531312 8354 531321
rect 8298 531247 8354 531256
rect 8312 524346 8340 531247
rect 8116 524340 8168 524346
rect 8116 524282 8168 524288
rect 8300 524340 8352 524346
rect 8300 524282 8352 524288
rect 8128 515438 8156 524282
rect 8116 515432 8168 515438
rect 8116 515374 8168 515380
rect 7564 509312 7616 509318
rect 7564 509254 7616 509260
rect 6184 509244 6236 509250
rect 6184 509186 6236 509192
rect 3790 481128 3846 481137
rect 3790 481063 3846 481072
rect 3700 448520 3752 448526
rect 3700 448462 3752 448468
rect 3606 438016 3662 438025
rect 3606 437951 3662 437960
rect 3516 418124 3568 418130
rect 3516 418066 3568 418072
rect 3620 409834 3648 437951
rect 3804 425066 3832 481063
rect 7576 440230 7604 509254
rect 8956 485790 8984 623766
rect 11704 594856 11756 594862
rect 11704 594798 11756 594804
rect 10324 567316 10376 567322
rect 10324 567258 10376 567264
rect 8944 485784 8996 485790
rect 8944 485726 8996 485732
rect 10336 463690 10364 567258
rect 11716 470558 11744 594798
rect 24780 515506 24808 699654
rect 41340 515574 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 72884 637560 72936 637566
rect 72884 637502 72936 637508
rect 72896 630578 72924 637502
rect 72896 630550 73108 630578
rect 73080 626550 73108 630550
rect 73068 626544 73120 626550
rect 73068 626486 73120 626492
rect 73068 616888 73120 616894
rect 73068 616830 73120 616836
rect 73080 611454 73108 616830
rect 73068 611448 73120 611454
rect 73068 611390 73120 611396
rect 72884 611312 72936 611318
rect 72884 611254 72936 611260
rect 72896 608546 72924 611254
rect 72974 608560 73030 608569
rect 72896 608518 72974 608546
rect 72974 608495 73030 608504
rect 73158 608560 73214 608569
rect 73158 608495 73214 608504
rect 73172 601594 73200 608495
rect 72976 601588 73028 601594
rect 72976 601530 73028 601536
rect 73160 601588 73212 601594
rect 73160 601530 73212 601536
rect 72988 598942 73016 601530
rect 72976 598936 73028 598942
rect 72976 598878 73028 598884
rect 72884 589348 72936 589354
rect 72884 589290 72936 589296
rect 72896 582418 72924 589290
rect 72700 582412 72752 582418
rect 72700 582354 72752 582360
rect 72884 582412 72936 582418
rect 72884 582354 72936 582360
rect 72712 579630 72740 582354
rect 72700 579624 72752 579630
rect 72700 579566 72752 579572
rect 72608 569968 72660 569974
rect 72608 569910 72660 569916
rect 72620 563106 72648 569910
rect 72608 563100 72660 563106
rect 72608 563042 72660 563048
rect 72700 562964 72752 562970
rect 72700 562906 72752 562912
rect 72712 560250 72740 562906
rect 72700 560244 72752 560250
rect 72700 560186 72752 560192
rect 72884 550656 72936 550662
rect 72884 550598 72936 550604
rect 72896 543658 72924 550598
rect 72700 543652 72752 543658
rect 72700 543594 72752 543600
rect 72884 543652 72936 543658
rect 72884 543594 72936 543600
rect 72712 534070 72740 543594
rect 72700 534064 72752 534070
rect 72700 534006 72752 534012
rect 72884 534064 72936 534070
rect 72884 534006 72936 534012
rect 72896 531298 72924 534006
rect 72804 531270 72924 531298
rect 72804 524482 72832 531270
rect 72792 524476 72844 524482
rect 72792 524418 72844 524424
rect 72792 521688 72844 521694
rect 72792 521630 72844 521636
rect 72804 515642 72832 521630
rect 89640 515710 89668 699654
rect 106200 515778 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 129004 624436 129056 624442
rect 129004 624378 129056 624384
rect 106188 515772 106240 515778
rect 106188 515714 106240 515720
rect 89628 515704 89680 515710
rect 89628 515646 89680 515652
rect 72792 515636 72844 515642
rect 72792 515578 72844 515584
rect 41328 515568 41380 515574
rect 41328 515510 41380 515516
rect 24768 515500 24820 515506
rect 24768 515442 24820 515448
rect 128360 509244 128412 509250
rect 128360 509186 128412 509192
rect 128372 508609 128400 509186
rect 128358 508600 128414 508609
rect 128358 508535 128414 508544
rect 128360 502308 128412 502314
rect 128360 502250 128412 502256
rect 128372 500993 128400 502250
rect 128358 500984 128414 500993
rect 128358 500919 128414 500928
rect 129016 493377 129044 624378
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 137756 596222 137784 605798
rect 154316 596222 154344 605798
rect 137744 596216 137796 596222
rect 137928 596216 137980 596222
rect 137744 596158 137796 596164
rect 137848 596164 137928 596170
rect 137848 596158 137980 596164
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 137848 596142 137968 596158
rect 154408 596142 154528 596158
rect 137848 591954 137876 596142
rect 154408 591954 154436 596142
rect 137756 591926 137876 591954
rect 154316 591926 154436 591954
rect 137756 589286 137784 591926
rect 154316 589286 154344 591926
rect 137744 589280 137796 589286
rect 137744 589222 137796 589228
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 137744 579760 137796 579766
rect 137664 579708 137744 579714
rect 154304 579760 154356 579766
rect 137664 579702 137796 579708
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 137664 579686 137784 579702
rect 154224 579686 154344 579702
rect 137664 579630 137692 579686
rect 154224 579630 154252 579686
rect 137652 579624 137704 579630
rect 137652 579566 137704 579572
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 137560 569968 137612 569974
rect 137560 569910 137612 569916
rect 137572 563106 137600 569910
rect 137560 563100 137612 563106
rect 137560 563042 137612 563048
rect 154408 562970 154436 579566
rect 137652 562964 137704 562970
rect 137652 562906 137704 562912
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 137664 560250 137692 562906
rect 137652 560244 137704 560250
rect 137652 560186 137704 560192
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 137836 550656 137888 550662
rect 137836 550598 137888 550604
rect 137848 543658 137876 550598
rect 154316 550594 154344 553302
rect 154304 550588 154356 550594
rect 154304 550530 154356 550536
rect 154488 543788 154540 543794
rect 154488 543730 154540 543736
rect 137652 543652 137704 543658
rect 137652 543594 137704 543600
rect 137836 543652 137888 543658
rect 137836 543594 137888 543600
rect 137664 534070 137692 543594
rect 154500 540977 154528 543730
rect 154210 540968 154266 540977
rect 154210 540903 154266 540912
rect 154486 540968 154542 540977
rect 154486 540903 154542 540912
rect 137652 534064 137704 534070
rect 137652 534006 137704 534012
rect 137836 534064 137888 534070
rect 137836 534006 137888 534012
rect 137848 531298 137876 534006
rect 154224 531350 154252 540903
rect 137756 531270 137876 531298
rect 154212 531344 154264 531350
rect 154212 531286 154264 531292
rect 154304 531344 154356 531350
rect 154304 531286 154356 531292
rect 137756 524482 137784 531270
rect 154316 524482 154344 531286
rect 137744 524476 137796 524482
rect 137744 524418 137796 524424
rect 154304 524476 154356 524482
rect 154304 524418 154356 524424
rect 154396 524340 154448 524346
rect 154396 524282 154448 524288
rect 137744 521688 137796 521694
rect 137744 521630 137796 521636
rect 137756 518922 137784 521630
rect 137756 518894 137968 518922
rect 137940 515522 137968 518894
rect 137940 515494 138060 515522
rect 154408 515506 154436 524282
rect 171060 515574 171088 700198
rect 196808 515772 196860 515778
rect 196808 515714 196860 515720
rect 185032 515704 185084 515710
rect 185032 515646 185084 515652
rect 173256 515636 173308 515642
rect 173256 515578 173308 515584
rect 161480 515568 161532 515574
rect 161480 515510 161532 515516
rect 171048 515568 171100 515574
rect 171048 515510 171100 515516
rect 138032 515438 138060 515494
rect 149704 515500 149756 515506
rect 149704 515442 149756 515448
rect 154396 515500 154448 515506
rect 154396 515442 154448 515448
rect 137928 515432 137980 515438
rect 137928 515374 137980 515380
rect 138020 515432 138072 515438
rect 138020 515374 138072 515380
rect 137940 512380 137968 515374
rect 149716 512380 149744 515442
rect 161492 512380 161520 515510
rect 173268 512380 173296 515578
rect 185044 512380 185072 515646
rect 196820 512380 196848 515714
rect 202800 515642 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 218992 579630 219020 582354
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 218992 560250 219020 562906
rect 218980 560244 219032 560250
rect 218980 560186 219032 560192
rect 219164 550656 219216 550662
rect 219164 550598 219216 550604
rect 219176 543658 219204 550598
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 219164 543652 219216 543658
rect 219164 543594 219216 543600
rect 218992 534070 219020 543594
rect 218980 534064 219032 534070
rect 218980 534006 219032 534012
rect 219164 534064 219216 534070
rect 219164 534006 219216 534012
rect 219176 531298 219204 534006
rect 219084 531270 219204 531298
rect 219084 524482 219112 531270
rect 219072 524476 219124 524482
rect 219072 524418 219124 524424
rect 219072 521688 219124 521694
rect 219072 521630 219124 521636
rect 202788 515636 202840 515642
rect 202788 515578 202840 515584
rect 219084 515438 219112 521630
rect 232228 515568 232280 515574
rect 232228 515510 232280 515516
rect 220452 515500 220504 515506
rect 220452 515442 220504 515448
rect 208584 515432 208636 515438
rect 208584 515374 208636 515380
rect 219072 515432 219124 515438
rect 219072 515374 219124 515380
rect 208596 512380 208624 515374
rect 220464 512380 220492 515442
rect 232240 512380 232268 515510
rect 235920 515506 235948 699654
rect 244004 515636 244056 515642
rect 244004 515578 244056 515584
rect 235908 515500 235960 515506
rect 235908 515442 235960 515448
rect 244016 512380 244044 515578
rect 267556 515500 267608 515506
rect 267556 515442 267608 515448
rect 255780 515432 255832 515438
rect 255780 515374 255832 515380
rect 255792 512380 255820 515374
rect 267568 512380 267596 515442
rect 267660 515438 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654158 284064 663734
rect 284024 654152 284076 654158
rect 284024 654094 284076 654100
rect 284208 654152 284260 654158
rect 284208 654094 284260 654100
rect 284220 644450 284248 654094
rect 284036 644422 284248 644450
rect 284036 634846 284064 644422
rect 284024 634840 284076 634846
rect 284024 634782 284076 634788
rect 284208 634840 284260 634846
rect 284208 634782 284260 634788
rect 284220 625138 284248 634782
rect 284036 625110 284248 625138
rect 284036 615534 284064 625110
rect 284024 615528 284076 615534
rect 284024 615470 284076 615476
rect 284208 615528 284260 615534
rect 284208 615470 284260 615476
rect 284220 605826 284248 615470
rect 284036 605798 284248 605826
rect 284036 596222 284064 605798
rect 284024 596216 284076 596222
rect 284208 596216 284260 596222
rect 284024 596158 284076 596164
rect 284128 596164 284208 596170
rect 284128 596158 284260 596164
rect 284128 596142 284248 596158
rect 284128 591954 284156 596142
rect 284036 591926 284156 591954
rect 284036 589286 284064 591926
rect 284024 589280 284076 589286
rect 284024 589222 284076 589228
rect 284024 579760 284076 579766
rect 283944 579708 284024 579714
rect 283944 579702 284076 579708
rect 283944 579686 284064 579702
rect 283944 579630 283972 579686
rect 283932 579624 283984 579630
rect 283932 579566 283984 579572
rect 284116 579624 284168 579630
rect 284116 579566 284168 579572
rect 284128 562970 284156 579566
rect 283932 562964 283984 562970
rect 283932 562906 283984 562912
rect 284116 562964 284168 562970
rect 284116 562906 284168 562912
rect 283944 553330 283972 562906
rect 283944 553302 284064 553330
rect 284036 550594 284064 553302
rect 284024 550588 284076 550594
rect 284024 550530 284076 550536
rect 284208 543788 284260 543794
rect 284208 543730 284260 543736
rect 284220 540977 284248 543730
rect 284206 540968 284262 540977
rect 284206 540903 284262 540912
rect 284390 540968 284446 540977
rect 284390 540903 284446 540912
rect 284404 533882 284432 540903
rect 284128 533854 284432 533882
rect 284128 531321 284156 533854
rect 284114 531312 284170 531321
rect 284114 531247 284170 531256
rect 284298 531312 284354 531321
rect 284298 531247 284354 531256
rect 284312 524346 284340 531247
rect 284116 524340 284168 524346
rect 284116 524282 284168 524288
rect 284300 524340 284352 524346
rect 284300 524282 284352 524288
rect 284128 516118 284156 524282
rect 284116 516112 284168 516118
rect 284116 516054 284168 516060
rect 291108 516112 291160 516118
rect 291108 516054 291160 516060
rect 267648 515432 267700 515438
rect 267648 515374 267700 515380
rect 279332 515432 279384 515438
rect 279332 515374 279384 515380
rect 279344 512380 279372 515374
rect 291120 512380 291148 516054
rect 300780 514894 300808 699654
rect 332520 697610 332548 703520
rect 348804 703474 348832 703520
rect 364996 703474 365024 703520
rect 348804 703446 348924 703474
rect 364996 703446 365116 703474
rect 331220 697604 331272 697610
rect 331220 697546 331272 697552
rect 332508 697604 332560 697610
rect 332508 697546 332560 697552
rect 326528 515500 326580 515506
rect 326528 515442 326580 515448
rect 314752 515432 314804 515438
rect 314752 515374 314804 515380
rect 300768 514888 300820 514894
rect 300768 514830 300820 514836
rect 302976 514888 303028 514894
rect 302976 514830 303028 514836
rect 302988 512380 303016 514830
rect 314764 512380 314792 515374
rect 326540 512380 326568 515442
rect 331232 515438 331260 697546
rect 348896 692850 348924 703446
rect 365088 692850 365116 703446
rect 347780 692844 347832 692850
rect 347780 692786 347832 692792
rect 348884 692844 348936 692850
rect 348884 692786 348936 692792
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 347792 683074 347820 692786
rect 364352 683074 364380 692786
rect 347792 683046 348004 683074
rect 364352 683046 364564 683074
rect 347976 673538 348004 683046
rect 364536 673538 364564 683046
rect 347780 673532 347832 673538
rect 347780 673474 347832 673480
rect 347964 673532 348016 673538
rect 347964 673474 348016 673480
rect 364340 673532 364392 673538
rect 364340 673474 364392 673480
rect 364524 673532 364576 673538
rect 364524 673474 364576 673480
rect 347792 663762 347820 673474
rect 364352 663762 364380 673474
rect 347792 663734 348004 663762
rect 364352 663734 364564 663762
rect 347976 654158 348004 663734
rect 364536 654158 364564 663734
rect 347780 654152 347832 654158
rect 347780 654094 347832 654100
rect 347964 654152 348016 654158
rect 347964 654094 348016 654100
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 347792 644450 347820 654094
rect 364352 644450 364380 654094
rect 347792 644422 348004 644450
rect 364352 644422 364564 644450
rect 347976 634846 348004 644422
rect 364536 634846 364564 644422
rect 347780 634840 347832 634846
rect 347780 634782 347832 634788
rect 347964 634840 348016 634846
rect 347964 634782 348016 634788
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 347792 625138 347820 634782
rect 364352 625138 364380 634782
rect 347792 625110 348004 625138
rect 364352 625110 364564 625138
rect 347976 615534 348004 625110
rect 364536 615534 364564 625110
rect 347780 615528 347832 615534
rect 347780 615470 347832 615476
rect 347964 615528 348016 615534
rect 347964 615470 348016 615476
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 347792 605826 347820 615470
rect 364352 605826 364380 615470
rect 347792 605798 348004 605826
rect 364352 605798 364564 605826
rect 347976 596222 348004 605798
rect 364536 596222 364564 605798
rect 347780 596216 347832 596222
rect 347964 596216 348016 596222
rect 347832 596164 347912 596170
rect 347780 596158 347912 596164
rect 347964 596158 348016 596164
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 347792 596142 347912 596158
rect 364352 596142 364472 596158
rect 347884 596034 347912 596142
rect 364444 596034 364472 596142
rect 347884 596006 348004 596034
rect 364444 596006 364564 596034
rect 347976 591954 348004 596006
rect 364536 591954 364564 596006
rect 347884 591926 348004 591954
rect 364444 591926 364564 591954
rect 347884 589286 347912 591926
rect 364444 589286 364472 591926
rect 347872 589280 347924 589286
rect 347872 589222 347924 589228
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 347780 579692 347832 579698
rect 347780 579634 347832 579640
rect 364340 579692 364392 579698
rect 364340 579634 364392 579640
rect 347792 572642 347820 579634
rect 364352 572642 364380 579634
rect 347792 572614 347912 572642
rect 364352 572614 364472 572642
rect 347884 569906 347912 572614
rect 364444 569906 364472 572614
rect 347872 569900 347924 569906
rect 347872 569842 347924 569848
rect 364432 569900 364484 569906
rect 364432 569842 364484 569848
rect 348056 563100 348108 563106
rect 348056 563042 348108 563048
rect 364616 563100 364668 563106
rect 364616 563042 364668 563048
rect 348068 560289 348096 563042
rect 364628 560289 364656 563042
rect 347870 560280 347926 560289
rect 347870 560215 347926 560224
rect 348054 560280 348110 560289
rect 348054 560215 348110 560224
rect 364430 560280 364486 560289
rect 364430 560215 364486 560224
rect 364614 560280 364670 560289
rect 364614 560215 364670 560224
rect 347884 550662 347912 560215
rect 364444 550662 364472 560215
rect 347872 550656 347924 550662
rect 347872 550598 347924 550604
rect 348148 550656 348200 550662
rect 348148 550598 348200 550604
rect 364432 550656 364484 550662
rect 364432 550598 364484 550604
rect 364708 550656 364760 550662
rect 364708 550598 364760 550604
rect 348160 543862 348188 550598
rect 364720 543862 364748 550598
rect 348148 543856 348200 543862
rect 348148 543798 348200 543804
rect 364708 543856 364760 543862
rect 364708 543798 364760 543804
rect 348056 543720 348108 543726
rect 348056 543662 348108 543668
rect 364616 543720 364668 543726
rect 364616 543662 364668 543668
rect 348068 540977 348096 543662
rect 364628 540977 364656 543662
rect 347870 540968 347926 540977
rect 347870 540903 347926 540912
rect 348054 540968 348110 540977
rect 348054 540903 348110 540912
rect 364430 540968 364486 540977
rect 364430 540903 364486 540912
rect 364614 540968 364670 540977
rect 364614 540903 364670 540912
rect 347884 531350 347912 540903
rect 364444 531350 364472 540903
rect 347872 531344 347924 531350
rect 347872 531286 347924 531292
rect 348148 531344 348200 531350
rect 348148 531286 348200 531292
rect 364432 531344 364484 531350
rect 364432 531286 364484 531292
rect 364708 531344 364760 531350
rect 364708 531286 364760 531292
rect 348160 521694 348188 531286
rect 364720 521694 364748 531286
rect 347964 521688 348016 521694
rect 347964 521630 348016 521636
rect 348148 521688 348200 521694
rect 348148 521630 348200 521636
rect 364524 521688 364576 521694
rect 364524 521630 364576 521636
rect 364708 521688 364760 521694
rect 364708 521630 364760 521636
rect 347976 515506 348004 521630
rect 350080 515568 350132 515574
rect 350080 515510 350132 515516
rect 347964 515500 348016 515506
rect 347964 515442 348016 515448
rect 331220 515432 331272 515438
rect 331220 515374 331272 515380
rect 338304 515432 338356 515438
rect 338304 515374 338356 515380
rect 338316 512380 338344 515374
rect 350092 512380 350120 515510
rect 361856 515500 361908 515506
rect 361856 515442 361908 515448
rect 361868 512380 361896 515442
rect 364536 515438 364564 521630
rect 385500 515772 385552 515778
rect 385500 515714 385552 515720
rect 364524 515432 364576 515438
rect 364524 515374 364576 515380
rect 373632 515432 373684 515438
rect 373632 515374 373684 515380
rect 373644 512380 373672 515374
rect 385512 512380 385540 515714
rect 397276 515704 397328 515710
rect 397276 515646 397328 515652
rect 397288 512380 397316 515646
rect 397472 515574 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 413756 698290 413784 703446
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 429856 684486 429884 703520
rect 429200 684480 429252 684486
rect 429200 684422 429252 684428
rect 429844 684480 429896 684486
rect 429844 684422 429896 684428
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 429212 683126 429240 684422
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 429200 683120 429252 683126
rect 429200 683062 429252 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 413112 659682 413140 666538
rect 429672 659682 429700 666538
rect 412928 659654 413140 659682
rect 429488 659654 429700 659682
rect 412928 647290 412956 659654
rect 429488 647290 429516 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 412836 640422 412864 647226
rect 429396 640422 429424 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 412928 630698 412956 640358
rect 429488 630698 429516 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 412744 630578 412772 630634
rect 429304 630578 429332 630634
rect 412744 630550 412864 630578
rect 429304 630550 429424 630578
rect 412836 621058 412864 630550
rect 429396 621058 429424 630550
rect 412836 621030 412956 621058
rect 429396 621030 429516 621058
rect 412928 611386 412956 621030
rect 429488 611386 429516 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 412744 611266 412772 611322
rect 429304 611266 429332 611322
rect 412744 611238 412864 611266
rect 429304 611238 429424 611266
rect 412836 608598 412864 611238
rect 429396 608598 429424 611238
rect 412824 608592 412876 608598
rect 412824 608534 412876 608540
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 413008 601724 413060 601730
rect 413008 601666 413060 601672
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 413020 598942 413048 601666
rect 429580 598942 429608 601666
rect 413008 598936 413060 598942
rect 413008 598878 413060 598884
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 413100 589348 413152 589354
rect 413100 589290 413152 589296
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 413112 582486 413140 589290
rect 429672 582486 429700 589290
rect 413100 582480 413152 582486
rect 413100 582422 413152 582428
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 413008 582344 413060 582350
rect 413008 582286 413060 582292
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 413020 572642 413048 582286
rect 429580 572642 429608 582286
rect 412836 572614 413048 572642
rect 429396 572614 429608 572642
rect 412836 569922 412864 572614
rect 429396 569922 429424 572614
rect 412744 569894 412864 569922
rect 429304 569894 429424 569922
rect 412744 563174 412772 569894
rect 429304 563174 429332 569894
rect 412732 563168 412784 563174
rect 412732 563110 412784 563116
rect 429292 563168 429344 563174
rect 429292 563110 429344 563116
rect 412732 563032 412784 563038
rect 412732 562974 412784 562980
rect 429292 563032 429344 563038
rect 429292 562974 429344 562980
rect 412744 560250 412772 562974
rect 429304 560250 429332 562974
rect 412732 560244 412784 560250
rect 412732 560186 412784 560192
rect 429292 560244 429344 560250
rect 429292 560186 429344 560192
rect 412916 550656 412968 550662
rect 412916 550598 412968 550604
rect 429476 550656 429528 550662
rect 429476 550598 429528 550604
rect 412928 543658 412956 550598
rect 429488 543658 429516 550598
rect 412732 543652 412784 543658
rect 412732 543594 412784 543600
rect 412916 543652 412968 543658
rect 412916 543594 412968 543600
rect 429292 543652 429344 543658
rect 429292 543594 429344 543600
rect 429476 543652 429528 543658
rect 429476 543594 429528 543600
rect 412744 534018 412772 543594
rect 429304 534018 429332 543594
rect 412744 533990 412864 534018
rect 429304 533990 429424 534018
rect 412836 524498 412864 533990
rect 429396 524498 429424 533990
rect 412836 524470 412956 524498
rect 429396 524470 429516 524498
rect 409052 515636 409104 515642
rect 409052 515578 409104 515584
rect 397460 515568 397512 515574
rect 397460 515510 397512 515516
rect 409064 512380 409092 515578
rect 412928 515506 412956 524470
rect 420828 515568 420880 515574
rect 420828 515510 420880 515516
rect 412916 515500 412968 515506
rect 412916 515442 412968 515448
rect 420840 512380 420868 515510
rect 429488 515438 429516 524470
rect 462332 515778 462360 703520
rect 478524 703474 478552 703520
rect 494808 703474 494836 703520
rect 478524 703446 478644 703474
rect 494808 703446 494928 703474
rect 476764 696992 476816 696998
rect 476764 696934 476816 696940
rect 475384 650072 475436 650078
rect 475384 650014 475436 650020
rect 471244 603152 471296 603158
rect 471244 603094 471296 603100
rect 467104 556232 467156 556238
rect 467104 556174 467156 556180
rect 462320 515772 462372 515778
rect 462320 515714 462372 515720
rect 432604 515500 432656 515506
rect 432604 515442 432656 515448
rect 429476 515432 429528 515438
rect 429476 515374 429528 515380
rect 432616 512380 432644 515442
rect 444380 515432 444432 515438
rect 444380 515374 444432 515380
rect 444392 512380 444420 515374
rect 462964 509312 463016 509318
rect 462964 509254 463016 509260
rect 453212 509244 453264 509250
rect 453212 509186 453264 509192
rect 453224 508881 453252 509186
rect 453210 508872 453266 508881
rect 453210 508807 453266 508816
rect 453396 502308 453448 502314
rect 453396 502250 453448 502256
rect 453408 501809 453436 502250
rect 453394 501800 453450 501809
rect 453394 501735 453450 501744
rect 460204 498228 460256 498234
rect 460204 498170 460256 498176
rect 453948 495440 454000 495446
rect 453948 495382 454000 495388
rect 453960 494601 453988 495382
rect 453946 494592 454002 494601
rect 453946 494527 454002 494536
rect 129002 493368 129058 493377
rect 129002 493303 129058 493312
rect 453764 488504 453816 488510
rect 453764 488446 453816 488452
rect 453776 487529 453804 488446
rect 453762 487520 453818 487529
rect 453762 487455 453818 487464
rect 456064 485852 456116 485858
rect 456064 485794 456116 485800
rect 128360 485784 128412 485790
rect 128358 485752 128360 485761
rect 128412 485752 128414 485761
rect 128358 485687 128414 485696
rect 453764 481636 453816 481642
rect 453764 481578 453816 481584
rect 453776 480457 453804 481578
rect 453762 480448 453818 480457
rect 453762 480383 453818 480392
rect 128360 478848 128412 478854
rect 128360 478790 128412 478796
rect 128372 478145 128400 478790
rect 128358 478136 128414 478145
rect 128358 478071 128414 478080
rect 453948 473340 454000 473346
rect 453948 473282 454000 473288
rect 453960 473249 453988 473282
rect 453946 473240 454002 473249
rect 453946 473175 454002 473184
rect 11704 470552 11756 470558
rect 128360 470552 128412 470558
rect 11704 470494 11756 470500
rect 128358 470520 128360 470529
rect 128412 470520 128414 470529
rect 128358 470455 128414 470464
rect 452752 466404 452804 466410
rect 452752 466346 452804 466352
rect 452764 466177 452792 466346
rect 452750 466168 452806 466177
rect 452750 466103 452806 466112
rect 10324 463684 10376 463690
rect 10324 463626 10376 463632
rect 128360 463684 128412 463690
rect 128360 463626 128412 463632
rect 128372 462913 128400 463626
rect 128358 462904 128414 462913
rect 128358 462839 128414 462848
rect 453396 459536 453448 459542
rect 453396 459478 453448 459484
rect 453408 459105 453436 459478
rect 453394 459096 453450 459105
rect 453394 459031 453450 459040
rect 128360 455388 128412 455394
rect 128360 455330 128412 455336
rect 128372 455297 128400 455330
rect 128358 455288 128414 455297
rect 128358 455223 128414 455232
rect 453948 452600 454000 452606
rect 453948 452542 454000 452548
rect 453960 451897 453988 452542
rect 453946 451888 454002 451897
rect 453946 451823 454002 451832
rect 128360 448520 128412 448526
rect 128360 448462 128412 448468
rect 128372 447681 128400 448462
rect 128358 447672 128414 447681
rect 128358 447607 128414 447616
rect 453672 445732 453724 445738
rect 453672 445674 453724 445680
rect 453684 444825 453712 445674
rect 453670 444816 453726 444825
rect 453670 444751 453726 444760
rect 7564 440224 7616 440230
rect 7564 440166 7616 440172
rect 128360 440224 128412 440230
rect 128360 440166 128412 440172
rect 128372 440065 128400 440166
rect 128358 440056 128414 440065
rect 128358 439991 128414 440000
rect 453304 438932 453356 438938
rect 453304 438874 453356 438880
rect 128360 433288 128412 433294
rect 128360 433230 128412 433236
rect 128372 432313 128400 433230
rect 128358 432304 128414 432313
rect 128358 432239 128414 432248
rect 3792 425060 3844 425066
rect 3792 425002 3844 425008
rect 128360 425060 128412 425066
rect 128360 425002 128412 425008
rect 128372 424697 128400 425002
rect 128358 424688 128414 424697
rect 128358 424623 128414 424632
rect 128360 418124 128412 418130
rect 128360 418066 128412 418072
rect 128372 417081 128400 418066
rect 128358 417072 128414 417081
rect 128358 417007 128414 417016
rect 3608 409828 3660 409834
rect 3608 409770 3660 409776
rect 128360 409828 128412 409834
rect 128360 409770 128412 409776
rect 128372 409465 128400 409770
rect 128358 409456 128414 409465
rect 128358 409391 128414 409400
rect 3424 402960 3476 402966
rect 3424 402902 3476 402908
rect 128360 402960 128412 402966
rect 128360 402902 128412 402908
rect 128372 401849 128400 402902
rect 128358 401840 128414 401849
rect 128358 401775 128414 401784
rect 3422 395040 3478 395049
rect 3422 394975 3478 394984
rect 3436 394670 3464 394975
rect 3424 394664 3476 394670
rect 3424 394606 3476 394612
rect 128360 394664 128412 394670
rect 128360 394606 128412 394612
rect 128372 394233 128400 394606
rect 128358 394224 128414 394233
rect 128358 394159 128414 394168
rect 453316 387841 453344 438874
rect 453764 438864 453816 438870
rect 453764 438806 453816 438812
rect 453776 437753 453804 438806
rect 453762 437744 453818 437753
rect 453762 437679 453818 437688
rect 453948 430568 454000 430574
rect 453946 430536 453948 430545
rect 454000 430536 454002 430545
rect 453946 430471 454002 430480
rect 453948 423632 454000 423638
rect 453948 423574 454000 423580
rect 453960 423473 453988 423574
rect 453946 423464 454002 423473
rect 453946 423399 454002 423408
rect 453948 416424 454000 416430
rect 453946 416392 453948 416401
rect 454000 416392 454002 416401
rect 453946 416327 454002 416336
rect 456076 409426 456104 485794
rect 460216 416430 460244 498170
rect 462976 423638 463004 509254
rect 467116 445738 467144 556174
rect 471256 466410 471284 603094
rect 475396 488510 475424 650014
rect 476776 509250 476804 696934
rect 478616 692850 478644 703446
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 477512 683074 477540 692786
rect 494900 685914 494928 703446
rect 494244 685908 494296 685914
rect 494244 685850 494296 685856
rect 494888 685908 494940 685914
rect 494888 685850 494940 685856
rect 477512 683046 477724 683074
rect 477696 673538 477724 683046
rect 494256 678994 494284 685850
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 483664 673532 483716 673538
rect 483664 673474 483716 673480
rect 477512 663762 477540 673474
rect 477512 663734 477724 663762
rect 477696 654158 477724 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 477512 644450 477540 654094
rect 477512 644422 477724 644450
rect 477696 634846 477724 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 477512 625138 477540 634782
rect 479524 626612 479576 626618
rect 479524 626554 479576 626560
rect 477512 625110 477724 625138
rect 477696 615534 477724 625110
rect 477500 615528 477552 615534
rect 477500 615470 477552 615476
rect 477684 615528 477736 615534
rect 477684 615470 477736 615476
rect 477512 605826 477540 615470
rect 477512 605798 477724 605826
rect 477696 596222 477724 605798
rect 477500 596216 477552 596222
rect 477684 596216 477736 596222
rect 477552 596164 477632 596170
rect 477500 596158 477632 596164
rect 477684 596158 477736 596164
rect 477512 596142 477632 596158
rect 477604 596034 477632 596142
rect 477604 596006 477724 596034
rect 477696 591954 477724 596006
rect 477604 591926 477724 591954
rect 477604 589286 477632 591926
rect 477592 589280 477644 589286
rect 477592 589222 477644 589228
rect 477500 579692 477552 579698
rect 477500 579634 477552 579640
rect 477512 572642 477540 579634
rect 477512 572614 477632 572642
rect 477604 569906 477632 572614
rect 477592 569900 477644 569906
rect 477592 569842 477644 569848
rect 477776 563100 477828 563106
rect 477776 563042 477828 563048
rect 477788 560289 477816 563042
rect 477590 560280 477646 560289
rect 477590 560215 477646 560224
rect 477774 560280 477830 560289
rect 477774 560215 477830 560224
rect 477604 550662 477632 560215
rect 477592 550656 477644 550662
rect 477592 550598 477644 550604
rect 477868 550656 477920 550662
rect 477868 550598 477920 550604
rect 477880 543862 477908 550598
rect 477868 543856 477920 543862
rect 477868 543798 477920 543804
rect 477776 543720 477828 543726
rect 477776 543662 477828 543668
rect 477788 540977 477816 543662
rect 477590 540968 477646 540977
rect 477590 540903 477646 540912
rect 477774 540968 477830 540977
rect 477774 540903 477830 540912
rect 477604 531350 477632 540903
rect 477592 531344 477644 531350
rect 477592 531286 477644 531292
rect 477868 531344 477920 531350
rect 477868 531286 477920 531292
rect 477880 521694 477908 531286
rect 477684 521688 477736 521694
rect 477684 521630 477736 521636
rect 477868 521688 477920 521694
rect 477868 521630 477920 521636
rect 477696 515710 477724 521630
rect 477684 515704 477736 515710
rect 477684 515646 477736 515652
rect 476764 509244 476816 509250
rect 476764 509186 476816 509192
rect 475384 488504 475436 488510
rect 475384 488446 475436 488452
rect 479536 473346 479564 626554
rect 482284 592068 482336 592074
rect 482284 592010 482336 592016
rect 480904 545148 480956 545154
rect 480904 545090 480956 545096
rect 479524 473340 479576 473346
rect 479524 473282 479576 473288
rect 471244 466404 471296 466410
rect 471244 466346 471296 466352
rect 467104 445732 467156 445738
rect 467104 445674 467156 445680
rect 480916 438870 480944 545090
rect 482296 459542 482324 592010
rect 483676 495446 483704 673474
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 494164 659682 494192 666538
rect 494164 659654 494284 659682
rect 494256 654158 494284 659654
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 494072 644450 494100 654094
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 494072 625110 494284 625138
rect 494256 615534 494284 625110
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 494072 605826 494100 615470
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579737 493916 589222
rect 493874 579728 493930 579737
rect 489184 579692 489236 579698
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 489184 579634 489236 579640
rect 485044 532772 485096 532778
rect 485044 532714 485096 532720
rect 483664 495440 483716 495446
rect 483664 495382 483716 495388
rect 482284 459536 482336 459542
rect 482284 459478 482336 459484
rect 480904 438864 480956 438870
rect 480904 438806 480956 438812
rect 485056 430574 485084 532714
rect 489196 452606 489224 579634
rect 494072 572642 494100 579663
rect 494072 572614 494192 572642
rect 494164 569906 494192 572614
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 494348 560289 494376 563042
rect 494150 560280 494206 560289
rect 494150 560215 494206 560224
rect 494334 560280 494390 560289
rect 494334 560215 494390 560224
rect 494164 550662 494192 560215
rect 494152 550656 494204 550662
rect 494152 550598 494204 550604
rect 494428 550656 494480 550662
rect 494428 550598 494480 550604
rect 494440 543862 494468 550598
rect 494428 543856 494480 543862
rect 494428 543798 494480 543804
rect 494336 543720 494388 543726
rect 494336 543662 494388 543668
rect 494348 540977 494376 543662
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 494164 531350 494192 540903
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 494440 521694 494468 531286
rect 494244 521688 494296 521694
rect 494244 521630 494296 521636
rect 494428 521688 494480 521694
rect 494428 521630 494480 521636
rect 494256 515642 494284 521630
rect 494244 515636 494296 515642
rect 494244 515578 494296 515584
rect 527192 515574 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 694142 542768 698226
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 692782 542584 694078
rect 542544 692776 542596 692782
rect 542544 692718 542596 692724
rect 542728 692776 542780 692782
rect 542728 692718 542780 692724
rect 542740 683233 542768 692718
rect 559668 684486 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 558920 684480 558972 684486
rect 558920 684422 558972 684428
rect 559656 684480 559708 684486
rect 559656 684422 559708 684428
rect 542358 683224 542414 683233
rect 542358 683159 542414 683168
rect 542726 683224 542782 683233
rect 542726 683159 542782 683168
rect 542372 683126 542400 683159
rect 558932 683126 558960 684422
rect 542360 683120 542412 683126
rect 542360 683062 542412 683068
rect 558920 683120 558972 683126
rect 558920 683062 558972 683068
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 542832 659682 542860 666538
rect 559392 659682 559420 666538
rect 542648 659654 542860 659682
rect 559208 659654 559420 659682
rect 542648 647290 542676 659654
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 542556 640422 542584 647226
rect 559116 640422 559144 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 542648 630698 542676 640358
rect 559208 630698 559236 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 542464 630578 542492 630634
rect 559024 630578 559052 630634
rect 542464 630550 542584 630578
rect 559024 630550 559144 630578
rect 542556 621058 542584 630550
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 559116 621030 559236 621058
rect 542648 611386 542676 621030
rect 559208 611386 559236 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 542464 611266 542492 611322
rect 559024 611266 559052 611322
rect 542464 611238 542584 611266
rect 559024 611238 559144 611266
rect 542556 608598 542584 611238
rect 559116 608598 559144 611238
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 542740 598942 542768 601666
rect 559300 598942 559328 601666
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 579894 592512 579950 592521
rect 579894 592447 579950 592456
rect 579908 592074 579936 592447
rect 579896 592068 579948 592074
rect 579896 592010 579948 592016
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 542832 582486 542860 589290
rect 559392 582486 559420 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 542740 572642 542768 582286
rect 559300 572642 559328 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 542556 572614 542768 572642
rect 559116 572614 559328 572642
rect 542556 569922 542584 572614
rect 559116 569922 559144 572614
rect 542464 569894 542584 569922
rect 559024 569894 559144 569922
rect 542464 563174 542492 569894
rect 559024 563174 559052 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 542464 560250 542492 562974
rect 559024 560250 559052 562974
rect 542452 560244 542504 560250
rect 542452 560186 542504 560192
rect 559012 560244 559064 560250
rect 559012 560186 559064 560192
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 542636 550656 542688 550662
rect 542636 550598 542688 550604
rect 559196 550656 559248 550662
rect 559196 550598 559248 550604
rect 542648 543658 542676 550598
rect 559208 543658 559236 550598
rect 579894 545592 579950 545601
rect 579894 545527 579950 545536
rect 579908 545154 579936 545527
rect 579896 545148 579948 545154
rect 579896 545090 579948 545096
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542636 543652 542688 543658
rect 542636 543594 542688 543600
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559196 543652 559248 543658
rect 559196 543594 559248 543600
rect 542464 534018 542492 543594
rect 559024 534018 559052 543594
rect 542464 533990 542584 534018
rect 559024 533990 559144 534018
rect 542556 524498 542584 533990
rect 559116 524498 559144 533990
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 542556 524470 542676 524498
rect 559116 524470 559236 524498
rect 527180 515568 527232 515574
rect 527180 515510 527232 515516
rect 542648 515506 542676 524470
rect 542636 515500 542688 515506
rect 542636 515442 542688 515448
rect 559208 515438 559236 524470
rect 559196 515432 559248 515438
rect 559196 515374 559248 515380
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580276 502314 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580264 502308 580316 502314
rect 580264 502250 580316 502256
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580368 481642 580396 639367
rect 580356 481636 580408 481642
rect 580356 481578 580408 481584
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 543004 462392 543056 462398
rect 543004 462334 543056 462340
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 489184 452600 489236 452606
rect 489184 452542 489236 452548
rect 485044 430568 485096 430574
rect 485044 430510 485096 430516
rect 462964 423632 463016 423638
rect 462964 423574 463016 423580
rect 460204 416424 460256 416430
rect 460204 416366 460256 416372
rect 453396 409420 453448 409426
rect 453396 409362 453448 409368
rect 456064 409420 456116 409426
rect 456064 409362 456116 409368
rect 453408 409193 453436 409362
rect 453394 409184 453450 409193
rect 453394 409119 453450 409128
rect 543016 402966 543044 462334
rect 580262 451752 580318 451761
rect 580262 451687 580318 451696
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 579908 438938 579936 439855
rect 579896 438932 579948 438938
rect 579896 438874 579948 438880
rect 578882 416528 578938 416537
rect 578882 416463 578938 416472
rect 453948 402960 454000 402966
rect 453948 402902 454000 402908
rect 543004 402960 543056 402966
rect 543004 402902 543056 402908
rect 453960 402121 453988 402902
rect 453946 402112 454002 402121
rect 453946 402047 454002 402056
rect 453764 396024 453816 396030
rect 453764 395966 453816 395972
rect 453776 394913 453804 395966
rect 453762 394904 453818 394913
rect 453762 394839 453818 394848
rect 460204 392012 460256 392018
rect 460204 391954 460256 391960
rect 453302 387832 453358 387841
rect 453302 387767 453358 387776
rect 129002 386608 129058 386617
rect 129002 386543 129058 386552
rect 129016 380866 129044 386543
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 129004 380860 129056 380866
rect 129004 380802 129056 380808
rect 453948 380860 454000 380866
rect 453948 380802 454000 380808
rect 3252 380633 3280 380802
rect 453960 380769 453988 380802
rect 453946 380760 454002 380769
rect 453946 380695 454002 380704
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 129002 378992 129058 379001
rect 129002 378927 129058 378936
rect 129016 367062 129044 378927
rect 453396 373992 453448 373998
rect 453396 373934 453448 373940
rect 453408 373561 453436 373934
rect 453394 373552 453450 373561
rect 453394 373487 453450 373496
rect 129278 371376 129334 371385
rect 129278 371311 129334 371320
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 129004 367056 129056 367062
rect 129004 366998 129056 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 129002 363760 129058 363769
rect 129002 363695 129058 363704
rect 128358 348392 128414 348401
rect 128358 348327 128414 348336
rect 128372 347818 128400 348327
rect 3424 347812 3476 347818
rect 3424 347754 3476 347760
rect 128360 347812 128412 347818
rect 128360 347754 128412 347760
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3436 294409 3464 347754
rect 3516 338088 3568 338094
rect 3516 338030 3568 338036
rect 3528 337521 3556 338030
rect 3514 337512 3570 337521
rect 3514 337447 3570 337456
rect 128358 333160 128414 333169
rect 128358 333095 128414 333104
rect 128372 332654 128400 333095
rect 8944 332648 8996 332654
rect 8944 332590 8996 332596
rect 128360 332648 128412 332654
rect 128360 332590 128412 332596
rect 7564 324352 7616 324358
rect 7564 324294 7616 324300
rect 3516 324284 3568 324290
rect 3516 324226 3568 324232
rect 3528 323105 3556 324226
rect 3514 323096 3570 323105
rect 3514 323031 3570 323040
rect 6184 302252 6236 302258
rect 6184 302194 6236 302200
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 3424 278044 3476 278050
rect 3424 277986 3476 277992
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3148 208208 3200 208214
rect 3146 208176 3148 208185
rect 3200 208176 3202 208185
rect 3146 208111 3202 208120
rect 2872 194540 2924 194546
rect 2872 194482 2924 194488
rect 2884 193905 2912 194482
rect 2870 193896 2926 193905
rect 2870 193831 2926 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3436 165073 3464 277986
rect 3516 266076 3568 266082
rect 3516 266018 3568 266024
rect 3528 265713 3556 266018
rect 3514 265704 3570 265713
rect 3514 265639 3570 265648
rect 3516 251660 3568 251666
rect 3516 251602 3568 251608
rect 3528 251297 3556 251602
rect 3514 251288 3570 251297
rect 3514 251223 3570 251232
rect 3516 237380 3568 237386
rect 3516 237322 3568 237328
rect 3528 237017 3556 237322
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 6196 208214 6224 302194
rect 7576 251666 7604 324294
rect 8956 266082 8984 332590
rect 128358 325544 128414 325553
rect 128358 325479 128414 325488
rect 128372 324358 128400 325479
rect 128360 324352 128412 324358
rect 128360 324294 128412 324300
rect 129016 324290 129044 363695
rect 129186 356144 129242 356153
rect 129186 356079 129242 356088
rect 129094 340776 129150 340785
rect 129094 340711 129150 340720
rect 129004 324284 129056 324290
rect 129004 324226 129056 324232
rect 129002 317928 129058 317937
rect 129002 317863 129058 317872
rect 128358 310312 128414 310321
rect 128358 310247 128414 310256
rect 128372 309194 128400 310247
rect 11704 309188 11756 309194
rect 11704 309130 11756 309136
rect 128360 309188 128412 309194
rect 128360 309130 128412 309136
rect 8944 266076 8996 266082
rect 8944 266018 8996 266024
rect 8944 263628 8996 263634
rect 8944 263570 8996 263576
rect 7564 251660 7616 251666
rect 7564 251602 7616 251608
rect 7564 211200 7616 211206
rect 7564 211142 7616 211148
rect 6184 208208 6236 208214
rect 6184 208150 6236 208156
rect 6184 194608 6236 194614
rect 6184 194550 6236 194556
rect 3422 165064 3478 165073
rect 3422 164999 3478 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3424 136536 3476 136542
rect 3424 136478 3476 136484
rect 3436 136377 3464 136478
rect 3422 136368 3478 136377
rect 3422 136303 3478 136312
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3424 80028 3476 80034
rect 3424 79970 3476 79976
rect 3436 78985 3464 79970
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 6196 8158 6224 194550
rect 7576 35902 7604 211142
rect 8956 136542 8984 263570
rect 10324 256760 10376 256766
rect 10324 256702 10376 256708
rect 8944 136536 8996 136542
rect 8944 136478 8996 136484
rect 10336 122806 10364 256702
rect 11716 223582 11744 309130
rect 128358 302696 128414 302705
rect 128358 302631 128414 302640
rect 128372 302258 128400 302631
rect 128360 302252 128412 302258
rect 128360 302194 128412 302200
rect 128358 287464 128414 287473
rect 128358 287399 128414 287408
rect 128372 287094 128400 287399
rect 13084 287088 13136 287094
rect 13084 287030 13136 287036
rect 128360 287088 128412 287094
rect 128360 287030 128412 287036
rect 11704 223576 11756 223582
rect 11704 223518 11756 223524
rect 11704 218068 11756 218074
rect 11704 218010 11756 218016
rect 10324 122800 10376 122806
rect 10324 122742 10376 122748
rect 11716 51066 11744 218010
rect 13096 180810 13124 287030
rect 128266 279848 128322 279857
rect 128266 279783 128322 279792
rect 128280 278050 128308 279783
rect 128268 278044 128320 278050
rect 128268 277986 128320 277992
rect 128358 264480 128414 264489
rect 128358 264415 128414 264424
rect 128372 263634 128400 264415
rect 128360 263628 128412 263634
rect 128360 263570 128412 263576
rect 128358 256864 128414 256873
rect 128358 256799 128414 256808
rect 128372 256766 128400 256799
rect 128360 256760 128412 256766
rect 128360 256702 128412 256708
rect 128358 241632 128414 241641
rect 128358 241567 128414 241576
rect 128372 241534 128400 241567
rect 15844 241528 15896 241534
rect 15844 241470 15896 241476
rect 128360 241528 128412 241534
rect 128360 241470 128412 241476
rect 14464 233300 14516 233306
rect 14464 233242 14516 233248
rect 13084 180804 13136 180810
rect 13084 180746 13136 180752
rect 14476 80034 14504 233242
rect 15856 93838 15884 241470
rect 129016 237386 129044 317863
rect 129108 280158 129136 340711
rect 129200 309126 129228 356079
rect 129292 338094 129320 371311
rect 460216 366722 460244 391954
rect 578896 380866 578924 416463
rect 580276 396030 580304 451687
rect 580354 404832 580410 404841
rect 580354 404767 580410 404776
rect 580264 396024 580316 396030
rect 580264 395966 580316 395972
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 578884 380860 578936 380866
rect 578884 380802 578936 380808
rect 580368 373998 580396 404767
rect 580356 373992 580408 373998
rect 580356 373934 580408 373940
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 453948 366716 454000 366722
rect 453948 366658 454000 366664
rect 460204 366716 460256 366722
rect 460204 366658 460256 366664
rect 453960 366489 453988 366658
rect 453946 366480 454002 366489
rect 453946 366415 454002 366424
rect 580276 360194 580304 369543
rect 453948 360188 454000 360194
rect 453948 360130 454000 360136
rect 580264 360188 580316 360194
rect 580264 360130 580316 360136
rect 453960 359417 453988 360130
rect 453946 359408 454002 359417
rect 453946 359343 454002 359352
rect 580262 357912 580318 357921
rect 580262 357847 580318 357856
rect 580276 353258 580304 357847
rect 453764 353252 453816 353258
rect 453764 353194 453816 353200
rect 580264 353252 580316 353258
rect 580264 353194 580316 353200
rect 453776 352209 453804 353194
rect 453762 352200 453818 352209
rect 453762 352135 453818 352144
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345710 580212 346015
rect 453948 345704 454000 345710
rect 453948 345646 454000 345652
rect 580172 345704 580224 345710
rect 580172 345646 580224 345652
rect 453960 345137 453988 345646
rect 453946 345128 454002 345137
rect 453946 345063 454002 345072
rect 129280 338088 129332 338094
rect 129280 338030 129332 338036
rect 453486 338056 453542 338065
rect 453486 337991 453542 338000
rect 453394 330848 453450 330857
rect 453394 330783 453450 330792
rect 453302 323776 453358 323785
rect 453302 323711 453358 323720
rect 129188 309120 129240 309126
rect 129188 309062 129240 309068
rect 453316 299470 453344 323711
rect 453408 311846 453436 330783
rect 453500 322930 453528 337991
rect 453488 322924 453540 322930
rect 453488 322866 453540 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 453578 316704 453634 316713
rect 453578 316639 453634 316648
rect 453396 311840 453448 311846
rect 453396 311782 453448 311788
rect 453486 309496 453542 309505
rect 453486 309431 453542 309440
rect 453304 299464 453356 299470
rect 453304 299406 453356 299412
rect 453394 295216 453450 295225
rect 453394 295151 453450 295160
rect 129370 295080 129426 295089
rect 129370 295015 129426 295024
rect 129096 280152 129148 280158
rect 129096 280094 129148 280100
rect 129278 272096 129334 272105
rect 129278 272031 129334 272040
rect 129186 249248 129242 249257
rect 129186 249183 129242 249192
rect 129004 237380 129056 237386
rect 129004 237322 129056 237328
rect 128358 234016 128414 234025
rect 128358 233951 128414 233960
rect 128372 233306 128400 233951
rect 128360 233300 128412 233306
rect 128360 233242 128412 233248
rect 129094 226400 129150 226409
rect 129094 226335 129150 226344
rect 128358 218784 128414 218793
rect 128358 218719 128414 218728
rect 128372 218074 128400 218719
rect 128360 218068 128412 218074
rect 128360 218010 128412 218016
rect 128360 211200 128412 211206
rect 128358 211168 128360 211177
rect 128412 211168 128414 211177
rect 128358 211103 128414 211112
rect 129002 203552 129058 203561
rect 129002 203487 129058 203496
rect 128634 195936 128690 195945
rect 128634 195871 128690 195880
rect 128648 194614 128676 195871
rect 128636 194608 128688 194614
rect 128636 194550 128688 194556
rect 15844 93832 15896 93838
rect 15844 93774 15896 93780
rect 14464 80028 14516 80034
rect 14464 79970 14516 79976
rect 11704 51060 11756 51066
rect 11704 51002 11756 51008
rect 7564 35896 7616 35902
rect 7564 35838 7616 35844
rect 129016 22098 129044 203487
rect 129108 64870 129136 226335
rect 129200 109002 129228 249183
rect 129292 151774 129320 272031
rect 129384 194546 129412 295015
rect 453302 288144 453358 288153
rect 453302 288079 453358 288088
rect 453026 252512 453082 252521
rect 453026 252447 453082 252456
rect 453040 251258 453068 252447
rect 453028 251252 453080 251258
rect 453028 251194 453080 251200
rect 453118 231160 453174 231169
rect 453118 231095 453174 231104
rect 453132 230518 453160 231095
rect 453120 230512 453172 230518
rect 453120 230454 453172 230460
rect 453316 218006 453344 288079
rect 453408 229090 453436 295151
rect 453500 264926 453528 309431
rect 453592 276010 453620 316639
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 453670 302424 453726 302433
rect 453670 302359 453672 302368
rect 453724 302359 453726 302368
rect 456064 302388 456116 302394
rect 453672 302330 453724 302336
rect 456064 302330 456116 302336
rect 453946 281072 454002 281081
rect 453946 281007 454002 281016
rect 453960 280226 453988 281007
rect 453948 280220 454000 280226
rect 453948 280162 454000 280168
rect 453580 276004 453632 276010
rect 453580 275946 453632 275952
rect 453670 273864 453726 273873
rect 453670 273799 453726 273808
rect 453578 266792 453634 266801
rect 453578 266727 453634 266736
rect 453488 264920 453540 264926
rect 453488 264862 453540 264868
rect 453486 245440 453542 245449
rect 453486 245375 453542 245384
rect 453396 229084 453448 229090
rect 453396 229026 453448 229032
rect 453394 224088 453450 224097
rect 453394 224023 453450 224032
rect 453304 218000 453356 218006
rect 453304 217942 453356 217948
rect 453302 202736 453358 202745
rect 453302 202671 453358 202680
rect 129372 194540 129424 194546
rect 129372 194482 129424 194488
rect 135732 192222 136482 192250
rect 139872 192222 140622 192250
rect 131132 192086 132434 192114
rect 132512 192086 133170 192114
rect 133892 192086 133998 192114
rect 134168 192086 134826 192114
rect 135272 192086 135654 192114
rect 129280 151768 129332 151774
rect 129280 151710 129332 151716
rect 129188 108996 129240 109002
rect 129188 108938 129240 108944
rect 129096 64864 129148 64870
rect 129096 64806 129148 64812
rect 129004 22092 129056 22098
rect 129004 22034 129056 22040
rect 2780 8152 2832 8158
rect 2780 8094 2832 8100
rect 6184 8152 6236 8158
rect 6184 8094 6236 8100
rect 2792 7177 2820 8094
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 127808 4140 127860 4146
rect 127808 4082 127860 4088
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 126612 3120 126664 3126
rect 126612 3062 126664 3068
rect 126624 480 126652 3062
rect 127820 480 127848 4082
rect 130200 4072 130252 4078
rect 130200 4014 130252 4020
rect 129004 4004 129056 4010
rect 129004 3946 129056 3952
rect 129016 480 129044 3946
rect 130212 480 130240 4014
rect 131132 3466 131160 192086
rect 132512 3534 132540 192086
rect 132592 3596 132644 3602
rect 132592 3538 132644 3544
rect 132500 3528 132552 3534
rect 132500 3470 132552 3476
rect 131120 3460 131172 3466
rect 131120 3402 131172 3408
rect 131396 3052 131448 3058
rect 131396 2994 131448 3000
rect 131408 480 131436 2994
rect 132604 480 132632 3538
rect 133788 3256 133840 3262
rect 133788 3198 133840 3204
rect 133800 480 133828 3198
rect 133892 3126 133920 192086
rect 134168 4146 134196 192086
rect 134156 4140 134208 4146
rect 134156 4082 134208 4088
rect 135272 4010 135300 192086
rect 135732 189258 135760 192222
rect 135640 189230 135760 189258
rect 136652 192086 137310 192114
rect 138032 192086 138138 192114
rect 138308 192086 138966 192114
rect 139412 192086 139794 192114
rect 135640 186266 135668 189230
rect 135548 186238 135668 186266
rect 135548 183530 135576 186238
rect 135536 183524 135588 183530
rect 135536 183466 135588 183472
rect 135628 183524 135680 183530
rect 135628 183466 135680 183472
rect 135640 166954 135668 183466
rect 135456 166926 135668 166954
rect 135456 159338 135484 166926
rect 135364 159310 135484 159338
rect 135364 154562 135392 159310
rect 135352 154556 135404 154562
rect 135352 154498 135404 154504
rect 135444 147620 135496 147626
rect 135444 147562 135496 147568
rect 135456 143546 135484 147562
rect 135444 143540 135496 143546
rect 135444 143482 135496 143488
rect 135628 131504 135680 131510
rect 135628 131446 135680 131452
rect 135640 124166 135668 131446
rect 135628 124160 135680 124166
rect 135628 124102 135680 124108
rect 135812 124160 135864 124166
rect 135812 124102 135864 124108
rect 135824 122806 135852 124102
rect 135812 122800 135864 122806
rect 135812 122742 135864 122748
rect 135628 106208 135680 106214
rect 135628 106150 135680 106156
rect 135640 104854 135668 106150
rect 135628 104848 135680 104854
rect 135628 104790 135680 104796
rect 135536 89684 135588 89690
rect 135536 89626 135588 89632
rect 135548 86986 135576 89626
rect 135456 86970 135576 86986
rect 135444 86964 135576 86970
rect 135496 86958 135576 86964
rect 135720 86964 135772 86970
rect 135444 86906 135496 86912
rect 135720 86906 135772 86912
rect 135732 85542 135760 86906
rect 135720 85536 135772 85542
rect 135720 85478 135772 85484
rect 135720 77308 135772 77314
rect 135720 77250 135772 77256
rect 135732 66298 135760 77250
rect 135444 66292 135496 66298
rect 135444 66234 135496 66240
rect 135720 66292 135772 66298
rect 135720 66234 135772 66240
rect 135456 60858 135484 66234
rect 135444 60852 135496 60858
rect 135444 60794 135496 60800
rect 135444 57928 135496 57934
rect 135444 57870 135496 57876
rect 135456 43466 135484 57870
rect 135456 43438 135576 43466
rect 135548 31634 135576 43438
rect 135456 31606 135576 31634
rect 135456 27606 135484 31606
rect 135444 27600 135496 27606
rect 135444 27542 135496 27548
rect 135536 11756 135588 11762
rect 135536 11698 135588 11704
rect 135548 4078 135576 11698
rect 135536 4072 135588 4078
rect 135536 4014 135588 4020
rect 135260 4004 135312 4010
rect 135260 3946 135312 3952
rect 134892 3460 134944 3466
rect 134892 3402 134944 3408
rect 133880 3120 133932 3126
rect 133880 3062 133932 3068
rect 134904 480 134932 3402
rect 136088 3392 136140 3398
rect 136088 3334 136140 3340
rect 136100 480 136128 3334
rect 136652 3058 136680 192086
rect 138032 3602 138060 192086
rect 138020 3596 138072 3602
rect 138020 3538 138072 3544
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 136640 3052 136692 3058
rect 136640 2994 136692 3000
rect 137296 480 137324 3470
rect 138308 3262 138336 192086
rect 138480 3596 138532 3602
rect 138480 3538 138532 3544
rect 138296 3256 138348 3262
rect 138296 3198 138348 3204
rect 138492 480 138520 3538
rect 139412 3466 139440 192086
rect 139872 189258 139900 192222
rect 139780 189230 139900 189258
rect 140792 192086 141450 192114
rect 139780 176746 139808 189230
rect 139688 176718 139808 176746
rect 139688 176610 139716 176718
rect 139596 176582 139716 176610
rect 139596 167090 139624 176582
rect 139504 167062 139624 167090
rect 139400 3460 139452 3466
rect 139400 3402 139452 3408
rect 139504 3398 139532 167062
rect 139676 3936 139728 3942
rect 139676 3878 139728 3884
rect 139492 3392 139544 3398
rect 139492 3334 139544 3340
rect 139688 480 139716 3878
rect 140792 3534 140820 192086
rect 142160 181484 142212 181490
rect 142160 181426 142212 181432
rect 140872 4072 140924 4078
rect 140872 4014 140924 4020
rect 140780 3528 140832 3534
rect 140780 3470 140832 3476
rect 140884 480 140912 4014
rect 142172 3942 142200 181426
rect 142160 3936 142212 3942
rect 142160 3878 142212 3884
rect 142068 3868 142120 3874
rect 142068 3810 142120 3816
rect 142080 480 142108 3810
rect 142264 3602 142292 192100
rect 142816 192086 143106 192114
rect 143552 192086 143934 192114
rect 144012 192086 144762 192114
rect 144932 192086 145590 192114
rect 142816 181490 142844 192086
rect 142804 181484 142856 181490
rect 142804 181426 142856 181432
rect 143552 4078 143580 192086
rect 144012 183569 144040 192086
rect 143998 183560 144054 183569
rect 143998 183495 144054 183504
rect 144182 183560 144238 183569
rect 144182 183495 144238 183504
rect 144196 173942 144224 183495
rect 143908 173936 143960 173942
rect 143908 173878 143960 173884
rect 144184 173936 144236 173942
rect 144184 173878 144236 173884
rect 143920 166954 143948 173878
rect 143828 166926 143948 166954
rect 143828 164218 143856 166926
rect 143632 164212 143684 164218
rect 143632 164154 143684 164160
rect 143816 164212 143868 164218
rect 143816 164154 143868 164160
rect 143644 154601 143672 164154
rect 143630 154592 143686 154601
rect 143630 154527 143686 154536
rect 143906 154592 143962 154601
rect 143906 154527 143962 154536
rect 143920 147642 143948 154527
rect 143828 147614 143948 147642
rect 143828 143546 143856 147614
rect 143816 143540 143868 143546
rect 143816 143482 143868 143488
rect 143816 128308 143868 128314
rect 143816 128250 143868 128256
rect 143828 120714 143856 128250
rect 143644 120686 143856 120714
rect 143644 115977 143672 120686
rect 143630 115968 143686 115977
rect 143630 115903 143686 115912
rect 143906 115968 143962 115977
rect 143906 115903 143962 115912
rect 143920 109018 143948 115903
rect 143828 108990 143948 109018
rect 143828 101402 143856 108990
rect 143644 101374 143856 101402
rect 143644 96665 143672 101374
rect 143630 96656 143686 96665
rect 143630 96591 143686 96600
rect 143906 96656 143962 96665
rect 143906 96591 143962 96600
rect 143920 89706 143948 96591
rect 143736 89678 143948 89706
rect 143736 86970 143764 89678
rect 143724 86964 143776 86970
rect 143724 86906 143776 86912
rect 143632 77308 143684 77314
rect 143632 77250 143684 77256
rect 143644 70258 143672 77250
rect 143644 70230 143764 70258
rect 143736 60722 143764 70230
rect 143724 60716 143776 60722
rect 143724 60658 143776 60664
rect 143908 60716 143960 60722
rect 143908 60658 143960 60664
rect 143920 57934 143948 60658
rect 143908 57928 143960 57934
rect 143908 57870 143960 57876
rect 143724 48340 143776 48346
rect 143724 48282 143776 48288
rect 143736 38690 143764 48282
rect 143724 38684 143776 38690
rect 143724 38626 143776 38632
rect 143908 38684 143960 38690
rect 143908 38626 143960 38632
rect 143920 29050 143948 38626
rect 143736 29022 143948 29050
rect 143736 27606 143764 29022
rect 143724 27600 143776 27606
rect 143724 27542 143776 27548
rect 144000 27600 144052 27606
rect 144000 27542 144052 27548
rect 144012 12458 144040 27542
rect 143920 12430 144040 12458
rect 143540 4072 143592 4078
rect 143540 4014 143592 4020
rect 143920 3874 143948 12430
rect 144460 4140 144512 4146
rect 144460 4082 144512 4088
rect 143908 3868 143960 3874
rect 143908 3810 143960 3816
rect 143264 3800 143316 3806
rect 143264 3742 143316 3748
rect 142252 3596 142304 3602
rect 142252 3538 142304 3544
rect 143276 480 143304 3742
rect 144472 480 144500 4082
rect 144932 3806 144960 192086
rect 146300 180940 146352 180946
rect 146300 180882 146352 180888
rect 144920 3800 144972 3806
rect 144920 3742 144972 3748
rect 146312 3330 146340 180882
rect 146404 4146 146432 192100
rect 146864 192086 147246 192114
rect 147784 192086 148074 192114
rect 148520 192086 148902 192114
rect 149072 192086 149730 192114
rect 146864 180946 146892 192086
rect 147680 185632 147732 185638
rect 147680 185574 147732 185580
rect 146852 180940 146904 180946
rect 146852 180882 146904 180888
rect 146392 4140 146444 4146
rect 146392 4082 146444 4088
rect 146852 3596 146904 3602
rect 146852 3538 146904 3544
rect 145656 3324 145708 3330
rect 145656 3266 145708 3272
rect 146300 3324 146352 3330
rect 146300 3266 146352 3272
rect 145668 480 145696 3266
rect 146864 480 146892 3538
rect 147692 3482 147720 185574
rect 147784 3602 147812 192086
rect 148520 185638 148548 192086
rect 148508 185632 148560 185638
rect 148508 185574 148560 185580
rect 147772 3596 147824 3602
rect 147772 3538 147824 3544
rect 147692 3454 148088 3482
rect 148060 480 148088 3454
rect 149072 3346 149100 192086
rect 150440 185632 150492 185638
rect 150440 185574 150492 185580
rect 150452 3602 150480 185574
rect 150440 3596 150492 3602
rect 150440 3538 150492 3544
rect 150544 3482 150572 192100
rect 151096 192086 151386 192114
rect 151832 192086 152214 192114
rect 153042 192086 153148 192114
rect 153870 192086 154528 192114
rect 151096 185638 151124 192086
rect 151084 185632 151136 185638
rect 151084 185574 151136 185580
rect 151544 3596 151596 3602
rect 151544 3538 151596 3544
rect 150452 3454 150572 3482
rect 149072 3318 149284 3346
rect 149256 480 149284 3318
rect 150452 480 150480 3454
rect 151556 480 151584 3538
rect 151832 3534 151860 192086
rect 153120 3534 153148 192086
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 152740 3528 152792 3534
rect 152740 3470 152792 3476
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 153936 3528 153988 3534
rect 153936 3470 153988 3476
rect 152752 480 152780 3470
rect 153948 480 153976 3470
rect 154500 3466 154528 192086
rect 154684 190126 154712 192100
rect 155434 192086 155908 192114
rect 154672 190120 154724 190126
rect 154672 190062 154724 190068
rect 155776 190120 155828 190126
rect 155776 190062 155828 190068
rect 155788 3534 155816 190062
rect 155776 3528 155828 3534
rect 155776 3470 155828 3476
rect 154488 3460 154540 3466
rect 154488 3402 154540 3408
rect 155132 3460 155184 3466
rect 155132 3402 155184 3408
rect 155144 480 155172 3402
rect 155880 3330 155908 192086
rect 156248 189378 156276 192100
rect 157090 192086 157196 192114
rect 156236 189372 156288 189378
rect 156236 189314 156288 189320
rect 156328 3528 156380 3534
rect 156328 3470 156380 3476
rect 155868 3324 155920 3330
rect 155868 3266 155920 3272
rect 156340 480 156368 3470
rect 157168 3058 157196 192086
rect 157248 189372 157300 189378
rect 157248 189314 157300 189320
rect 157260 3534 157288 189314
rect 157904 189106 157932 192100
rect 158732 189854 158760 192100
rect 159574 192086 160048 192114
rect 158720 189848 158772 189854
rect 158720 189790 158772 189796
rect 159916 189848 159968 189854
rect 159916 189790 159968 189796
rect 157892 189100 157944 189106
rect 157892 189042 157944 189048
rect 158628 189100 158680 189106
rect 158628 189042 158680 189048
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 158640 3466 158668 189042
rect 159928 4078 159956 189790
rect 160020 4146 160048 192086
rect 160388 189174 160416 192100
rect 161230 192086 161336 192114
rect 162058 192086 162808 192114
rect 160376 189168 160428 189174
rect 160376 189110 160428 189116
rect 160008 4140 160060 4146
rect 160008 4082 160060 4088
rect 159916 4072 159968 4078
rect 159916 4014 159968 4020
rect 158720 3528 158772 3534
rect 158720 3470 158772 3476
rect 158628 3460 158680 3466
rect 158628 3402 158680 3408
rect 157524 3324 157576 3330
rect 157524 3266 157576 3272
rect 157156 3052 157208 3058
rect 157156 2994 157208 3000
rect 157536 480 157564 3266
rect 158732 480 158760 3470
rect 161308 3466 161336 192086
rect 161388 189168 161440 189174
rect 161388 189110 161440 189116
rect 161400 3602 161428 189110
rect 162308 4072 162360 4078
rect 162308 4014 162360 4020
rect 161388 3596 161440 3602
rect 161388 3538 161440 3544
rect 161112 3460 161164 3466
rect 161112 3402 161164 3408
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 159916 3052 159968 3058
rect 159916 2994 159968 3000
rect 159928 480 159956 2994
rect 161124 480 161152 3402
rect 162320 480 162348 4014
rect 162780 3534 162808 192086
rect 162872 189990 162900 192100
rect 163714 192086 164188 192114
rect 162860 189984 162912 189990
rect 162860 189926 162912 189932
rect 164056 189984 164108 189990
rect 164056 189926 164108 189932
rect 163504 4140 163556 4146
rect 163504 4082 163556 4088
rect 162768 3528 162820 3534
rect 162768 3470 162820 3476
rect 163516 480 163544 4082
rect 164068 3330 164096 189926
rect 164056 3324 164108 3330
rect 164056 3266 164108 3272
rect 164160 3194 164188 192086
rect 164528 190126 164556 192100
rect 165370 192086 165568 192114
rect 164516 190120 164568 190126
rect 164516 190062 164568 190068
rect 165436 190120 165488 190126
rect 165436 190062 165488 190068
rect 165448 3602 165476 190062
rect 164700 3596 164752 3602
rect 164700 3538 164752 3544
rect 165436 3596 165488 3602
rect 165436 3538 165488 3544
rect 164148 3188 164200 3194
rect 164148 3130 164200 3136
rect 164712 480 164740 3538
rect 165540 3058 165568 192086
rect 166184 189106 166212 192100
rect 167012 189106 167040 192100
rect 167854 192086 168328 192114
rect 166172 189100 166224 189106
rect 166172 189042 166224 189048
rect 166908 189100 166960 189106
rect 166908 189042 166960 189048
rect 167000 189100 167052 189106
rect 167000 189042 167052 189048
rect 168196 189100 168248 189106
rect 168196 189042 168248 189048
rect 166920 4146 166948 189042
rect 166908 4140 166960 4146
rect 166908 4082 166960 4088
rect 168208 3670 168236 189042
rect 168196 3664 168248 3670
rect 168196 3606 168248 3612
rect 168300 3534 168328 192086
rect 168668 190330 168696 192100
rect 169510 192086 169708 192114
rect 170338 192086 171088 192114
rect 168656 190324 168708 190330
rect 168656 190266 168708 190272
rect 169576 190324 169628 190330
rect 169576 190266 169628 190272
rect 169588 3942 169616 190266
rect 169576 3936 169628 3942
rect 169576 3878 169628 3884
rect 169680 3874 169708 192086
rect 169668 3868 169720 3874
rect 169668 3810 169720 3816
rect 170588 3596 170640 3602
rect 170588 3538 170640 3544
rect 167092 3528 167144 3534
rect 167092 3470 167144 3476
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 165896 3460 165948 3466
rect 165896 3402 165948 3408
rect 165528 3052 165580 3058
rect 165528 2994 165580 3000
rect 165908 480 165936 3402
rect 167104 480 167132 3470
rect 168196 3324 168248 3330
rect 168196 3266 168248 3272
rect 168208 480 168236 3266
rect 169392 3188 169444 3194
rect 169392 3130 169444 3136
rect 169404 480 169432 3130
rect 170600 480 170628 3538
rect 171060 3466 171088 192086
rect 171152 189106 171180 192100
rect 171994 192086 172376 192114
rect 171140 189100 171192 189106
rect 171140 189042 171192 189048
rect 172348 3602 172376 192086
rect 172808 189378 172836 192100
rect 173650 192086 173756 192114
rect 172796 189372 172848 189378
rect 172796 189314 172848 189320
rect 172428 189100 172480 189106
rect 172428 189042 172480 189048
rect 172336 3596 172388 3602
rect 172336 3538 172388 3544
rect 171048 3460 171100 3466
rect 171048 3402 171100 3408
rect 171784 3052 171836 3058
rect 171784 2994 171836 3000
rect 171796 480 171824 2994
rect 172440 2990 172468 189042
rect 173728 4826 173756 192086
rect 173808 189372 173860 189378
rect 173808 189314 173860 189320
rect 173716 4820 173768 4826
rect 173716 4762 173768 4768
rect 172980 4140 173032 4146
rect 172980 4082 173032 4088
rect 172428 2984 172480 2990
rect 172428 2926 172480 2932
rect 172992 480 173020 4082
rect 173820 3738 173848 189314
rect 174464 189106 174492 192100
rect 175292 189310 175320 192100
rect 176134 192086 176516 192114
rect 175280 189304 175332 189310
rect 175280 189246 175332 189252
rect 174452 189100 174504 189106
rect 174452 189042 174504 189048
rect 175188 189100 175240 189106
rect 175188 189042 175240 189048
rect 173808 3732 173860 3738
rect 173808 3674 173860 3680
rect 175200 3670 175228 189042
rect 176488 6186 176516 192086
rect 176568 189304 176620 189310
rect 176568 189246 176620 189252
rect 176476 6180 176528 6186
rect 176476 6122 176528 6128
rect 176580 4010 176608 189246
rect 176948 189106 176976 192100
rect 177790 192086 177988 192114
rect 176936 189100 176988 189106
rect 176936 189042 176988 189048
rect 177856 189100 177908 189106
rect 177856 189042 177908 189048
rect 176568 4004 176620 4010
rect 176568 3946 176620 3952
rect 177868 3942 177896 189042
rect 176476 3936 176528 3942
rect 177856 3936 177908 3942
rect 176528 3884 176608 3890
rect 176476 3878 176608 3884
rect 177856 3878 177908 3884
rect 176488 3862 176608 3878
rect 174176 3664 174228 3670
rect 174176 3606 174228 3612
rect 175188 3664 175240 3670
rect 175188 3606 175240 3612
rect 174188 480 174216 3606
rect 175372 3528 175424 3534
rect 175372 3470 175424 3476
rect 175384 480 175412 3470
rect 176580 480 176608 3862
rect 177764 3868 177816 3874
rect 177764 3810 177816 3816
rect 177776 480 177804 3810
rect 177960 3534 177988 192086
rect 178512 189854 178540 192100
rect 178500 189848 178552 189854
rect 178500 189790 178552 189796
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179340 3466 179368 192100
rect 180182 192086 180748 192114
rect 180720 3738 180748 192086
rect 180996 189786 181024 192100
rect 181838 192086 182128 192114
rect 180984 189780 181036 189786
rect 180984 189722 181036 189728
rect 182100 3874 182128 192086
rect 182652 189446 182680 192100
rect 183388 192086 183494 192114
rect 184322 192086 184888 192114
rect 182640 189440 182692 189446
rect 182640 189382 182692 189388
rect 183388 7614 183416 192086
rect 183468 189440 183520 189446
rect 183468 189382 183520 189388
rect 183376 7608 183428 7614
rect 183376 7550 183428 7556
rect 182088 3868 182140 3874
rect 182088 3810 182140 3816
rect 183480 3806 183508 189382
rect 184860 11762 184888 192086
rect 185136 189310 185164 192100
rect 185978 192086 186176 192114
rect 185124 189304 185176 189310
rect 185124 189246 185176 189252
rect 184848 11756 184900 11762
rect 184848 11698 184900 11704
rect 186148 6254 186176 192086
rect 186228 189304 186280 189310
rect 186228 189246 186280 189252
rect 186136 6248 186188 6254
rect 186136 6190 186188 6196
rect 183744 4820 183796 4826
rect 183744 4762 183796 4768
rect 182548 3800 182600 3806
rect 182548 3742 182600 3748
rect 183468 3800 183520 3806
rect 183468 3742 183520 3748
rect 180708 3732 180760 3738
rect 180708 3674 180760 3680
rect 181352 3596 181404 3602
rect 181352 3538 181404 3544
rect 178960 3460 179012 3466
rect 178960 3402 179012 3408
rect 179328 3460 179380 3466
rect 179328 3402 179380 3408
rect 178972 480 179000 3402
rect 180156 2984 180208 2990
rect 180156 2926 180208 2932
rect 180168 480 180196 2926
rect 181364 480 181392 3538
rect 182560 480 182588 3742
rect 183756 480 183784 4762
rect 186044 4004 186096 4010
rect 186044 3946 186096 3952
rect 184848 3664 184900 3670
rect 184848 3606 184900 3612
rect 184860 480 184888 3606
rect 186056 480 186084 3946
rect 186240 3670 186268 189246
rect 186792 189106 186820 192100
rect 186780 189100 186832 189106
rect 186780 189042 186832 189048
rect 187516 189100 187568 189106
rect 187516 189042 187568 189048
rect 187528 13122 187556 189042
rect 187516 13116 187568 13122
rect 187516 13058 187568 13064
rect 187240 6180 187292 6186
rect 187240 6122 187292 6128
rect 186228 3664 186280 3670
rect 186228 3606 186280 3612
rect 187252 480 187280 6122
rect 187620 3602 187648 192100
rect 188462 192086 189028 192114
rect 188344 189848 188396 189854
rect 188344 189790 188396 189796
rect 188356 4894 188384 189790
rect 189000 10334 189028 192086
rect 189276 189106 189304 192100
rect 190118 192086 190408 192114
rect 189264 189100 189316 189106
rect 189264 189042 189316 189048
rect 190276 189100 190328 189106
rect 190276 189042 190328 189048
rect 190288 14482 190316 189042
rect 190276 14476 190328 14482
rect 190276 14418 190328 14424
rect 188988 10328 189040 10334
rect 188988 10270 189040 10276
rect 188344 4888 188396 4894
rect 188344 4830 188396 4836
rect 188436 3936 188488 3942
rect 188436 3878 188488 3884
rect 187608 3596 187660 3602
rect 187608 3538 187660 3544
rect 188448 480 188476 3878
rect 190380 3534 190408 192086
rect 190932 189106 190960 192100
rect 191668 192086 191774 192114
rect 192602 192086 193168 192114
rect 190920 189100 190972 189106
rect 190920 189042 190972 189048
rect 191668 15910 191696 192086
rect 192484 189780 192536 189786
rect 192484 189722 192536 189728
rect 191748 189100 191800 189106
rect 191748 189042 191800 189048
rect 191656 15904 191708 15910
rect 191656 15846 191708 15852
rect 191760 8974 191788 189042
rect 191748 8968 191800 8974
rect 191748 8910 191800 8916
rect 190828 4888 190880 4894
rect 190828 4830 190880 4836
rect 189632 3528 189684 3534
rect 189632 3470 189684 3476
rect 190368 3528 190420 3534
rect 190368 3470 190420 3476
rect 189644 480 189672 3470
rect 190840 480 190868 4830
rect 192496 4214 192524 189722
rect 192484 4208 192536 4214
rect 192484 4150 192536 4156
rect 193140 3466 193168 192086
rect 193416 189310 193444 192100
rect 194258 192086 194456 192114
rect 193404 189304 193456 189310
rect 193404 189246 193456 189252
rect 194428 17270 194456 192086
rect 194508 189304 194560 189310
rect 194508 189246 194560 189252
rect 194416 17264 194468 17270
rect 194416 17206 194468 17212
rect 194520 4826 194548 189246
rect 195072 189106 195100 192100
rect 195900 189786 195928 192100
rect 196742 192086 197308 192114
rect 195888 189780 195940 189786
rect 195888 189722 195940 189728
rect 195060 189100 195112 189106
rect 195060 189042 195112 189048
rect 195888 189100 195940 189106
rect 195888 189042 195940 189048
rect 194508 4820 194560 4826
rect 194508 4762 194560 4768
rect 194416 4208 194468 4214
rect 194416 4150 194468 4156
rect 193220 3732 193272 3738
rect 193220 3674 193272 3680
rect 192024 3460 192076 3466
rect 192024 3402 192076 3408
rect 193128 3460 193180 3466
rect 193128 3402 193180 3408
rect 192036 480 192064 3402
rect 193232 480 193260 3674
rect 194428 480 194456 4150
rect 195900 3942 195928 189042
rect 197280 18698 197308 192086
rect 197556 189378 197584 192100
rect 198398 192086 198596 192114
rect 197544 189372 197596 189378
rect 197544 189314 197596 189320
rect 197268 18692 197320 18698
rect 197268 18634 197320 18640
rect 198568 7614 198596 192086
rect 198648 189372 198700 189378
rect 198648 189314 198700 189320
rect 198004 7608 198056 7614
rect 198004 7550 198056 7556
rect 198556 7608 198608 7614
rect 198556 7550 198608 7556
rect 195888 3936 195940 3942
rect 195888 3878 195940 3884
rect 195612 3868 195664 3874
rect 195612 3810 195664 3816
rect 195624 480 195652 3810
rect 196808 3800 196860 3806
rect 196808 3742 196860 3748
rect 196820 480 196848 3742
rect 198016 480 198044 7550
rect 198660 3874 198688 189314
rect 199212 189106 199240 192100
rect 199200 189100 199252 189106
rect 199200 189042 199252 189048
rect 198740 11756 198792 11762
rect 198740 11698 198792 11704
rect 198648 3868 198700 3874
rect 198648 3810 198700 3816
rect 198752 3346 198780 11698
rect 200040 3806 200068 192100
rect 200790 192086 201448 192114
rect 200764 189100 200816 189106
rect 200764 189042 200816 189048
rect 200776 20058 200804 189042
rect 200764 20052 200816 20058
rect 200764 19994 200816 20000
rect 201420 6186 201448 192086
rect 201604 190262 201632 192100
rect 202446 192086 202828 192114
rect 201592 190256 201644 190262
rect 201592 190198 201644 190204
rect 201500 13116 201552 13122
rect 201500 13058 201552 13064
rect 201408 6180 201460 6186
rect 201408 6122 201460 6128
rect 200028 3800 200080 3806
rect 200028 3742 200080 3748
rect 200396 3664 200448 3670
rect 200396 3606 200448 3612
rect 198752 3318 199240 3346
rect 199212 480 199240 3318
rect 200408 480 200436 3606
rect 201512 3534 201540 13058
rect 201592 6248 201644 6254
rect 201592 6190 201644 6196
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 201604 3346 201632 6190
rect 202800 3670 202828 192086
rect 203260 189446 203288 192100
rect 203248 189440 203300 189446
rect 203248 189382 203300 189388
rect 204088 22778 204116 192100
rect 204930 192086 205588 192114
rect 204904 190256 204956 190262
rect 204904 190198 204956 190204
rect 204168 189440 204220 189446
rect 204168 189382 204220 189388
rect 204076 22772 204128 22778
rect 204076 22714 204128 22720
rect 204180 11762 204208 189382
rect 204916 21486 204944 190198
rect 204904 21480 204956 21486
rect 204904 21422 204956 21428
rect 204168 11756 204220 11762
rect 204168 11698 204220 11704
rect 204260 10328 204312 10334
rect 204260 10270 204312 10276
rect 202788 3664 202840 3670
rect 202788 3606 202840 3612
rect 203892 3596 203944 3602
rect 203892 3538 203944 3544
rect 202696 3528 202748 3534
rect 202696 3470 202748 3476
rect 201512 3318 201632 3346
rect 201512 480 201540 3318
rect 202708 480 202736 3470
rect 203904 480 203932 3538
rect 204272 3346 204300 10270
rect 205560 3738 205588 192086
rect 205744 189310 205772 192100
rect 206586 192086 206876 192114
rect 205732 189304 205784 189310
rect 205732 189246 205784 189252
rect 206848 24138 206876 192086
rect 206928 189304 206980 189310
rect 206928 189246 206980 189252
rect 206836 24132 206888 24138
rect 206836 24074 206888 24080
rect 205640 14476 205692 14482
rect 205640 14418 205692 14424
rect 205548 3732 205600 3738
rect 205548 3674 205600 3680
rect 205652 3346 205680 14418
rect 206940 10334 206968 189246
rect 207400 189106 207428 192100
rect 207388 189100 207440 189106
rect 207388 189042 207440 189048
rect 208228 13122 208256 192100
rect 209070 192086 209728 192114
rect 208308 189100 208360 189106
rect 208308 189042 208360 189048
rect 208216 13116 208268 13122
rect 208216 13058 208268 13064
rect 206928 10328 206980 10334
rect 206928 10270 206980 10276
rect 208320 3602 208348 189042
rect 209700 15978 209728 192086
rect 209884 189310 209912 192100
rect 210726 192086 211016 192114
rect 209872 189304 209924 189310
rect 209872 189246 209924 189252
rect 209688 15972 209740 15978
rect 209688 15914 209740 15920
rect 209872 15904 209924 15910
rect 209872 15846 209924 15852
rect 208676 8968 208728 8974
rect 208676 8910 208728 8916
rect 208308 3596 208360 3602
rect 208308 3538 208360 3544
rect 207480 3392 207532 3398
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 207480 3334 207532 3340
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3334
rect 208688 480 208716 8910
rect 209884 480 209912 15846
rect 210988 8974 211016 192086
rect 211068 189304 211120 189310
rect 211068 189246 211120 189252
rect 210976 8968 211028 8974
rect 210976 8910 211028 8916
rect 211080 3618 211108 189246
rect 211540 189106 211568 192100
rect 212382 192086 212488 192114
rect 213210 192086 213592 192114
rect 211528 189100 211580 189106
rect 211528 189042 211580 189048
rect 212356 189100 212408 189106
rect 212356 189042 212408 189048
rect 212368 25634 212396 189042
rect 212356 25628 212408 25634
rect 212356 25570 212408 25576
rect 212264 4820 212316 4826
rect 212264 4762 212316 4768
rect 211080 3590 211200 3618
rect 211172 3534 211200 3590
rect 211160 3528 211212 3534
rect 211160 3470 211212 3476
rect 211068 3460 211120 3466
rect 211068 3402 211120 3408
rect 211080 480 211108 3402
rect 212276 480 212304 4762
rect 212460 3466 212488 192086
rect 213184 189780 213236 189786
rect 213184 189722 213236 189728
rect 212540 17264 212592 17270
rect 212540 17206 212592 17212
rect 212552 3618 212580 17206
rect 213196 4214 213224 189722
rect 213564 189174 213592 192086
rect 214024 189378 214052 192100
rect 214866 192086 215156 192114
rect 214012 189372 214064 189378
rect 214012 189314 214064 189320
rect 213552 189168 213604 189174
rect 213552 189110 213604 189116
rect 215128 32434 215156 192086
rect 215208 189372 215260 189378
rect 215208 189314 215260 189320
rect 215116 32428 215168 32434
rect 215116 32370 215168 32376
rect 215220 17270 215248 189314
rect 215680 189106 215708 192100
rect 215668 189100 215720 189106
rect 215668 189042 215720 189048
rect 216508 18630 216536 192100
rect 217350 192086 218008 192114
rect 216588 189100 216640 189106
rect 216588 189042 216640 189048
rect 216496 18624 216548 18630
rect 216496 18566 216548 18572
rect 215208 17264 215260 17270
rect 215208 17206 215260 17212
rect 216600 14482 216628 189042
rect 217980 33794 218008 192086
rect 218164 189106 218192 192100
rect 219006 192086 219296 192114
rect 218152 189100 218204 189106
rect 218152 189042 218204 189048
rect 217968 33788 218020 33794
rect 217968 33730 218020 33736
rect 219268 19990 219296 192086
rect 219820 189446 219848 192100
rect 220662 192086 220768 192114
rect 219808 189440 219860 189446
rect 219808 189382 219860 189388
rect 220636 189440 220688 189446
rect 220636 189382 220688 189388
rect 219348 189100 219400 189106
rect 219348 189042 219400 189048
rect 219256 19984 219308 19990
rect 219256 19926 219308 19932
rect 216680 18692 216732 18698
rect 216680 18634 216732 18640
rect 216588 14476 216640 14482
rect 216588 14418 216640 14424
rect 213184 4208 213236 4214
rect 213184 4150 213236 4156
rect 215852 4208 215904 4214
rect 215852 4150 215904 4156
rect 214656 3936 214708 3942
rect 214656 3878 214708 3884
rect 212552 3590 213500 3618
rect 212448 3460 212500 3466
rect 212448 3402 212500 3408
rect 213472 480 213500 3590
rect 214668 480 214696 3878
rect 215864 480 215892 4150
rect 216692 3482 216720 18634
rect 219360 7614 219388 189042
rect 220648 36582 220676 189382
rect 220740 188358 220768 192086
rect 221476 189310 221504 192100
rect 222304 189514 222332 192100
rect 223132 189786 223160 192100
rect 223120 189780 223172 189786
rect 223120 189722 223172 189728
rect 222292 189508 222344 189514
rect 222292 189450 222344 189456
rect 223488 189508 223540 189514
rect 223488 189450 223540 189456
rect 221464 189304 221516 189310
rect 221464 189246 221516 189252
rect 222844 189304 222896 189310
rect 222844 189246 222896 189252
rect 221464 189168 221516 189174
rect 221464 189110 221516 189116
rect 220728 188352 220780 188358
rect 220728 188294 220780 188300
rect 220636 36576 220688 36582
rect 220636 36518 220688 36524
rect 219440 20052 219492 20058
rect 219440 19994 219492 20000
rect 219348 7608 219400 7614
rect 219348 7550 219400 7556
rect 219348 7404 219400 7410
rect 219348 7346 219400 7352
rect 218152 3868 218204 3874
rect 218152 3810 218204 3816
rect 216692 3454 217088 3482
rect 217060 480 217088 3454
rect 218164 480 218192 3810
rect 219360 480 219388 7346
rect 219452 3346 219480 19994
rect 221476 4826 221504 189110
rect 222856 21418 222884 189246
rect 223500 178702 223528 189450
rect 223868 189310 223896 192100
rect 224710 192086 224816 192114
rect 225538 192086 226288 192114
rect 223856 189304 223908 189310
rect 223856 189246 223908 189252
rect 223488 178696 223540 178702
rect 223488 178638 223540 178644
rect 224788 39370 224816 192086
rect 224868 189304 224920 189310
rect 224868 189246 224920 189252
rect 224776 39364 224828 39370
rect 224776 39306 224828 39312
rect 224880 26926 224908 189246
rect 224868 26920 224920 26926
rect 224868 26862 224920 26868
rect 223580 21480 223632 21486
rect 223580 21422 223632 21428
rect 222844 21412 222896 21418
rect 222844 21354 222896 21360
rect 222936 6180 222988 6186
rect 222936 6122 222988 6128
rect 221464 4820 221516 4826
rect 221464 4762 221516 4768
rect 221740 3800 221792 3806
rect 221740 3742 221792 3748
rect 219452 3318 220584 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3742
rect 222948 480 222976 6122
rect 223592 3346 223620 21422
rect 226260 6186 226288 192086
rect 226352 190058 226380 192100
rect 227194 192086 227668 192114
rect 226340 190052 226392 190058
rect 226340 189994 226392 190000
rect 227536 190052 227588 190058
rect 227536 189994 227588 190000
rect 227548 177342 227576 189994
rect 227536 177336 227588 177342
rect 227536 177278 227588 177284
rect 227640 40730 227668 192086
rect 228008 189106 228036 192100
rect 228850 192086 228956 192114
rect 227996 189100 228048 189106
rect 227996 189042 228048 189048
rect 227628 40724 227680 40730
rect 227628 40666 227680 40672
rect 228928 22778 228956 192086
rect 229664 189718 229692 192100
rect 229652 189712 229704 189718
rect 229652 189654 229704 189660
rect 230388 189712 230440 189718
rect 230388 189654 230440 189660
rect 229008 189100 229060 189106
rect 229008 189042 229060 189048
rect 227812 22772 227864 22778
rect 227812 22714 227864 22720
rect 228916 22772 228968 22778
rect 228916 22714 228968 22720
rect 226340 11756 226392 11762
rect 226340 11698 226392 11704
rect 226248 6180 226300 6186
rect 226248 6122 226300 6128
rect 225328 3664 225380 3670
rect 225328 3606 225380 3612
rect 223592 3318 224172 3346
rect 224144 480 224172 3318
rect 225340 480 225368 3606
rect 226352 3346 226380 11698
rect 226352 3318 226564 3346
rect 226536 480 226564 3318
rect 227824 1442 227852 22714
rect 229020 11762 229048 189042
rect 230400 42090 230428 189654
rect 230492 189310 230520 192100
rect 231334 192086 231716 192114
rect 230480 189304 230532 189310
rect 230480 189246 230532 189252
rect 230388 42084 230440 42090
rect 230388 42026 230440 42032
rect 231688 24138 231716 192086
rect 231768 189304 231820 189310
rect 231768 189246 231820 189252
rect 230480 24132 230532 24138
rect 230480 24074 230532 24080
rect 231676 24132 231728 24138
rect 231676 24074 231728 24080
rect 229008 11756 229060 11762
rect 229008 11698 229060 11704
rect 229100 10328 229152 10334
rect 229100 10270 229152 10276
rect 228916 3732 228968 3738
rect 228916 3674 228968 3680
rect 227732 1414 227852 1442
rect 227732 480 227760 1414
rect 228928 480 228956 3674
rect 229112 3482 229140 10270
rect 230492 3482 230520 24074
rect 231780 10334 231808 189246
rect 232148 189106 232176 192100
rect 232990 192086 233188 192114
rect 233818 192086 234568 192114
rect 232136 189100 232188 189106
rect 232136 189042 232188 189048
rect 233056 189100 233108 189106
rect 233056 189042 233108 189048
rect 233068 44878 233096 189042
rect 233056 44872 233108 44878
rect 233056 44814 233108 44820
rect 233160 15910 233188 192086
rect 234540 28286 234568 192086
rect 234632 189310 234660 192100
rect 234620 189304 234672 189310
rect 234620 189246 234672 189252
rect 235460 186998 235488 192100
rect 236288 189378 236316 192100
rect 237130 192086 237236 192114
rect 236276 189372 236328 189378
rect 236276 189314 236328 189320
rect 235908 189304 235960 189310
rect 235908 189246 235960 189252
rect 235448 186992 235500 186998
rect 235448 186934 235500 186940
rect 235920 46238 235948 189246
rect 237208 47598 237236 192086
rect 237944 189990 237972 192100
rect 237932 189984 237984 189990
rect 237932 189926 237984 189932
rect 238668 189984 238720 189990
rect 238668 189926 238720 189932
rect 237288 189372 237340 189378
rect 237288 189314 237340 189320
rect 237196 47592 237248 47598
rect 237196 47534 237248 47540
rect 235908 46232 235960 46238
rect 235908 46174 235960 46180
rect 234528 28280 234580 28286
rect 234528 28222 234580 28228
rect 237300 25566 237328 189314
rect 237380 25628 237432 25634
rect 237380 25570 237432 25576
rect 237288 25560 237340 25566
rect 237288 25502 237340 25508
rect 234620 15972 234672 15978
rect 234620 15914 234672 15920
rect 233148 15904 233200 15910
rect 233148 15846 233200 15852
rect 233240 13116 233292 13122
rect 233240 13058 233292 13064
rect 231768 10328 231820 10334
rect 231768 10270 231820 10276
rect 232504 3596 232556 3602
rect 232504 3538 232556 3544
rect 229112 3454 230152 3482
rect 230492 3454 231348 3482
rect 230124 480 230152 3454
rect 231320 480 231348 3454
rect 232516 480 232544 3538
rect 233252 3482 233280 13058
rect 234632 3482 234660 15914
rect 237196 8968 237248 8974
rect 237196 8910 237248 8916
rect 236000 3528 236052 3534
rect 233252 3454 233740 3482
rect 234632 3454 234844 3482
rect 236000 3470 236052 3476
rect 233712 480 233740 3454
rect 234816 480 234844 3454
rect 236012 480 236040 3470
rect 237208 480 237236 8910
rect 237392 3482 237420 25570
rect 238680 9042 238708 189926
rect 238772 189310 238800 192100
rect 239614 192086 239996 192114
rect 238760 189304 238812 189310
rect 238760 189246 238812 189252
rect 239968 49026 239996 192086
rect 240428 189854 240456 192100
rect 241270 192086 241468 192114
rect 242098 192086 242848 192114
rect 240416 189848 240468 189854
rect 240416 189790 240468 189796
rect 240048 189304 240100 189310
rect 240048 189246 240100 189252
rect 239956 49020 240008 49026
rect 239956 48962 240008 48968
rect 240060 29646 240088 189246
rect 241440 31074 241468 192086
rect 242164 189780 242216 189786
rect 242164 189722 242216 189728
rect 241428 31068 241480 31074
rect 241428 31010 241480 31016
rect 240048 29640 240100 29646
rect 240048 29582 240100 29588
rect 241520 17264 241572 17270
rect 241520 17206 241572 17212
rect 238668 9036 238720 9042
rect 238668 8978 238720 8984
rect 240784 4820 240836 4826
rect 240784 4762 240836 4768
rect 237392 3454 238432 3482
rect 238404 480 238432 3454
rect 239588 3460 239640 3466
rect 239588 3402 239640 3408
rect 239600 480 239628 3402
rect 240796 480 240824 4762
rect 241532 3482 241560 17206
rect 242176 4826 242204 189722
rect 242820 50386 242848 192086
rect 242912 189106 242940 192100
rect 243754 192086 244136 192114
rect 242900 189100 242952 189106
rect 242900 189042 242952 189048
rect 242808 50380 242860 50386
rect 242808 50322 242860 50328
rect 244108 32434 244136 192086
rect 244568 190126 244596 192100
rect 245410 192086 245608 192114
rect 244556 190120 244608 190126
rect 244556 190062 244608 190068
rect 245476 190120 245528 190126
rect 245476 190062 245528 190068
rect 244188 189100 244240 189106
rect 244188 189042 244240 189048
rect 242900 32428 242952 32434
rect 242900 32370 242952 32376
rect 244096 32428 244148 32434
rect 244096 32370 244148 32376
rect 242164 4820 242216 4826
rect 242164 4762 242216 4768
rect 242912 3482 242940 32370
rect 244200 13122 244228 189042
rect 245488 51746 245516 190062
rect 245476 51740 245528 51746
rect 245476 51682 245528 51688
rect 244280 18624 244332 18630
rect 244280 18566 244332 18572
rect 244188 13116 244240 13122
rect 244188 13058 244240 13064
rect 244292 3534 244320 18566
rect 245580 14482 245608 192086
rect 246132 189106 246160 192100
rect 246868 192086 246974 192114
rect 247802 192086 248368 192114
rect 246120 189100 246172 189106
rect 246120 189042 246172 189048
rect 246868 53106 246896 192086
rect 246948 189100 247000 189106
rect 246948 189042 247000 189048
rect 246856 53100 246908 53106
rect 246856 53042 246908 53048
rect 246960 33862 246988 189042
rect 246948 33856 247000 33862
rect 246948 33798 247000 33804
rect 245660 33788 245712 33794
rect 245660 33730 245712 33736
rect 244372 14476 244424 14482
rect 244372 14418 244424 14424
rect 245568 14476 245620 14482
rect 245568 14418 245620 14424
rect 244280 3528 244332 3534
rect 241532 3454 242020 3482
rect 242912 3454 243216 3482
rect 244280 3470 244332 3476
rect 241992 480 242020 3454
rect 243188 480 243216 3454
rect 244384 480 244412 14418
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245672 3482 245700 33730
rect 248340 7614 248368 192086
rect 248616 189310 248644 192100
rect 249458 192086 249656 192114
rect 248604 189304 248656 189310
rect 248604 189246 248656 189252
rect 249628 54534 249656 192086
rect 250272 189514 250300 192100
rect 251008 192086 251114 192114
rect 251942 192086 252508 192114
rect 250260 189508 250312 189514
rect 250260 189450 250312 189456
rect 249708 189304 249760 189310
rect 249708 189246 249760 189252
rect 249616 54528 249668 54534
rect 249616 54470 249668 54476
rect 249720 35222 249748 189246
rect 251008 36582 251036 192086
rect 251088 189508 251140 189514
rect 251088 189450 251140 189456
rect 249800 36576 249852 36582
rect 249800 36518 249852 36524
rect 250996 36576 251048 36582
rect 250996 36518 251048 36524
rect 249708 35216 249760 35222
rect 249708 35158 249760 35164
rect 248420 19984 248472 19990
rect 248420 19926 248472 19932
rect 247960 7608 248012 7614
rect 247960 7550 248012 7556
rect 248328 7608 248380 7614
rect 248328 7550 248380 7556
rect 245580 480 245608 3470
rect 245672 3454 246804 3482
rect 246776 480 246804 3454
rect 247972 480 248000 7550
rect 248432 3482 248460 19926
rect 249812 3482 249840 36518
rect 251100 17338 251128 189450
rect 251180 188352 251232 188358
rect 251180 188294 251232 188300
rect 251088 17332 251140 17338
rect 251088 17274 251140 17280
rect 251192 3482 251220 188294
rect 252480 55894 252508 192086
rect 252756 188358 252784 192100
rect 253584 190126 253612 192100
rect 254426 192086 255176 192114
rect 253572 190120 253624 190126
rect 253572 190062 253624 190068
rect 252744 188352 252796 188358
rect 252744 188294 252796 188300
rect 252560 178696 252612 178702
rect 252560 178638 252612 178644
rect 252468 55888 252520 55894
rect 252468 55830 252520 55836
rect 252572 3534 252600 178638
rect 255148 57254 255176 192086
rect 255136 57248 255188 57254
rect 255136 57190 255188 57196
rect 252652 21412 252704 21418
rect 252652 21354 252704 21360
rect 252560 3528 252612 3534
rect 248432 3454 249196 3482
rect 249812 3454 250392 3482
rect 251192 3454 251496 3482
rect 252560 3470 252612 3476
rect 249168 480 249196 3454
rect 250364 480 250392 3454
rect 251468 480 251496 3454
rect 252664 480 252692 21354
rect 255240 18630 255268 192100
rect 256082 192086 256648 192114
rect 255964 189848 256016 189854
rect 255964 189790 256016 189796
rect 255320 26920 255372 26926
rect 255320 26862 255372 26868
rect 255228 18624 255280 18630
rect 255228 18566 255280 18572
rect 255044 4820 255096 4826
rect 255044 4762 255096 4768
rect 253848 3528 253900 3534
rect 253848 3470 253900 3476
rect 253860 480 253888 3470
rect 255056 480 255084 4762
rect 255332 3618 255360 26862
rect 255976 4826 256004 189790
rect 256620 37942 256648 192086
rect 256896 189106 256924 192100
rect 257344 190120 257396 190126
rect 257344 190062 257396 190068
rect 256884 189100 256936 189106
rect 256884 189042 256936 189048
rect 256700 39364 256752 39370
rect 256700 39306 256752 39312
rect 256608 37936 256660 37942
rect 256608 37878 256660 37884
rect 255964 4820 256016 4826
rect 255964 4762 256016 4768
rect 255332 3590 256280 3618
rect 256252 480 256280 3590
rect 256712 3482 256740 39306
rect 257356 26926 257384 190062
rect 257724 189854 257752 192100
rect 257712 189848 257764 189854
rect 257712 189790 257764 189796
rect 258552 189106 258580 192100
rect 257988 189100 258040 189106
rect 257988 189042 258040 189048
rect 258540 189100 258592 189106
rect 258540 189042 258592 189048
rect 259276 189100 259328 189106
rect 259276 189042 259328 189048
rect 258000 58682 258028 189042
rect 259288 178702 259316 189042
rect 259276 178696 259328 178702
rect 259276 178638 259328 178644
rect 257988 58676 258040 58682
rect 257988 58618 258040 58624
rect 259380 28354 259408 192100
rect 260222 192086 260788 192114
rect 259460 177336 259512 177342
rect 259460 177278 259512 177284
rect 259368 28348 259420 28354
rect 259368 28290 259420 28296
rect 257344 26920 257396 26926
rect 257344 26862 257396 26868
rect 258632 6180 258684 6186
rect 258632 6122 258684 6128
rect 256712 3454 257476 3482
rect 257448 480 257476 3454
rect 258644 480 258672 6122
rect 259472 3482 259500 177278
rect 260760 6186 260788 192086
rect 261036 189378 261064 192100
rect 261878 192086 262076 192114
rect 261024 189372 261076 189378
rect 261024 189314 261076 189320
rect 262048 61402 262076 192086
rect 262128 189372 262180 189378
rect 262128 189314 262180 189320
rect 262036 61396 262088 61402
rect 262036 61338 262088 61344
rect 260840 40724 260892 40730
rect 260840 40666 260892 40672
rect 260748 6180 260800 6186
rect 260748 6122 260800 6128
rect 260852 3482 260880 40666
rect 262140 39438 262168 189314
rect 262692 189106 262720 192100
rect 263428 192086 263534 192114
rect 264362 192086 264928 192114
rect 262680 189100 262732 189106
rect 262680 189042 262732 189048
rect 263428 40730 263456 192086
rect 263508 189100 263560 189106
rect 263508 189042 263560 189048
rect 263416 40724 263468 40730
rect 263416 40666 263468 40672
rect 262128 39432 262180 39438
rect 262128 39374 262180 39380
rect 262220 22772 262272 22778
rect 262220 22714 262272 22720
rect 262232 3602 262260 22714
rect 263520 11762 263548 189042
rect 264900 64190 264928 192086
rect 265176 189310 265204 192100
rect 266018 192086 266216 192114
rect 265164 189304 265216 189310
rect 265164 189246 265216 189252
rect 264888 64184 264940 64190
rect 264888 64126 264940 64132
rect 266188 42158 266216 192086
rect 266268 189304 266320 189310
rect 266268 189246 266320 189252
rect 266176 42152 266228 42158
rect 266176 42094 266228 42100
rect 263600 42084 263652 42090
rect 263600 42026 263652 42032
rect 262312 11756 262364 11762
rect 262312 11698 262364 11704
rect 263508 11756 263560 11762
rect 263508 11698 263560 11704
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 262324 3482 262352 11698
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 259472 3454 259868 3482
rect 260852 3454 261064 3482
rect 259840 480 259868 3454
rect 261036 480 261064 3454
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3538
rect 263612 3482 263640 42026
rect 266280 19990 266308 189246
rect 266832 189106 266860 192100
rect 266820 189100 266872 189106
rect 266820 189042 266872 189048
rect 267556 189100 267608 189106
rect 267556 189042 267608 189048
rect 267568 65550 267596 189042
rect 267556 65544 267608 65550
rect 267556 65486 267608 65492
rect 266360 24132 266412 24138
rect 266360 24074 266412 24080
rect 266268 19984 266320 19990
rect 266268 19926 266320 19932
rect 264980 10328 265032 10334
rect 264980 10270 265032 10276
rect 264992 3482 265020 10270
rect 266372 3482 266400 24074
rect 267660 10334 267688 192100
rect 268502 192086 269068 192114
rect 267740 44872 267792 44878
rect 267740 44814 267792 44820
rect 267648 10328 267700 10334
rect 267648 10270 267700 10276
rect 267752 3482 267780 44814
rect 269040 43450 269068 192086
rect 269224 189990 269252 192100
rect 270066 192086 270448 192114
rect 269212 189984 269264 189990
rect 269212 189926 269264 189932
rect 270316 189984 270368 189990
rect 270316 189926 270368 189932
rect 270328 66910 270356 189926
rect 270316 66904 270368 66910
rect 270316 66846 270368 66852
rect 269028 43444 269080 43450
rect 269028 43386 269080 43392
rect 270420 15910 270448 192086
rect 270880 189310 270908 192100
rect 271722 192086 271828 192114
rect 272550 192086 273208 192114
rect 270868 189304 270920 189310
rect 270868 189246 270920 189252
rect 271800 68338 271828 192086
rect 271972 189304 272024 189310
rect 271972 189246 272024 189252
rect 271984 186998 272012 189246
rect 271880 186992 271932 186998
rect 271880 186934 271932 186940
rect 271972 186992 272024 186998
rect 271972 186934 272024 186940
rect 271788 68332 271840 68338
rect 271788 68274 271840 68280
rect 270500 46232 270552 46238
rect 270500 46174 270552 46180
rect 269120 15904 269172 15910
rect 269120 15846 269172 15852
rect 270408 15904 270460 15910
rect 270408 15846 270460 15852
rect 269132 3482 269160 15846
rect 270512 3602 270540 46174
rect 270592 28280 270644 28286
rect 270592 28222 270644 28228
rect 270500 3596 270552 3602
rect 270500 3538 270552 3544
rect 270604 3482 270632 28222
rect 271696 3596 271748 3602
rect 271696 3538 271748 3544
rect 263612 3454 264652 3482
rect 264992 3454 265848 3482
rect 266372 3454 267044 3482
rect 267752 3454 268148 3482
rect 269132 3454 269344 3482
rect 264624 480 264652 3454
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 268120 480 268148 3454
rect 269316 480 269344 3454
rect 270512 3454 270632 3482
rect 270512 480 270540 3454
rect 271708 480 271736 3538
rect 271892 3482 271920 186934
rect 273180 8974 273208 192086
rect 273364 189106 273392 192100
rect 274206 192086 274496 192114
rect 273352 189100 273404 189106
rect 273352 189042 273404 189048
rect 274468 69698 274496 192086
rect 275020 189786 275048 192100
rect 275862 192086 275968 192114
rect 276690 192086 277348 192114
rect 275008 189780 275060 189786
rect 275008 189722 275060 189728
rect 274548 189100 274600 189106
rect 274548 189042 274600 189048
rect 274456 69692 274508 69698
rect 274456 69634 274508 69640
rect 274560 44946 274588 189042
rect 275940 47598 275968 192086
rect 277320 71058 277348 192086
rect 277504 189378 277532 192100
rect 278346 192086 278636 192114
rect 277492 189372 277544 189378
rect 277492 189314 277544 189320
rect 277308 71052 277360 71058
rect 277308 70994 277360 71000
rect 274640 47592 274692 47598
rect 274640 47534 274692 47540
rect 275928 47592 275980 47598
rect 275928 47534 275980 47540
rect 274548 44940 274600 44946
rect 274548 44882 274600 44888
rect 273260 25560 273312 25566
rect 273260 25502 273312 25508
rect 273168 8968 273220 8974
rect 273168 8910 273220 8916
rect 273272 3482 273300 25502
rect 274652 3482 274680 47534
rect 278608 46238 278636 192086
rect 278688 189372 278740 189378
rect 278688 189314 278740 189320
rect 278596 46232 278648 46238
rect 278596 46174 278648 46180
rect 277400 29640 277452 29646
rect 277400 29582 277452 29588
rect 276480 9036 276532 9042
rect 276480 8978 276532 8984
rect 271892 3454 272932 3482
rect 273272 3454 274128 3482
rect 274652 3454 275324 3482
rect 272904 480 272932 3454
rect 274100 480 274128 3454
rect 275296 480 275324 3454
rect 276492 480 276520 8978
rect 277412 3346 277440 29582
rect 278700 21486 278728 189314
rect 279160 189106 279188 192100
rect 280002 192086 280108 192114
rect 280830 192086 281488 192114
rect 279148 189100 279200 189106
rect 279148 189042 279200 189048
rect 279976 189100 280028 189106
rect 279976 189042 280028 189048
rect 279988 73846 280016 189042
rect 279976 73840 280028 73846
rect 279976 73782 280028 73788
rect 278780 49020 278832 49026
rect 278780 48962 278832 48968
rect 278688 21480 278740 21486
rect 278688 21422 278740 21428
rect 278792 3482 278820 48962
rect 280080 22778 280108 192086
rect 280804 189780 280856 189786
rect 280804 189722 280856 189728
rect 280160 31068 280212 31074
rect 280160 31010 280212 31016
rect 280068 22772 280120 22778
rect 280068 22714 280120 22720
rect 280068 4820 280120 4826
rect 280068 4762 280120 4768
rect 278792 3454 278912 3482
rect 277412 3318 277716 3346
rect 277688 480 277716 3318
rect 278884 480 278912 3454
rect 280080 480 280108 4762
rect 280172 3346 280200 31010
rect 280816 4962 280844 189722
rect 281460 31074 281488 192086
rect 281644 190194 281672 192100
rect 282486 192086 282868 192114
rect 281632 190188 281684 190194
rect 281632 190130 281684 190136
rect 282736 190188 282788 190194
rect 282736 190130 282788 190136
rect 282748 72486 282776 190130
rect 282736 72480 282788 72486
rect 282736 72422 282788 72428
rect 281540 50380 281592 50386
rect 281540 50322 281592 50328
rect 281448 31068 281500 31074
rect 281448 31010 281500 31016
rect 280804 4956 280856 4962
rect 280804 4898 280856 4904
rect 281552 3346 281580 50322
rect 282840 24138 282868 192086
rect 283300 189446 283328 192100
rect 283288 189440 283340 189446
rect 283288 189382 283340 189388
rect 284128 75206 284156 192100
rect 284970 192086 285628 192114
rect 284208 189440 284260 189446
rect 284208 189382 284260 189388
rect 284116 75200 284168 75206
rect 284116 75142 284168 75148
rect 284220 49026 284248 189382
rect 284208 49020 284260 49026
rect 284208 48962 284260 48968
rect 284300 32428 284352 32434
rect 284300 32370 284352 32376
rect 282828 24132 282880 24138
rect 282828 24074 282880 24080
rect 282920 13116 282972 13122
rect 282920 13058 282972 13064
rect 282932 3346 282960 13058
rect 284312 3346 284340 32370
rect 285600 13122 285628 192086
rect 285784 189514 285812 192100
rect 286626 192086 286916 192114
rect 285772 189508 285824 189514
rect 285772 189450 285824 189456
rect 286888 76566 286916 192086
rect 286968 189508 287020 189514
rect 286968 189450 287020 189456
rect 286876 76560 286928 76566
rect 286876 76502 286928 76508
rect 285680 51740 285732 51746
rect 285680 51682 285732 51688
rect 285588 13116 285640 13122
rect 285588 13058 285640 13064
rect 285692 3346 285720 51682
rect 286980 33794 287008 189450
rect 287440 189106 287468 192100
rect 287428 189100 287480 189106
rect 287428 189042 287480 189048
rect 288268 50454 288296 192100
rect 289110 192086 289768 192114
rect 288348 189100 288400 189106
rect 288348 189042 288400 189048
rect 288256 50448 288308 50454
rect 288256 50390 288308 50396
rect 287060 33856 287112 33862
rect 287060 33798 287112 33804
rect 286968 33788 287020 33794
rect 286968 33730 287020 33736
rect 287072 3534 287100 33798
rect 288360 14550 288388 189042
rect 289740 77994 289768 192086
rect 289924 189106 289952 192100
rect 290766 192086 291056 192114
rect 289912 189100 289964 189106
rect 289912 189042 289964 189048
rect 289728 77988 289780 77994
rect 289728 77930 289780 77936
rect 288440 53100 288492 53106
rect 288440 53042 288492 53048
rect 288348 14544 288400 14550
rect 288348 14486 288400 14492
rect 287152 14476 287204 14482
rect 287152 14418 287204 14424
rect 287060 3528 287112 3534
rect 287060 3470 287112 3476
rect 280172 3318 281304 3346
rect 281552 3318 282500 3346
rect 282932 3318 283696 3346
rect 284312 3318 284800 3346
rect 285692 3318 285996 3346
rect 281276 480 281304 3318
rect 282472 480 282500 3318
rect 283668 480 283696 3318
rect 284772 480 284800 3318
rect 285968 480 285996 3318
rect 287164 480 287192 14418
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288452 3482 288480 53042
rect 291028 51814 291056 192086
rect 291580 189106 291608 192100
rect 292330 192086 292528 192114
rect 291108 189100 291160 189106
rect 291108 189042 291160 189048
rect 291568 189100 291620 189106
rect 291568 189042 291620 189048
rect 292396 189100 292448 189106
rect 292396 189042 292448 189048
rect 291016 51808 291068 51814
rect 291016 51750 291068 51756
rect 291120 7614 291148 189042
rect 292408 79354 292436 189042
rect 292396 79348 292448 79354
rect 292396 79290 292448 79296
rect 291200 35216 291252 35222
rect 291200 35158 291252 35164
rect 290740 7608 290792 7614
rect 290740 7550 290792 7556
rect 291108 7608 291160 7614
rect 291108 7550 291160 7556
rect 288360 480 288388 3470
rect 288452 3454 289584 3482
rect 289556 480 289584 3454
rect 290752 480 290780 7550
rect 291212 3482 291240 35158
rect 292500 17270 292528 192086
rect 293144 189106 293172 192100
rect 293972 189446 294000 192100
rect 294800 189786 294828 192100
rect 294788 189780 294840 189786
rect 294788 189722 294840 189728
rect 293960 189440 294012 189446
rect 293960 189382 294012 189388
rect 295248 189440 295300 189446
rect 295248 189382 295300 189388
rect 293132 189100 293184 189106
rect 293132 189042 293184 189048
rect 293868 189100 293920 189106
rect 293868 189042 293920 189048
rect 292580 54528 292632 54534
rect 292580 54470 292632 54476
rect 292488 17264 292540 17270
rect 292488 17206 292540 17212
rect 292592 3482 292620 54470
rect 293880 53106 293908 189042
rect 295260 80714 295288 189382
rect 295628 189106 295656 192100
rect 296470 192086 296576 192114
rect 297298 192086 298048 192114
rect 295616 189100 295668 189106
rect 295616 189042 295668 189048
rect 295248 80708 295300 80714
rect 295248 80650 295300 80656
rect 293868 53100 293920 53106
rect 293868 53042 293920 53048
rect 296548 39370 296576 192086
rect 296628 189100 296680 189106
rect 296628 189042 296680 189048
rect 296536 39364 296588 39370
rect 296536 39306 296588 39312
rect 296640 36650 296668 189042
rect 296720 188352 296772 188358
rect 296720 188294 296772 188300
rect 296628 36644 296680 36650
rect 296628 36586 296680 36592
rect 295340 36576 295392 36582
rect 295340 36518 295392 36524
rect 293960 17332 294012 17338
rect 293960 17274 294012 17280
rect 293972 3482 294000 17274
rect 295352 3482 295380 36518
rect 296732 3534 296760 188294
rect 296812 55888 296864 55894
rect 296812 55830 296864 55836
rect 296720 3528 296772 3534
rect 291212 3454 291976 3482
rect 292592 3454 293172 3482
rect 293972 3454 294368 3482
rect 295352 3454 295564 3482
rect 296720 3470 296772 3476
rect 291948 480 291976 3454
rect 293144 480 293172 3454
rect 294340 480 294368 3454
rect 295536 480 295564 3454
rect 296824 1442 296852 55830
rect 298020 25566 298048 192086
rect 298112 189106 298140 192100
rect 298954 192086 299336 192114
rect 298100 189100 298152 189106
rect 298100 189042 298152 189048
rect 299308 82142 299336 192086
rect 299768 189378 299796 192100
rect 300610 192086 300716 192114
rect 299756 189372 299808 189378
rect 299756 189314 299808 189320
rect 299388 189100 299440 189106
rect 299388 189042 299440 189048
rect 299296 82136 299348 82142
rect 299296 82078 299348 82084
rect 299400 54534 299428 189042
rect 299480 57248 299532 57254
rect 299480 57190 299532 57196
rect 299388 54528 299440 54534
rect 299388 54470 299440 54476
rect 298100 26920 298152 26926
rect 298100 26862 298152 26868
rect 298008 25560 298060 25566
rect 298008 25502 298060 25508
rect 297916 3528 297968 3534
rect 297916 3470 297968 3476
rect 298112 3482 298140 26862
rect 299492 3482 299520 57190
rect 300688 55894 300716 192086
rect 300768 189372 300820 189378
rect 300768 189314 300820 189320
rect 300676 55888 300728 55894
rect 300676 55830 300728 55836
rect 300780 26926 300808 189314
rect 301424 189106 301452 192100
rect 301504 189848 301556 189854
rect 301504 189790 301556 189796
rect 301412 189100 301464 189106
rect 301412 189042 301464 189048
rect 300768 26920 300820 26926
rect 300768 26862 300820 26868
rect 301516 19310 301544 189790
rect 302252 189310 302280 192100
rect 303094 192086 303476 192114
rect 302240 189304 302292 189310
rect 302240 189246 302292 189252
rect 302148 189100 302200 189106
rect 302148 189042 302200 189048
rect 302160 83502 302188 189042
rect 302148 83496 302200 83502
rect 302148 83438 302200 83444
rect 303448 57254 303476 192086
rect 303908 190398 303936 192100
rect 304750 192086 304948 192114
rect 305578 192086 306328 192114
rect 303896 190392 303948 190398
rect 303896 190334 303948 190340
rect 304816 190392 304868 190398
rect 304816 190334 304868 190340
rect 303528 189304 303580 189310
rect 303528 189246 303580 189252
rect 303436 57248 303488 57254
rect 303436 57190 303488 57196
rect 302240 37936 302292 37942
rect 302240 37878 302292 37884
rect 301504 19304 301556 19310
rect 301504 19246 301556 19252
rect 300860 18624 300912 18630
rect 300860 18566 300912 18572
rect 300872 3482 300900 18566
rect 302252 3482 302280 37878
rect 303540 28286 303568 189246
rect 304828 86290 304856 190334
rect 304816 86284 304868 86290
rect 304816 86226 304868 86232
rect 303620 58676 303672 58682
rect 303620 58618 303672 58624
rect 303528 28280 303580 28286
rect 303528 28222 303580 28228
rect 303632 3482 303660 58618
rect 304920 29646 304948 192086
rect 305000 178696 305052 178702
rect 305000 178638 305052 178644
rect 304908 29640 304960 29646
rect 304908 29582 304960 29588
rect 305012 3534 305040 178638
rect 306300 58682 306328 192086
rect 306392 189310 306420 192100
rect 306380 189304 306432 189310
rect 306380 189246 306432 189252
rect 307220 189174 307248 192100
rect 307668 189304 307720 189310
rect 307668 189246 307720 189252
rect 307208 189168 307260 189174
rect 307208 189110 307260 189116
rect 307680 84862 307708 189246
rect 308048 189106 308076 192100
rect 308890 192086 309088 192114
rect 308036 189100 308088 189106
rect 308036 189042 308088 189048
rect 308956 189100 309008 189106
rect 308956 189042 309008 189048
rect 307668 84856 307720 84862
rect 307668 84798 307720 84804
rect 308968 60042 308996 189042
rect 308956 60036 309008 60042
rect 308956 59978 309008 59984
rect 306288 58676 306340 58682
rect 306288 58618 306340 58624
rect 306380 28348 306432 28354
rect 306380 28290 306432 28296
rect 305092 19304 305144 19310
rect 305092 19246 305144 19252
rect 305000 3528 305052 3534
rect 296732 1414 296852 1442
rect 296732 480 296760 1414
rect 297928 480 297956 3470
rect 298112 3454 299152 3482
rect 299492 3454 300348 3482
rect 300872 3454 301452 3482
rect 302252 3454 302648 3482
rect 303632 3454 303844 3482
rect 305000 3470 305052 3476
rect 299124 480 299152 3454
rect 300320 480 300348 3454
rect 301424 480 301452 3454
rect 302620 480 302648 3454
rect 303816 480 303844 3454
rect 305104 1442 305132 19246
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 305012 1414 305132 1442
rect 305012 480 305040 1414
rect 306208 480 306236 3470
rect 306392 3346 306420 28290
rect 308588 6180 308640 6186
rect 308588 6122 308640 6128
rect 306392 3318 307432 3346
rect 307404 480 307432 3318
rect 308600 480 308628 6122
rect 309060 4826 309088 192086
rect 309704 189718 309732 192100
rect 310532 189922 310560 192100
rect 311374 192086 311848 192114
rect 310520 189916 310572 189922
rect 310520 189858 310572 189864
rect 309692 189712 309744 189718
rect 309692 189654 309744 189660
rect 310428 189712 310480 189718
rect 310428 189654 310480 189660
rect 309784 189168 309836 189174
rect 309784 189110 309836 189116
rect 309140 39432 309192 39438
rect 309140 39374 309192 39380
rect 309048 4820 309100 4826
rect 309048 4762 309100 4768
rect 309152 3346 309180 39374
rect 309796 6186 309824 189110
rect 310440 18630 310468 189654
rect 311820 89010 311848 192086
rect 312188 189310 312216 192100
rect 313030 192086 313136 192114
rect 313858 192086 314516 192114
rect 312176 189304 312228 189310
rect 312176 189246 312228 189252
rect 311808 89004 311860 89010
rect 311808 88946 311860 88952
rect 313108 62830 313136 192086
rect 313188 189304 313240 189310
rect 313188 189246 313240 189252
rect 313096 62824 313148 62830
rect 313096 62766 313148 62772
rect 310520 61396 310572 61402
rect 310520 61338 310572 61344
rect 310428 18624 310480 18630
rect 310428 18566 310480 18572
rect 309784 6180 309836 6186
rect 309784 6122 309836 6128
rect 310532 3346 310560 61338
rect 313200 11762 313228 189246
rect 314488 91798 314516 192086
rect 314476 91792 314528 91798
rect 314476 91734 314528 91740
rect 313280 64184 313332 64190
rect 313280 64126 313332 64132
rect 311900 11756 311952 11762
rect 311900 11698 311952 11704
rect 313188 11756 313240 11762
rect 313188 11698 313240 11704
rect 311912 3346 311940 11698
rect 313292 3534 313320 64126
rect 313372 40724 313424 40730
rect 313372 40666 313424 40672
rect 313280 3528 313332 3534
rect 313280 3470 313332 3476
rect 309152 3318 309824 3346
rect 310532 3318 311020 3346
rect 311912 3318 312216 3346
rect 309796 480 309824 3318
rect 310992 480 311020 3318
rect 312188 480 312216 3318
rect 313384 480 313412 40666
rect 314580 32434 314608 192100
rect 315422 192086 315988 192114
rect 315304 189916 315356 189922
rect 315304 189858 315356 189864
rect 315316 61402 315344 189858
rect 315304 61396 315356 61402
rect 315304 61338 315356 61344
rect 315960 42090 315988 192086
rect 316236 190126 316264 192100
rect 317078 192086 317368 192114
rect 317906 192086 318656 192114
rect 316224 190120 316276 190126
rect 316224 190062 316276 190068
rect 317236 190120 317288 190126
rect 317236 190062 317288 190068
rect 317248 93158 317276 190062
rect 317236 93152 317288 93158
rect 317236 93094 317288 93100
rect 316040 42152 316092 42158
rect 316040 42094 316092 42100
rect 315948 42084 316000 42090
rect 315948 42026 316000 42032
rect 314568 32428 314620 32434
rect 314568 32370 314620 32376
rect 314660 19984 314712 19990
rect 314660 19926 314712 19932
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 314580 480 314608 3470
rect 314672 3346 314700 19926
rect 316052 3482 316080 42094
rect 317340 35222 317368 192086
rect 318628 178702 318656 192086
rect 318616 178696 318668 178702
rect 318616 178638 318668 178644
rect 318720 94518 318748 192100
rect 319562 192086 320128 192114
rect 318708 94512 318760 94518
rect 318708 94454 318760 94460
rect 317420 65544 317472 65550
rect 317420 65486 317472 65492
rect 317328 35216 317380 35222
rect 317328 35158 317380 35164
rect 317432 3482 317460 65486
rect 320100 10334 320128 192086
rect 320376 189310 320404 192100
rect 321218 192086 321416 192114
rect 320364 189304 320416 189310
rect 320364 189246 320416 189252
rect 321388 95946 321416 192086
rect 322032 189514 322060 192100
rect 322768 192086 322874 192114
rect 323702 192086 324268 192114
rect 322020 189508 322072 189514
rect 322020 189450 322072 189456
rect 321468 189304 321520 189310
rect 321468 189246 321520 189252
rect 321376 95940 321428 95946
rect 321376 95882 321428 95888
rect 321480 64190 321508 189246
rect 321560 66904 321612 66910
rect 321560 66846 321612 66852
rect 321468 64184 321520 64190
rect 321468 64126 321520 64132
rect 320180 43444 320232 43450
rect 320180 43386 320232 43392
rect 318800 10328 318852 10334
rect 318800 10270 318852 10276
rect 320088 10328 320140 10334
rect 320088 10270 320140 10276
rect 318812 3482 318840 10270
rect 320192 3482 320220 43386
rect 321572 3482 321600 66846
rect 322768 65550 322796 192086
rect 322848 189508 322900 189514
rect 322848 189450 322900 189456
rect 322756 65544 322808 65550
rect 322756 65486 322808 65492
rect 322860 15910 322888 189450
rect 322940 186992 322992 186998
rect 322940 186934 322992 186940
rect 321652 15904 321704 15910
rect 321652 15846 321704 15852
rect 322848 15904 322900 15910
rect 322848 15846 322900 15852
rect 321664 3602 321692 15846
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 316052 3454 317000 3482
rect 317432 3454 318104 3482
rect 318812 3454 319300 3482
rect 320192 3454 320496 3482
rect 321572 3454 321692 3482
rect 314672 3318 315804 3346
rect 315776 480 315804 3318
rect 316972 480 317000 3454
rect 318076 480 318104 3454
rect 319272 480 319300 3454
rect 320468 480 320496 3454
rect 321664 480 321692 3454
rect 322860 480 322888 3538
rect 322952 3482 322980 186934
rect 324240 97306 324268 192086
rect 324516 189106 324544 192100
rect 325358 192086 325648 192114
rect 326186 192086 326936 192114
rect 324504 189100 324556 189106
rect 324504 189042 324556 189048
rect 324228 97300 324280 97306
rect 324228 97242 324280 97248
rect 324320 68332 324372 68338
rect 324320 68274 324372 68280
rect 324332 3482 324360 68274
rect 325620 44878 325648 192086
rect 326908 98666 326936 192086
rect 326896 98660 326948 98666
rect 326896 98602 326948 98608
rect 325608 44872 325660 44878
rect 325608 44814 325660 44820
rect 327000 19990 327028 192100
rect 327842 192086 328408 192114
rect 327724 189100 327776 189106
rect 327724 189042 327776 189048
rect 327080 44940 327132 44946
rect 327080 44882 327132 44888
rect 326988 19984 327040 19990
rect 326988 19926 327040 19932
rect 326436 8968 326488 8974
rect 326436 8910 326488 8916
rect 322952 3454 324084 3482
rect 324332 3454 325280 3482
rect 324056 480 324084 3454
rect 325252 480 325280 3454
rect 326448 480 326476 8910
rect 327092 3482 327120 44882
rect 327736 8974 327764 189042
rect 328380 90370 328408 192086
rect 328656 189446 328684 192100
rect 329484 189990 329512 192100
rect 329472 189984 329524 189990
rect 329472 189926 329524 189932
rect 330312 189514 330340 192100
rect 331048 192086 331154 192114
rect 331982 192086 332548 192114
rect 330300 189508 330352 189514
rect 330300 189450 330352 189456
rect 328644 189440 328696 189446
rect 328644 189382 328696 189388
rect 329748 189440 329800 189446
rect 329748 189382 329800 189388
rect 329760 100026 329788 189382
rect 331048 108322 331076 192086
rect 331864 189984 331916 189990
rect 331864 189926 331916 189932
rect 331128 189508 331180 189514
rect 331128 189450 331180 189456
rect 331036 108316 331088 108322
rect 331036 108258 331088 108264
rect 329748 100020 329800 100026
rect 329748 99962 329800 99968
rect 328368 90364 328420 90370
rect 328368 90306 328420 90312
rect 328460 69692 328512 69698
rect 328460 69634 328512 69640
rect 327724 8968 327776 8974
rect 327724 8910 327776 8916
rect 328472 3482 328500 69634
rect 331140 47666 331168 189450
rect 331876 104174 331904 189926
rect 331864 104168 331916 104174
rect 331864 104110 331916 104116
rect 331220 71052 331272 71058
rect 331220 70994 331272 71000
rect 331128 47660 331180 47666
rect 331128 47602 331180 47608
rect 330024 4888 330076 4894
rect 330024 4830 330076 4836
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330036 480 330064 4830
rect 331232 3602 331260 70994
rect 331312 47592 331364 47598
rect 331312 47534 331364 47540
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 331324 3482 331352 47534
rect 332520 21418 332548 192086
rect 332796 190262 332824 192100
rect 333638 192086 333836 192114
rect 334466 192086 335216 192114
rect 332784 190256 332836 190262
rect 332784 190198 332836 190204
rect 333808 109750 333836 192086
rect 333888 190256 333940 190262
rect 333888 190198 333940 190204
rect 333796 109744 333848 109750
rect 333796 109686 333848 109692
rect 333900 66910 333928 190198
rect 335188 177342 335216 192086
rect 335176 177336 335228 177342
rect 335176 177278 335228 177284
rect 335280 68338 335308 192100
rect 336122 192086 336688 192114
rect 336660 101454 336688 192086
rect 336936 189310 336964 192100
rect 337686 192086 337976 192114
rect 336924 189304 336976 189310
rect 336924 189246 336976 189252
rect 336648 101448 336700 101454
rect 336648 101390 336700 101396
rect 335360 73840 335412 73846
rect 335360 73782 335412 73788
rect 335268 68332 335320 68338
rect 335268 68274 335320 68280
rect 333888 66904 333940 66910
rect 333888 66846 333940 66852
rect 333980 46232 334032 46238
rect 333980 46174 334032 46180
rect 332600 21480 332652 21486
rect 332600 21422 332652 21428
rect 332508 21412 332560 21418
rect 332508 21354 332560 21360
rect 332416 3596 332468 3602
rect 332416 3538 332468 3544
rect 331232 3454 331352 3482
rect 331232 480 331260 3454
rect 332428 480 332456 3538
rect 332612 3482 332640 21422
rect 333992 3482 334020 46174
rect 335372 3482 335400 73782
rect 337948 69698 337976 192086
rect 338028 189304 338080 189310
rect 338028 189246 338080 189252
rect 337936 69692 337988 69698
rect 337936 69634 337988 69640
rect 338040 22778 338068 189246
rect 338500 189106 338528 192100
rect 339342 192086 339448 192114
rect 340170 192086 340828 192114
rect 338488 189100 338540 189106
rect 338488 189042 338540 189048
rect 339316 189100 339368 189106
rect 339316 189042 339368 189048
rect 339328 102814 339356 189042
rect 339316 102808 339368 102814
rect 339316 102750 339368 102756
rect 338120 31068 338172 31074
rect 338120 31010 338172 31016
rect 336740 22772 336792 22778
rect 336740 22714 336792 22720
rect 338028 22772 338080 22778
rect 338028 22714 338080 22720
rect 336752 3482 336780 22714
rect 338132 3482 338160 31010
rect 339420 24206 339448 192086
rect 339500 72480 339552 72486
rect 339500 72422 339552 72428
rect 339408 24200 339460 24206
rect 339408 24142 339460 24148
rect 332612 3454 333652 3482
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 333624 480 333652 3454
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339512 480 339540 72422
rect 340800 71058 340828 192086
rect 340984 189990 341012 192100
rect 341826 192086 342208 192114
rect 340972 189984 341024 189990
rect 340972 189926 341024 189932
rect 342076 189984 342128 189990
rect 342076 189926 342128 189932
rect 342088 106962 342116 189926
rect 342076 106956 342128 106962
rect 342076 106898 342128 106904
rect 340788 71052 340840 71058
rect 340788 70994 340840 71000
rect 340880 49020 340932 49026
rect 340880 48962 340932 48968
rect 339592 24132 339644 24138
rect 339592 24074 339644 24080
rect 339604 3482 339632 24074
rect 340892 3482 340920 48962
rect 342180 37942 342208 192086
rect 342640 189106 342668 192100
rect 343482 192086 343588 192114
rect 344310 192086 344968 192114
rect 342628 189100 342680 189106
rect 342628 189042 342680 189048
rect 343560 112470 343588 192086
rect 344284 189100 344336 189106
rect 344284 189042 344336 189048
rect 343548 112464 343600 112470
rect 343548 112406 343600 112412
rect 342260 75200 342312 75206
rect 342260 75142 342312 75148
rect 342168 37936 342220 37942
rect 342168 37878 342220 37884
rect 342272 3482 342300 75142
rect 344296 72486 344324 189042
rect 344284 72480 344336 72486
rect 344284 72422 344336 72428
rect 344940 14482 344968 192086
rect 345124 190126 345152 192100
rect 345966 192086 346348 192114
rect 345112 190120 345164 190126
rect 345112 190062 345164 190068
rect 346216 190120 346268 190126
rect 346216 190062 346268 190068
rect 346228 73846 346256 190062
rect 346216 73840 346268 73846
rect 346216 73782 346268 73788
rect 346320 50386 346348 192086
rect 346780 189106 346808 192100
rect 347622 192086 347728 192114
rect 348450 192086 349108 192114
rect 346768 189100 346820 189106
rect 346768 189042 346820 189048
rect 346400 76560 346452 76566
rect 346400 76502 346452 76508
rect 346308 50380 346360 50386
rect 346308 50322 346360 50328
rect 345020 33788 345072 33794
rect 345020 33730 345072 33736
rect 344928 14476 344980 14482
rect 344928 14418 344980 14424
rect 343640 13116 343692 13122
rect 343640 13058 343692 13064
rect 343652 3482 343680 13058
rect 345032 3482 345060 33730
rect 346412 3482 346440 76502
rect 347700 75206 347728 192086
rect 348424 189100 348476 189106
rect 348424 189042 348476 189048
rect 347688 75200 347740 75206
rect 347688 75142 347740 75148
rect 347780 50448 347832 50454
rect 347780 50390 347832 50396
rect 347792 3534 347820 50390
rect 348436 31074 348464 189042
rect 349080 105602 349108 192086
rect 349264 189854 349292 192100
rect 350106 192086 350488 192114
rect 349252 189848 349304 189854
rect 349252 189790 349304 189796
rect 349068 105596 349120 105602
rect 349068 105538 349120 105544
rect 349160 77988 349212 77994
rect 349160 77930 349212 77936
rect 348424 31068 348476 31074
rect 348424 31010 348476 31016
rect 347872 14544 347924 14550
rect 347872 14486 347924 14492
rect 347780 3528 347832 3534
rect 339604 3454 340736 3482
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 343652 3454 344324 3482
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 347780 3470 347832 3476
rect 340708 480 340736 3454
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 3454
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 14486
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 349172 3482 349200 77930
rect 350460 51746 350488 192086
rect 350920 189106 350948 192100
rect 351762 192086 351868 192114
rect 352590 192086 353248 192114
rect 350908 189100 350960 189106
rect 350908 189042 350960 189048
rect 351736 189100 351788 189106
rect 351736 189042 351788 189048
rect 351748 113830 351776 189042
rect 351736 113824 351788 113830
rect 351736 113766 351788 113772
rect 350448 51740 350500 51746
rect 350448 51682 350500 51688
rect 351840 33794 351868 192086
rect 352564 189780 352616 189786
rect 352564 189722 352616 189728
rect 351920 51808 351972 51814
rect 351920 51750 351972 51756
rect 351828 33788 351880 33794
rect 351828 33730 351880 33736
rect 351368 7608 351420 7614
rect 351368 7550 351420 7556
rect 349080 480 349108 3470
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 7550
rect 351932 3618 351960 51750
rect 352576 4894 352604 189722
rect 353220 76566 353248 192086
rect 353404 190126 353432 192100
rect 354246 192086 354628 192114
rect 353392 190120 353444 190126
rect 353392 190062 353444 190068
rect 354496 190120 354548 190126
rect 354496 190062 354548 190068
rect 354508 166326 354536 190062
rect 354496 166320 354548 166326
rect 354496 166262 354548 166268
rect 353300 79348 353352 79354
rect 353300 79290 353352 79296
rect 353208 76560 353260 76566
rect 353208 76502 353260 76508
rect 352564 4888 352616 4894
rect 352564 4830 352616 4836
rect 351932 3590 352604 3618
rect 352576 480 352604 3590
rect 353312 3482 353340 79290
rect 354600 40730 354628 192086
rect 355060 189106 355088 192100
rect 355902 192086 356008 192114
rect 356730 192086 357388 192114
rect 355048 189100 355100 189106
rect 355048 189042 355100 189048
rect 355876 189100 355928 189106
rect 355876 189042 355928 189048
rect 355888 79354 355916 189042
rect 355876 79348 355928 79354
rect 355876 79290 355928 79296
rect 354588 40724 354640 40730
rect 354588 40666 354640 40672
rect 354680 17264 354732 17270
rect 354680 17206 354732 17212
rect 353312 3454 353800 3482
rect 353772 480 353800 3454
rect 354692 3346 354720 17206
rect 355980 3466 356008 192086
rect 356060 80708 356112 80714
rect 356060 80650 356112 80656
rect 356072 3534 356100 80650
rect 356152 53100 356204 53106
rect 356152 53042 356204 53048
rect 356060 3528 356112 3534
rect 356060 3470 356112 3476
rect 355968 3460 356020 3466
rect 355968 3402 356020 3408
rect 354692 3318 354996 3346
rect 354968 480 354996 3318
rect 356164 480 356192 53042
rect 357360 36582 357388 192086
rect 357544 189990 357572 192100
rect 358386 192086 358768 192114
rect 357532 189984 357584 189990
rect 357532 189926 357584 189932
rect 358636 189984 358688 189990
rect 358636 189926 358688 189932
rect 358648 53106 358676 189926
rect 358636 53100 358688 53106
rect 358636 53042 358688 53048
rect 357348 36576 357400 36582
rect 357348 36518 357400 36524
rect 358544 4888 358596 4894
rect 358544 4830 358596 4836
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 357360 480 357388 3470
rect 358556 480 358584 4830
rect 358740 3466 358768 192086
rect 359200 189106 359228 192100
rect 359950 192086 360056 192114
rect 360778 192086 361528 192114
rect 359188 189100 359240 189106
rect 359188 189042 359240 189048
rect 360028 77994 360056 192086
rect 360108 189100 360160 189106
rect 360108 189042 360160 189048
rect 360016 77988 360068 77994
rect 360016 77930 360068 77936
rect 360120 43450 360148 189042
rect 360108 43444 360160 43450
rect 360108 43386 360160 43392
rect 360200 39364 360252 39370
rect 360200 39306 360252 39312
rect 358820 36644 358872 36650
rect 358820 36586 358872 36592
rect 358728 3460 358780 3466
rect 358728 3402 358780 3408
rect 358832 3346 358860 36586
rect 360212 3346 360240 39306
rect 361500 4146 361528 192086
rect 361592 189106 361620 192100
rect 362434 192086 362816 192114
rect 361580 189100 361632 189106
rect 361580 189042 361632 189048
rect 362788 80714 362816 192086
rect 363248 189106 363276 192100
rect 364090 192086 364196 192114
rect 362868 189100 362920 189106
rect 362868 189042 362920 189048
rect 363236 189100 363288 189106
rect 363236 189042 363288 189048
rect 362776 80708 362828 80714
rect 362776 80650 362828 80656
rect 362880 39370 362908 189042
rect 364168 163538 364196 192086
rect 364904 189106 364932 192100
rect 365732 189310 365760 192100
rect 366574 192086 366956 192114
rect 365720 189304 365772 189310
rect 365720 189246 365772 189252
rect 364248 189100 364300 189106
rect 364248 189042 364300 189048
rect 364892 189100 364944 189106
rect 364892 189042 364944 189048
rect 365628 189100 365680 189106
rect 365628 189042 365680 189048
rect 364156 163532 364208 163538
rect 364156 163474 364208 163480
rect 362960 54528 363012 54534
rect 362960 54470 363012 54476
rect 362868 39364 362920 39370
rect 362868 39306 362920 39312
rect 361580 25560 361632 25566
rect 361580 25502 361632 25508
rect 361488 4140 361540 4146
rect 361488 4082 361540 4088
rect 361592 3346 361620 25502
rect 362972 3346 363000 54470
rect 364260 4078 364288 189042
rect 365640 158030 365668 189042
rect 366928 162178 366956 192086
rect 367008 189304 367060 189310
rect 367008 189246 367060 189252
rect 366916 162172 366968 162178
rect 366916 162114 366968 162120
rect 365628 158024 365680 158030
rect 365628 157966 365680 157972
rect 364340 82136 364392 82142
rect 364340 82078 364392 82084
rect 364248 4072 364300 4078
rect 364248 4014 364300 4020
rect 358832 3318 359780 3346
rect 360212 3318 360976 3346
rect 361592 3318 362172 3346
rect 362972 3318 363368 3346
rect 359752 480 359780 3318
rect 360948 480 360976 3318
rect 362144 480 362172 3318
rect 363340 480 363368 3318
rect 364352 610 364380 82078
rect 365720 55888 365772 55894
rect 365720 55830 365772 55836
rect 365732 3602 365760 55830
rect 365812 26920 365864 26926
rect 365812 26862 365864 26868
rect 365720 3596 365772 3602
rect 365720 3538 365772 3544
rect 365824 3482 365852 26862
rect 367020 4010 367048 189246
rect 367388 181490 367416 192100
rect 368230 192086 368428 192114
rect 369058 192086 369808 192114
rect 367376 181484 367428 181490
rect 367376 181426 367428 181432
rect 367100 83496 367152 83502
rect 367100 83438 367152 83444
rect 367008 4004 367060 4010
rect 367008 3946 367060 3952
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 365732 3454 365852 3482
rect 364340 604 364392 610
rect 364340 546 364392 552
rect 364524 604 364576 610
rect 364524 546 364576 552
rect 364536 480 364564 546
rect 365732 480 365760 3454
rect 366928 480 366956 3538
rect 367112 610 367140 83438
rect 368400 3942 368428 192086
rect 369780 28286 369808 192086
rect 369872 190058 369900 192100
rect 370714 192086 371188 192114
rect 369860 190052 369912 190058
rect 369860 189994 369912 190000
rect 371056 190052 371108 190058
rect 371056 189994 371108 190000
rect 371068 140078 371096 189994
rect 371056 140072 371108 140078
rect 371056 140014 371108 140020
rect 369860 57248 369912 57254
rect 369860 57190 369912 57196
rect 368480 28280 368532 28286
rect 368480 28222 368532 28228
rect 369768 28280 369820 28286
rect 369768 28222 369820 28228
rect 368388 3936 368440 3942
rect 368388 3878 368440 3884
rect 368492 610 368520 28222
rect 369872 610 369900 57190
rect 371160 3806 371188 192086
rect 371528 189378 371556 192100
rect 372370 192086 372476 192114
rect 371516 189372 371568 189378
rect 371516 189314 371568 189320
rect 372448 111110 372476 192086
rect 373184 189990 373212 192100
rect 373172 189984 373224 189990
rect 373172 189926 373224 189932
rect 373908 189984 373960 189990
rect 373908 189926 373960 189932
rect 372528 189372 372580 189378
rect 372528 189314 372580 189320
rect 372436 111104 372488 111110
rect 372436 111046 372488 111052
rect 371240 86284 371292 86290
rect 371240 86226 371292 86232
rect 371148 3800 371200 3806
rect 371148 3742 371200 3748
rect 371252 626 371280 86226
rect 372540 26926 372568 189314
rect 372620 29640 372672 29646
rect 372620 29582 372672 29588
rect 372528 26920 372580 26926
rect 372528 26862 372580 26868
rect 367100 604 367152 610
rect 367100 546 367152 552
rect 368020 604 368072 610
rect 368020 546 368072 552
rect 368480 604 368532 610
rect 368480 546 368532 552
rect 369216 604 369268 610
rect 369216 546 369268 552
rect 369860 604 369912 610
rect 369860 546 369912 552
rect 370412 604 370464 610
rect 371252 598 371648 626
rect 372632 610 372660 29582
rect 373920 3874 373948 189926
rect 374012 189310 374040 192100
rect 374854 192086 375236 192114
rect 374000 189304 374052 189310
rect 374000 189246 374052 189252
rect 375208 87650 375236 192086
rect 375668 190262 375696 192100
rect 376510 192086 376616 192114
rect 377338 192086 378088 192114
rect 375656 190256 375708 190262
rect 375656 190198 375708 190204
rect 375288 189304 375340 189310
rect 375288 189246 375340 189252
rect 375196 87644 375248 87650
rect 375196 87586 375248 87592
rect 374000 84856 374052 84862
rect 374000 84798 374052 84804
rect 373908 3868 373960 3874
rect 373908 3810 373960 3816
rect 374012 3602 374040 84798
rect 374092 58676 374144 58682
rect 374092 58618 374144 58624
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 374104 3482 374132 58618
rect 375300 46238 375328 189246
rect 376588 160750 376616 192086
rect 376668 190256 376720 190262
rect 376668 190198 376720 190204
rect 376576 160744 376628 160750
rect 376576 160686 376628 160692
rect 375288 46232 375340 46238
rect 375288 46174 375340 46180
rect 376392 6180 376444 6186
rect 376392 6122 376444 6128
rect 375196 3596 375248 3602
rect 375196 3538 375248 3544
rect 374012 3454 374132 3482
rect 370412 546 370464 552
rect 368032 480 368060 546
rect 369228 480 369256 546
rect 370424 480 370452 546
rect 371620 480 371648 598
rect 372620 604 372672 610
rect 372620 546 372672 552
rect 372804 604 372856 610
rect 372804 546 372856 552
rect 372816 480 372844 546
rect 374012 480 374040 3454
rect 375208 480 375236 3538
rect 376404 480 376432 6122
rect 376680 3670 376708 190198
rect 376760 60036 376812 60042
rect 376760 59978 376812 59984
rect 376668 3664 376720 3670
rect 376668 3606 376720 3612
rect 376772 610 376800 59978
rect 378060 54534 378088 192086
rect 378152 189310 378180 192100
rect 378140 189304 378192 189310
rect 378140 189246 378192 189252
rect 378980 189174 379008 192100
rect 379428 189304 379480 189310
rect 379428 189246 379480 189252
rect 378968 189168 379020 189174
rect 378968 189110 379020 189116
rect 378048 54528 378100 54534
rect 378048 54470 378100 54476
rect 378784 4820 378836 4826
rect 378784 4762 378836 4768
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 377600 480 377628 546
rect 378796 480 378824 4762
rect 379440 3738 379468 189246
rect 379808 189106 379836 192100
rect 380650 192086 380848 192114
rect 379796 189100 379848 189106
rect 379796 189042 379848 189048
rect 380716 189100 380768 189106
rect 380716 189042 380768 189048
rect 380728 138718 380756 189042
rect 380716 138712 380768 138718
rect 380716 138654 380768 138660
rect 379520 18624 379572 18630
rect 379520 18566 379572 18572
rect 379428 3732 379480 3738
rect 379428 3674 379480 3680
rect 379532 610 379560 18566
rect 380820 3602 380848 192086
rect 381464 189106 381492 192100
rect 382292 189922 382320 192100
rect 383042 192086 383608 192114
rect 382280 189916 382332 189922
rect 382280 189858 382332 189864
rect 381544 189168 381596 189174
rect 381544 189110 381596 189116
rect 381452 189100 381504 189106
rect 381452 189042 381504 189048
rect 381556 159390 381584 189110
rect 382188 189100 382240 189106
rect 382188 189042 382240 189048
rect 381544 159384 381596 159390
rect 381544 159326 381596 159332
rect 380900 61396 380952 61402
rect 380900 61338 380952 61344
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 380912 626 380940 61338
rect 382200 4826 382228 189042
rect 382280 89004 382332 89010
rect 382280 88946 382332 88952
rect 382188 4820 382240 4826
rect 382188 4762 382240 4768
rect 382292 1578 382320 88946
rect 383580 57254 383608 192086
rect 383856 189786 383884 192100
rect 384698 192086 384988 192114
rect 384304 189848 384356 189854
rect 384304 189790 384356 189796
rect 383844 189780 383896 189786
rect 383844 189722 383896 189728
rect 383660 62824 383712 62830
rect 383660 62766 383712 62772
rect 383568 57248 383620 57254
rect 383568 57190 383620 57196
rect 382372 11756 382424 11762
rect 382372 11698 382424 11704
rect 382384 3398 382412 11698
rect 383672 3482 383700 62766
rect 384316 17270 384344 189790
rect 384960 155242 384988 192086
rect 385512 189106 385540 192100
rect 385500 189100 385552 189106
rect 385500 189042 385552 189048
rect 386236 189100 386288 189106
rect 386236 189042 386288 189048
rect 384948 155236 385000 155242
rect 384948 155178 385000 155184
rect 386248 137290 386276 189042
rect 386236 137284 386288 137290
rect 386236 137226 386288 137232
rect 385040 91792 385092 91798
rect 385040 91734 385092 91740
rect 384304 17264 384356 17270
rect 384304 17206 384356 17212
rect 385052 3482 385080 91734
rect 386340 6186 386368 192100
rect 387182 192086 387748 192114
rect 387064 189916 387116 189922
rect 387064 189858 387116 189864
rect 387076 156670 387104 189858
rect 387064 156664 387116 156670
rect 387064 156606 387116 156612
rect 387720 32434 387748 192086
rect 387996 189106 388024 192100
rect 387984 189100 388036 189106
rect 387984 189042 388036 189048
rect 388824 188358 388852 192100
rect 389652 189446 389680 192100
rect 390388 192086 390494 192114
rect 391322 192086 391888 192114
rect 389640 189440 389692 189446
rect 389640 189382 389692 189388
rect 388996 189100 389048 189106
rect 388996 189042 389048 189048
rect 388812 188352 388864 188358
rect 388812 188294 388864 188300
rect 389008 55894 389036 189042
rect 390388 135930 390416 192086
rect 390468 189440 390520 189446
rect 390468 189382 390520 189388
rect 390376 135924 390428 135930
rect 390376 135866 390428 135872
rect 389180 93152 389232 93158
rect 389180 93094 389232 93100
rect 388996 55888 389048 55894
rect 388996 55830 389048 55836
rect 387800 42084 387852 42090
rect 387800 42026 387852 42032
rect 386420 32428 386472 32434
rect 386420 32370 386472 32376
rect 387708 32428 387760 32434
rect 387708 32370 387760 32376
rect 386328 6180 386380 6186
rect 386328 6122 386380 6128
rect 386432 3482 386460 32370
rect 387812 3482 387840 42026
rect 389192 3482 389220 93094
rect 390480 18630 390508 189382
rect 390560 178696 390612 178702
rect 390560 178638 390612 178644
rect 390468 18624 390520 18630
rect 390468 18566 390520 18572
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 386432 3454 387104 3482
rect 387812 3454 388300 3482
rect 389192 3454 389496 3482
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 1550 382412 1578
rect 379520 604 379572 610
rect 379520 546 379572 552
rect 379980 604 380032 610
rect 380912 598 381216 626
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 598
rect 382384 480 382412 1550
rect 383580 480 383608 3334
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 3454
rect 388272 480 388300 3454
rect 389468 480 389496 3454
rect 390572 3398 390600 178638
rect 390652 35216 390704 35222
rect 390652 35158 390704 35164
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 35158
rect 391860 11762 391888 192086
rect 392136 190262 392164 192100
rect 392978 192086 393268 192114
rect 392124 190256 392176 190262
rect 392124 190198 392176 190204
rect 393136 190256 393188 190262
rect 393136 190198 393188 190204
rect 393148 153882 393176 190198
rect 393136 153876 393188 153882
rect 393136 153818 393188 153824
rect 391940 94512 391992 94518
rect 391940 94454 391992 94460
rect 391848 11756 391900 11762
rect 391848 11698 391900 11704
rect 391952 3482 391980 94454
rect 393240 58682 393268 192086
rect 393792 186998 393820 192100
rect 393780 186992 393832 186998
rect 393780 186934 393832 186940
rect 393228 58676 393280 58682
rect 393228 58618 393280 58624
rect 394620 35222 394648 192100
rect 395462 192086 396028 192114
rect 396000 82142 396028 192086
rect 396276 185638 396304 192100
rect 397118 192086 397408 192114
rect 397946 192086 398696 192114
rect 396264 185632 396316 185638
rect 396264 185574 396316 185580
rect 397380 152522 397408 192086
rect 397368 152516 397420 152522
rect 397368 152458 397420 152464
rect 398668 133210 398696 192086
rect 398656 133204 398708 133210
rect 398656 133146 398708 133152
rect 396080 95940 396132 95946
rect 396080 95882 396132 95888
rect 395988 82136 396040 82142
rect 395988 82078 396040 82084
rect 394700 64184 394752 64190
rect 394700 64126 394752 64132
rect 394608 35216 394660 35222
rect 394608 35158 394660 35164
rect 393320 10328 393372 10334
rect 393320 10270 393372 10276
rect 393332 3482 393360 10270
rect 394712 3482 394740 64126
rect 396092 3482 396120 95882
rect 397460 15904 397512 15910
rect 397460 15846 397512 15852
rect 397472 3482 397500 15846
rect 398760 7614 398788 192100
rect 399602 192086 400168 192114
rect 398840 65544 398892 65550
rect 398840 65486 398892 65492
rect 398748 7608 398800 7614
rect 398748 7550 398800 7556
rect 398852 3482 398880 65486
rect 400140 15910 400168 192086
rect 400416 189106 400444 192100
rect 400404 189100 400456 189106
rect 400404 189042 400456 189048
rect 401244 184210 401272 192100
rect 402072 189106 402100 192100
rect 402808 192086 402914 192114
rect 403742 192086 404308 192114
rect 401508 189100 401560 189106
rect 401508 189042 401560 189048
rect 402060 189100 402112 189106
rect 402060 189042 402112 189048
rect 401232 184204 401284 184210
rect 401232 184146 401284 184152
rect 401520 131782 401548 189042
rect 401508 131776 401560 131782
rect 401508 131718 401560 131724
rect 402808 130422 402836 192086
rect 402888 189100 402940 189106
rect 402888 189042 402940 189048
rect 402796 130416 402848 130422
rect 402796 130358 402848 130364
rect 400220 97300 400272 97306
rect 400220 97242 400272 97248
rect 400128 15904 400180 15910
rect 400128 15846 400180 15852
rect 391952 3454 393084 3482
rect 393332 3454 394280 3482
rect 394712 3454 395476 3482
rect 396092 3454 396672 3482
rect 397472 3454 397868 3482
rect 398852 3454 399064 3482
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 393056 480 393084 3454
rect 394252 480 394280 3454
rect 395448 480 395476 3454
rect 396644 480 396672 3454
rect 397840 480 397868 3454
rect 399036 480 399064 3454
rect 400232 480 400260 97242
rect 401600 44872 401652 44878
rect 401600 44814 401652 44820
rect 401324 8968 401376 8974
rect 401324 8910 401376 8916
rect 401336 480 401364 8910
rect 401612 3482 401640 44814
rect 402900 42090 402928 189042
rect 402980 98660 403032 98666
rect 402980 98602 403032 98608
rect 402888 42084 402940 42090
rect 402888 42026 402940 42032
rect 402992 3482 403020 98602
rect 404280 13122 404308 192086
rect 404556 189106 404584 192100
rect 405306 192086 405688 192114
rect 404544 189100 404596 189106
rect 404544 189042 404596 189048
rect 405556 189100 405608 189106
rect 405556 189042 405608 189048
rect 405568 151094 405596 189042
rect 405556 151088 405608 151094
rect 405556 151030 405608 151036
rect 405660 62830 405688 192086
rect 406120 182850 406148 192100
rect 406962 192086 407068 192114
rect 407790 192086 408448 192114
rect 406108 182844 406160 182850
rect 406108 182786 406160 182792
rect 405740 90364 405792 90370
rect 405740 90306 405792 90312
rect 405648 62824 405700 62830
rect 405648 62766 405700 62772
rect 404360 19984 404412 19990
rect 404360 19926 404412 19932
rect 404268 13116 404320 13122
rect 404268 13058 404320 13064
rect 404372 3482 404400 19926
rect 405752 3482 405780 90306
rect 407040 47598 407068 192086
rect 407120 100020 407172 100026
rect 407120 99962 407172 99968
rect 407028 47592 407080 47598
rect 407028 47534 407080 47540
rect 407132 3482 407160 99962
rect 408420 86290 408448 192086
rect 408604 190194 408632 192100
rect 409446 192086 409828 192114
rect 408592 190188 408644 190194
rect 408592 190130 408644 190136
rect 409696 190188 409748 190194
rect 409696 190130 409748 190136
rect 409708 180130 409736 190130
rect 409696 180124 409748 180130
rect 409696 180066 409748 180072
rect 408500 104168 408552 104174
rect 408500 104110 408552 104116
rect 408408 86284 408460 86290
rect 408408 86226 408460 86232
rect 401612 3454 402560 3482
rect 402992 3454 403756 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 407132 3454 407344 3482
rect 402532 480 402560 3454
rect 403728 480 403756 3454
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407316 480 407344 3454
rect 408512 480 408540 104110
rect 409800 49026 409828 192086
rect 410260 189106 410288 192100
rect 411088 189854 411116 192100
rect 411930 192086 412588 192114
rect 411076 189848 411128 189854
rect 411076 189790 411128 189796
rect 410248 189100 410300 189106
rect 410248 189042 410300 189048
rect 411168 189100 411220 189106
rect 411168 189042 411220 189048
rect 409880 108316 409932 108322
rect 409880 108258 409932 108264
rect 409788 49020 409840 49026
rect 409788 48962 409840 48968
rect 408592 47660 408644 47666
rect 408592 47602 408644 47608
rect 408604 3482 408632 47602
rect 409892 3482 409920 108258
rect 411180 60042 411208 189042
rect 411168 60036 411220 60042
rect 411168 59978 411220 59984
rect 412560 21418 412588 192086
rect 412744 189378 412772 192100
rect 413586 192086 413876 192114
rect 412732 189372 412784 189378
rect 412732 189314 412784 189320
rect 413848 178702 413876 192086
rect 413928 189372 413980 189378
rect 413928 189314 413980 189320
rect 413836 178696 413888 178702
rect 413836 178638 413888 178644
rect 412640 66904 412692 66910
rect 412640 66846 412692 66852
rect 411260 21412 411312 21418
rect 411260 21354 411312 21360
rect 412548 21412 412600 21418
rect 412548 21354 412600 21360
rect 411272 3482 411300 21354
rect 412652 3482 412680 66846
rect 413940 61402 413968 189314
rect 414400 189106 414428 192100
rect 415242 192086 415348 192114
rect 416070 192086 416728 192114
rect 414388 189100 414440 189106
rect 414388 189042 414440 189048
rect 415320 129062 415348 192086
rect 416044 189100 416096 189106
rect 416044 189042 416096 189048
rect 415400 177336 415452 177342
rect 415400 177278 415452 177284
rect 415308 129056 415360 129062
rect 415308 128998 415360 129004
rect 414020 109744 414072 109750
rect 414020 109686 414072 109692
rect 413928 61396 413980 61402
rect 413928 61338 413980 61344
rect 414032 3482 414060 109686
rect 415412 3482 415440 177278
rect 416056 149734 416084 189042
rect 416044 149728 416096 149734
rect 416044 149670 416096 149676
rect 416700 19990 416728 192086
rect 416884 190262 416912 192100
rect 417726 192086 418108 192114
rect 416872 190256 416924 190262
rect 416872 190198 416924 190204
rect 417976 190256 418028 190262
rect 417976 190198 418028 190204
rect 417988 148374 418016 190198
rect 417976 148368 418028 148374
rect 417976 148310 418028 148316
rect 416780 101448 416832 101454
rect 416780 101390 416832 101396
rect 416688 19984 416740 19990
rect 416688 19926 416740 19932
rect 408604 3454 409736 3482
rect 409892 3454 410932 3482
rect 411272 3454 412128 3482
rect 412652 3454 413324 3482
rect 414032 3454 414520 3482
rect 415412 3454 415716 3482
rect 409708 480 409736 3454
rect 410904 480 410932 3454
rect 412100 480 412128 3454
rect 413296 480 413324 3454
rect 414492 480 414520 3454
rect 415688 480 415716 3454
rect 416792 3398 416820 101390
rect 418080 68338 418108 192086
rect 418540 189106 418568 192100
rect 419382 192086 419488 192114
rect 420210 192086 420868 192114
rect 418528 189100 418580 189106
rect 418528 189042 418580 189048
rect 416872 68332 416924 68338
rect 416872 68274 416924 68280
rect 418068 68332 418120 68338
rect 418068 68274 418120 68280
rect 416780 3392 416832 3398
rect 416780 3334 416832 3340
rect 416884 480 416912 68274
rect 419460 22778 419488 192086
rect 420184 189100 420236 189106
rect 420184 189042 420236 189048
rect 420196 177342 420224 189042
rect 420184 177336 420236 177342
rect 420184 177278 420236 177284
rect 420840 83502 420868 192086
rect 421024 189106 421052 192100
rect 421866 192086 422248 192114
rect 421012 189100 421064 189106
rect 421012 189042 421064 189048
rect 422116 189100 422168 189106
rect 422116 189042 422168 189048
rect 422128 175982 422156 189042
rect 422116 175976 422168 175982
rect 422116 175918 422168 175924
rect 420920 102808 420972 102814
rect 420920 102750 420972 102756
rect 420828 83496 420880 83502
rect 420828 83438 420880 83444
rect 419540 69692 419592 69698
rect 419540 69634 419592 69640
rect 418160 22772 418212 22778
rect 418160 22714 418212 22720
rect 419448 22772 419500 22778
rect 419448 22714 419500 22720
rect 418172 3482 418200 22714
rect 419552 3482 419580 69634
rect 420932 3482 420960 102750
rect 422220 24138 422248 192086
rect 422680 189106 422708 192100
rect 423522 192086 423628 192114
rect 424350 192086 425008 192114
rect 422668 189100 422720 189106
rect 422668 189042 422720 189048
rect 423496 189100 423548 189106
rect 423496 189042 423548 189048
rect 423508 127634 423536 189042
rect 423496 127628 423548 127634
rect 423496 127570 423548 127576
rect 422300 24200 422352 24206
rect 422300 24142 422352 24148
rect 422208 24132 422260 24138
rect 422208 24074 422260 24080
rect 422312 3482 422340 24142
rect 423600 10334 423628 192086
rect 423680 71052 423732 71058
rect 423680 70994 423732 71000
rect 423588 10328 423640 10334
rect 423588 10270 423640 10276
rect 423692 3482 423720 70994
rect 424980 44878 425008 192086
rect 425164 189310 425192 192100
rect 426006 192086 426296 192114
rect 425152 189304 425204 189310
rect 425152 189246 425204 189252
rect 426268 174554 426296 192086
rect 426348 189304 426400 189310
rect 426348 189246 426400 189252
rect 426256 174548 426308 174554
rect 426256 174490 426308 174496
rect 425060 106956 425112 106962
rect 425060 106898 425112 106904
rect 424968 44872 425020 44878
rect 424968 44814 425020 44820
rect 425072 3482 425100 106898
rect 426360 65550 426388 189246
rect 426820 189106 426848 192100
rect 427662 192086 427768 192114
rect 426808 189100 426860 189106
rect 426808 189042 426860 189048
rect 427636 189100 427688 189106
rect 427636 189042 427688 189048
rect 427648 146946 427676 189042
rect 427636 146940 427688 146946
rect 427636 146882 427688 146888
rect 427740 84862 427768 192086
rect 428384 189106 428412 192100
rect 429212 189990 429240 192100
rect 430054 192086 430528 192114
rect 429200 189984 429252 189990
rect 429200 189926 429252 189932
rect 430396 189984 430448 189990
rect 430396 189926 430448 189932
rect 428372 189100 428424 189106
rect 428372 189042 428424 189048
rect 429108 189100 429160 189106
rect 429108 189042 429160 189048
rect 427820 112464 427872 112470
rect 427820 112406 427872 112412
rect 427728 84856 427780 84862
rect 427728 84798 427780 84804
rect 426440 72480 426492 72486
rect 426440 72422 426492 72428
rect 426348 65544 426400 65550
rect 426348 65486 426400 65492
rect 425152 37936 425204 37942
rect 425152 37878 425204 37884
rect 425164 4214 425192 37878
rect 425152 4208 425204 4214
rect 425152 4150 425204 4156
rect 426348 4208 426400 4214
rect 426348 4150 426400 4156
rect 418172 3454 419212 3482
rect 419552 3454 420408 3482
rect 420932 3454 421604 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 425072 3454 425192 3482
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 417988 480 418016 3334
rect 419184 480 419212 3454
rect 420380 480 420408 3454
rect 421576 480 421604 3454
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425164 480 425192 3454
rect 426360 480 426388 4150
rect 426452 3482 426480 72422
rect 427832 3482 427860 112406
rect 429120 25566 429148 189042
rect 430408 145586 430436 189926
rect 430396 145580 430448 145586
rect 430396 145522 430448 145528
rect 430500 66910 430528 192086
rect 430868 189106 430896 192100
rect 431710 192086 431908 192114
rect 432538 192086 433288 192114
rect 430856 189100 430908 189106
rect 430856 189042 430908 189048
rect 431776 189100 431828 189106
rect 431776 189042 431828 189048
rect 431788 173194 431816 189042
rect 431776 173188 431828 173194
rect 431776 173130 431828 173136
rect 430580 73840 430632 73846
rect 430580 73782 430632 73788
rect 430488 66904 430540 66910
rect 430488 66846 430540 66852
rect 429108 25560 429160 25566
rect 429108 25502 429160 25508
rect 429200 14476 429252 14482
rect 429200 14418 429252 14424
rect 429212 3482 429240 14418
rect 430592 3482 430620 73782
rect 431880 37942 431908 192086
rect 433260 126274 433288 192086
rect 433352 190126 433380 192100
rect 434194 192086 434668 192114
rect 433340 190120 433392 190126
rect 433340 190062 433392 190068
rect 434536 190120 434588 190126
rect 434536 190062 434588 190068
rect 434548 171834 434576 190062
rect 434536 171828 434588 171834
rect 434536 171770 434588 171776
rect 433248 126268 433300 126274
rect 433248 126210 433300 126216
rect 433340 75200 433392 75206
rect 433340 75142 433392 75148
rect 431960 50380 432012 50386
rect 431960 50322 432012 50328
rect 431868 37936 431920 37942
rect 431868 37878 431920 37884
rect 431972 3482 432000 50322
rect 426452 3454 427584 3482
rect 427832 3454 428780 3482
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 431972 3454 432368 3482
rect 427556 480 427584 3454
rect 428752 480 428780 3454
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3454
rect 433352 3398 433380 75142
rect 434640 50386 434668 192086
rect 435008 190262 435036 192100
rect 435850 192086 436048 192114
rect 434996 190256 435048 190262
rect 434996 190198 435048 190204
rect 435916 190256 435968 190262
rect 435916 190198 435968 190204
rect 435928 124914 435956 190198
rect 435916 124908 435968 124914
rect 435916 124850 435968 124856
rect 434720 105596 434772 105602
rect 434720 105538 434772 105544
rect 434628 50380 434680 50386
rect 434628 50322 434680 50328
rect 433432 31068 433484 31074
rect 433432 31010 433484 31016
rect 433444 3482 433472 31010
rect 434732 3482 434760 105538
rect 436020 14482 436048 192086
rect 436664 189106 436692 192100
rect 437492 189310 437520 192100
rect 438334 192086 438716 192114
rect 437480 189304 437532 189310
rect 437480 189246 437532 189252
rect 436652 189100 436704 189106
rect 436652 189042 436704 189048
rect 437388 189100 437440 189106
rect 437388 189042 437440 189048
rect 437400 144226 437428 189042
rect 438688 169046 438716 192086
rect 439148 189310 439176 192100
rect 439990 192086 440188 192114
rect 440818 192086 441568 192114
rect 438768 189304 438820 189310
rect 438768 189246 438820 189252
rect 439136 189304 439188 189310
rect 439136 189246 439188 189252
rect 440056 189304 440108 189310
rect 440056 189246 440108 189252
rect 438676 169040 438728 169046
rect 438676 168982 438728 168988
rect 437388 144220 437440 144226
rect 437388 144162 437440 144168
rect 438780 69698 438808 189246
rect 440068 142866 440096 189246
rect 440056 142860 440108 142866
rect 440056 142802 440108 142808
rect 438860 113824 438912 113830
rect 438860 113766 438912 113772
rect 438768 69692 438820 69698
rect 438768 69634 438820 69640
rect 437480 51740 437532 51746
rect 437480 51682 437532 51688
rect 436100 17264 436152 17270
rect 436100 17206 436152 17212
rect 436008 14476 436060 14482
rect 436008 14418 436060 14424
rect 436112 3482 436140 17206
rect 437492 3482 437520 51682
rect 438872 3482 438900 113766
rect 440160 71058 440188 192086
rect 440148 71052 440200 71058
rect 440148 70994 440200 71000
rect 440240 33788 440292 33794
rect 440240 33730 440292 33736
rect 440252 3482 440280 33730
rect 441540 31074 441568 192086
rect 441632 190194 441660 192100
rect 442474 192086 442948 192114
rect 441620 190188 441672 190194
rect 441620 190130 441672 190136
rect 442816 190188 442868 190194
rect 442816 190130 442868 190136
rect 442828 141438 442856 190130
rect 442816 141432 442868 141438
rect 442816 141374 442868 141380
rect 441620 76560 441672 76566
rect 441620 76502 441672 76508
rect 441528 31068 441580 31074
rect 441528 31010 441580 31016
rect 433444 3454 433564 3482
rect 434732 3454 435864 3482
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 440252 3454 440648 3482
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433536 480 433564 3454
rect 434628 3392 434680 3398
rect 434628 3334 434680 3340
rect 434640 480 434668 3334
rect 435836 480 435864 3454
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 3454
rect 441632 3346 441660 76502
rect 442920 72486 442948 192086
rect 443288 189106 443316 192100
rect 444130 192086 444328 192114
rect 443276 189100 443328 189106
rect 443276 189042 443328 189048
rect 444196 189100 444248 189106
rect 444196 189042 444248 189048
rect 444208 167686 444236 189042
rect 444196 167680 444248 167686
rect 444196 167622 444248 167628
rect 443000 166320 443052 166326
rect 443000 166262 443052 166268
rect 442908 72480 442960 72486
rect 442908 72422 442960 72428
rect 441632 3318 441844 3346
rect 441816 480 441844 3318
rect 443012 480 443040 166262
rect 444300 51746 444328 192086
rect 444944 189106 444972 192100
rect 445772 189990 445800 192100
rect 446614 192086 447088 192114
rect 445760 189984 445812 189990
rect 445760 189926 445812 189932
rect 446956 189984 447008 189990
rect 446956 189926 447008 189932
rect 444932 189100 444984 189106
rect 444932 189042 444984 189048
rect 445668 189100 445720 189106
rect 445668 189042 445720 189048
rect 445680 79354 445708 189042
rect 446968 166326 446996 189926
rect 446956 166320 447008 166326
rect 446956 166262 447008 166268
rect 444380 79348 444432 79354
rect 444380 79290 444432 79296
rect 445668 79348 445720 79354
rect 445668 79290 445720 79296
rect 444288 51740 444340 51746
rect 444288 51682 444340 51688
rect 443092 40724 443144 40730
rect 443092 40666 443144 40672
rect 443104 3346 443132 40666
rect 444392 3346 444420 79290
rect 447060 33794 447088 192086
rect 447428 189106 447456 192100
rect 448270 192086 448376 192114
rect 449098 192086 449848 192114
rect 447416 189100 447468 189106
rect 447416 189042 447468 189048
rect 448348 164898 448376 192086
rect 448428 189100 448480 189106
rect 448428 189042 448480 189048
rect 448336 164892 448388 164898
rect 448336 164834 448388 164840
rect 447140 36576 447192 36582
rect 447140 36518 447192 36524
rect 447048 33788 447100 33794
rect 447048 33730 447100 33736
rect 446588 3528 446640 3534
rect 446588 3470 446640 3476
rect 443104 3318 444236 3346
rect 444392 3318 445432 3346
rect 444208 480 444236 3318
rect 445404 480 445432 3318
rect 446600 480 446628 3470
rect 447152 3346 447180 36518
rect 448440 3534 448468 189042
rect 448520 53100 448572 53106
rect 448520 53042 448572 53048
rect 448428 3528 448480 3534
rect 448428 3470 448480 3476
rect 448532 3346 448560 53042
rect 449820 36582 449848 192086
rect 449912 189106 449940 192100
rect 451924 189848 451976 189854
rect 451924 189790 451976 189796
rect 449900 189100 449952 189106
rect 449900 189042 449952 189048
rect 451188 189100 451240 189106
rect 451188 189042 451240 189048
rect 449808 36576 449860 36582
rect 449808 36518 449860 36524
rect 451200 3466 451228 189042
rect 451280 77988 451332 77994
rect 451280 77930 451332 77936
rect 451292 4214 451320 77930
rect 451372 43444 451424 43450
rect 451372 43386 451424 43392
rect 451280 4208 451332 4214
rect 451280 4150 451332 4156
rect 451384 3482 451412 43386
rect 451936 8974 451964 189790
rect 453316 30326 453344 202671
rect 453408 77246 453436 224023
rect 453500 124166 453528 245375
rect 453592 171086 453620 266727
rect 453684 182170 453712 273799
rect 453946 259720 454002 259729
rect 453946 259655 454002 259664
rect 453960 259486 453988 259655
rect 453948 259480 454000 259486
rect 453948 259422 454000 259428
rect 456076 252550 456104 302330
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 461584 280220 461636 280226
rect 461584 280162 461636 280168
rect 456064 252544 456116 252550
rect 456064 252486 456116 252492
rect 457444 251252 457496 251258
rect 457444 251194 457496 251200
rect 453946 238368 454002 238377
rect 453946 238303 454002 238312
rect 453960 237454 453988 238303
rect 453948 237448 454000 237454
rect 453948 237390 454000 237396
rect 453762 217016 453818 217025
rect 453762 216951 453818 216960
rect 453776 216850 453804 216951
rect 453764 216844 453816 216850
rect 453764 216786 453816 216792
rect 456064 216844 456116 216850
rect 456064 216786 456116 216792
rect 453948 209840 454000 209846
rect 453946 209808 453948 209817
rect 454000 209808 454002 209817
rect 453946 209743 454002 209752
rect 453946 195664 454002 195673
rect 453946 195599 454002 195608
rect 453960 194614 453988 195599
rect 453948 194608 454000 194614
rect 453948 194550 454000 194556
rect 453672 182164 453724 182170
rect 453672 182106 453724 182112
rect 453580 171080 453632 171086
rect 453580 171022 453632 171028
rect 453488 124160 453540 124166
rect 453488 124102 453540 124108
rect 455420 80708 455472 80714
rect 455420 80650 455472 80656
rect 453396 77240 453448 77246
rect 453396 77182 453448 77188
rect 454040 39364 454092 39370
rect 454040 39306 454092 39312
rect 453304 30320 453356 30326
rect 453304 30262 453356 30268
rect 451924 8968 451976 8974
rect 451924 8910 451976 8916
rect 452476 4208 452528 4214
rect 452476 4150 452528 4156
rect 450176 3460 450228 3466
rect 450176 3402 450228 3408
rect 451188 3460 451240 3466
rect 451188 3402 451240 3408
rect 451292 3454 451412 3482
rect 447152 3318 447824 3346
rect 448532 3318 449020 3346
rect 447796 480 447824 3318
rect 448992 480 449020 3318
rect 450188 480 450216 3402
rect 451292 480 451320 3454
rect 452488 480 452516 4150
rect 453672 4140 453724 4146
rect 453672 4082 453724 4088
rect 453684 480 453712 4082
rect 454052 3482 454080 39306
rect 455432 3482 455460 80650
rect 456076 64870 456104 216786
rect 457456 135250 457484 251194
rect 461596 205630 461624 280162
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 471244 259480 471296 259486
rect 471244 259422 471296 259428
rect 469864 237448 469916 237454
rect 469864 237390 469916 237396
rect 461584 205624 461636 205630
rect 461584 205566 461636 205572
rect 462320 181484 462372 181490
rect 462320 181426 462372 181432
rect 458180 163532 458232 163538
rect 458180 163474 458232 163480
rect 457444 135244 457496 135250
rect 457444 135186 457496 135192
rect 456064 64864 456116 64870
rect 456064 64806 456116 64812
rect 457260 4072 457312 4078
rect 457260 4014 457312 4020
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 4014
rect 458192 3482 458220 163474
rect 460940 162172 460992 162178
rect 460940 162114 460992 162120
rect 459652 158024 459704 158030
rect 459652 157966 459704 157972
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 157966
rect 460848 4004 460900 4010
rect 460848 3946 460900 3952
rect 460860 480 460888 3946
rect 460952 3482 460980 162114
rect 462332 3482 462360 181426
rect 466460 140072 466512 140078
rect 466460 140014 466512 140020
rect 465080 28280 465132 28286
rect 465080 28222 465132 28228
rect 464436 3936 464488 3942
rect 464436 3878 464488 3884
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3878
rect 465092 3482 465120 28222
rect 466472 3482 466500 140014
rect 469876 111790 469904 237390
rect 471256 158710 471284 259422
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 474004 230512 474056 230518
rect 474004 230454 474056 230460
rect 471244 158704 471296 158710
rect 471244 158646 471296 158652
rect 469864 111784 469916 111790
rect 469864 111726 469916 111732
rect 469220 111104 469272 111110
rect 469220 111046 469272 111052
rect 467932 26920 467984 26926
rect 467932 26862 467984 26868
rect 467840 3800 467892 3806
rect 467840 3742 467892 3748
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 3210 467880 3742
rect 467944 3398 467972 26862
rect 469232 3482 469260 111046
rect 474016 88330 474044 230454
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 478144 209840 478196 209846
rect 478144 209782 478196 209788
rect 476120 160744 476172 160750
rect 476120 160686 476172 160692
rect 474004 88324 474056 88330
rect 474004 88266 474056 88272
rect 473360 87644 473412 87650
rect 473360 87586 473412 87592
rect 471980 46232 472032 46238
rect 471980 46174 472032 46180
rect 471520 3868 471572 3874
rect 471520 3810 471572 3816
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 3182 467972 3210
rect 467944 480 467972 3182
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3810
rect 471992 3482 472020 46174
rect 473372 3482 473400 87586
rect 475108 3664 475160 3670
rect 475108 3606 475160 3612
rect 471992 3454 472756 3482
rect 473372 3454 473952 3482
rect 472728 480 472756 3454
rect 473924 480 473952 3454
rect 475120 480 475148 3606
rect 476132 3482 476160 160686
rect 477592 54528 477644 54534
rect 477592 54470 477644 54476
rect 477604 3482 477632 54470
rect 478156 41410 478184 209782
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 483664 194608 483716 194614
rect 483664 194550 483716 194556
rect 478880 159384 478932 159390
rect 478880 159326 478932 159332
rect 478144 41404 478196 41410
rect 478144 41346 478196 41352
rect 478696 3732 478748 3738
rect 478696 3674 478748 3680
rect 476132 3454 476344 3482
rect 476316 480 476344 3454
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 3674
rect 478892 3482 478920 159326
rect 480260 138712 480312 138718
rect 480260 138654 480312 138660
rect 480272 3482 480300 138654
rect 483676 17950 483704 194550
rect 485780 189780 485832 189786
rect 485780 189722 485832 189728
rect 484400 156664 484452 156670
rect 484400 156606 484452 156612
rect 483664 17944 483716 17950
rect 483664 17886 483716 17892
rect 483480 4820 483532 4826
rect 483480 4762 483532 4768
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 478892 3454 479932 3482
rect 480272 3454 481128 3482
rect 479904 480 479932 3454
rect 481100 480 481128 3454
rect 482296 480 482324 3538
rect 483492 480 483520 4762
rect 484412 3482 484440 156606
rect 485792 3602 485820 189722
rect 494060 188352 494112 188358
rect 494060 188294 494112 188300
rect 487160 155236 487212 155242
rect 487160 155178 487212 155184
rect 485872 57248 485924 57254
rect 485872 57190 485924 57196
rect 485780 3596 485832 3602
rect 485780 3538 485832 3544
rect 485884 3482 485912 57190
rect 486976 3596 487028 3602
rect 486976 3538 487028 3544
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 3454 485912 3482
rect 485792 480 485820 3454
rect 486988 480 487016 3538
rect 487172 3482 487200 155178
rect 488540 137284 488592 137290
rect 488540 137226 488592 137232
rect 488552 3482 488580 137226
rect 492680 55888 492732 55894
rect 492680 55830 492732 55836
rect 491300 32428 491352 32434
rect 491300 32370 491352 32376
rect 490564 6180 490616 6186
rect 490564 6122 490616 6128
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 490576 480 490604 6122
rect 491312 1306 491340 32370
rect 492692 3482 492720 55830
rect 494072 3482 494100 188294
rect 500960 186992 501012 186998
rect 500960 186934 501012 186940
rect 498200 153876 498252 153882
rect 498200 153818 498252 153824
rect 495440 135924 495492 135930
rect 495440 135866 495492 135872
rect 494152 18624 494204 18630
rect 494152 18566 494204 18572
rect 494164 3602 494192 18566
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 492692 3454 492996 3482
rect 494072 3454 494192 3482
rect 491312 1278 491800 1306
rect 491772 480 491800 1278
rect 492968 480 492996 3454
rect 494164 480 494192 3454
rect 495360 480 495388 3538
rect 495452 3482 495480 135866
rect 496820 11756 496872 11762
rect 496820 11698 496872 11704
rect 496832 3482 496860 11698
rect 498212 3482 498240 153818
rect 499580 58676 499632 58682
rect 499580 58618 499632 58624
rect 495452 3454 496584 3482
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 496556 480 496584 3454
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 499592 610 499620 58618
rect 500972 610 501000 186934
rect 503720 185632 503772 185638
rect 503720 185574 503772 185580
rect 502340 82136 502392 82142
rect 502340 82078 502392 82084
rect 502352 2786 502380 82078
rect 502432 35216 502484 35222
rect 502432 35158 502484 35164
rect 502340 2780 502392 2786
rect 502340 2722 502392 2728
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500960 604 501012 610
rect 500960 546 501012 552
rect 501236 604 501288 610
rect 501236 546 501288 552
rect 500144 480 500172 546
rect 501248 480 501276 546
rect 502444 480 502472 35158
rect 503628 2780 503680 2786
rect 503628 2722 503680 2728
rect 503640 480 503668 2722
rect 503732 610 503760 185574
rect 512000 184204 512052 184210
rect 512000 184146 512052 184152
rect 505100 152516 505152 152522
rect 505100 152458 505152 152464
rect 505112 610 505140 152458
rect 506480 133204 506532 133210
rect 506480 133146 506532 133152
rect 506492 610 506520 133146
rect 510620 131776 510672 131782
rect 510620 131718 510672 131724
rect 509240 15904 509292 15910
rect 509240 15846 509292 15852
rect 508412 7608 508464 7614
rect 508412 7550 508464 7556
rect 503720 604 503772 610
rect 503720 546 503772 552
rect 504824 604 504876 610
rect 504824 546 504876 552
rect 505100 604 505152 610
rect 505100 546 505152 552
rect 506020 604 506072 610
rect 506020 546 506072 552
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 504836 480 504864 546
rect 506032 480 506060 546
rect 507228 480 507256 546
rect 508424 480 508452 7550
rect 509252 3482 509280 15846
rect 510632 3482 510660 131718
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 480 512040 184146
rect 518900 182844 518952 182850
rect 518900 182786 518952 182792
rect 516140 151088 516192 151094
rect 516140 151030 516192 151036
rect 513380 130416 513432 130422
rect 513380 130358 513432 130364
rect 512092 42084 512144 42090
rect 512092 42026 512144 42032
rect 512104 3482 512132 42026
rect 513392 3482 513420 130358
rect 514760 13116 514812 13122
rect 514760 13058 514812 13064
rect 514772 3482 514800 13058
rect 516152 3482 516180 151030
rect 517520 62824 517572 62830
rect 517520 62766 517572 62772
rect 517532 3482 517560 62766
rect 518912 3482 518940 182786
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 521660 180124 521712 180130
rect 521660 180066 521712 180072
rect 520280 86284 520332 86290
rect 520280 86226 520332 86232
rect 520292 3602 520320 86226
rect 520372 47592 520424 47598
rect 520372 47534 520424 47540
rect 520280 3596 520332 3602
rect 520280 3538 520332 3544
rect 512104 3454 513236 3482
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513208 480 513236 3454
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520384 1578 520412 47534
rect 521476 3596 521528 3602
rect 521476 3538 521528 3544
rect 520292 1550 520412 1578
rect 520292 480 520320 1550
rect 521488 480 521516 3538
rect 521672 3482 521700 180066
rect 528560 178696 528612 178702
rect 528560 178638 528612 178644
rect 524420 60036 524472 60042
rect 524420 59978 524472 59984
rect 523040 49020 523092 49026
rect 523040 48962 523092 48968
rect 523052 3482 523080 48962
rect 524432 3482 524460 59978
rect 527180 21412 527232 21418
rect 527180 21354 527232 21360
rect 526260 8968 526312 8974
rect 526260 8910 526312 8916
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 8910
rect 527192 3482 527220 21354
rect 528572 3602 528600 178638
rect 536840 177336 536892 177342
rect 536840 177278 536892 177284
rect 529940 149728 529992 149734
rect 529940 149670 529992 149676
rect 528652 61396 528704 61402
rect 528652 61338 528704 61344
rect 528560 3596 528612 3602
rect 528560 3538 528612 3544
rect 527192 3454 527496 3482
rect 527468 480 527496 3454
rect 528664 480 528692 61338
rect 529848 3596 529900 3602
rect 529848 3538 529900 3544
rect 529860 480 529888 3538
rect 529952 3482 529980 149670
rect 534080 148368 534132 148374
rect 534080 148310 534132 148316
rect 531320 129056 531372 129062
rect 531320 128998 531372 129004
rect 531332 3482 531360 128998
rect 532700 19984 532752 19990
rect 532700 19926 532752 19932
rect 532712 3482 532740 19926
rect 534092 3482 534120 148310
rect 535460 68332 535512 68338
rect 535460 68274 535512 68280
rect 535472 3482 535500 68274
rect 536852 3482 536880 177278
rect 539600 175976 539652 175982
rect 539600 175918 539652 175924
rect 538220 83496 538272 83502
rect 538220 83438 538272 83444
rect 536932 22772 536984 22778
rect 536932 22714 536984 22720
rect 536944 3602 536972 22714
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 538128 3596 538180 3602
rect 538128 3538 538180 3544
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 3538
rect 538232 3482 538260 83438
rect 539612 3482 539640 175918
rect 546500 174548 546552 174554
rect 546500 174490 546552 174496
rect 542360 127628 542412 127634
rect 542360 127570 542412 127576
rect 540980 24132 541032 24138
rect 540980 24074 541032 24080
rect 540992 3482 541020 24074
rect 542372 3482 542400 127570
rect 545120 44872 545172 44878
rect 545120 44814 545172 44820
rect 543740 10328 543792 10334
rect 543740 10270 543792 10276
rect 543752 3482 543780 10270
rect 545132 3482 545160 44814
rect 546512 3602 546540 174490
rect 554780 173188 554832 173194
rect 554780 173130 554832 173136
rect 547880 146940 547932 146946
rect 547880 146882 547932 146888
rect 546592 65544 546644 65550
rect 546592 65486 546644 65492
rect 546500 3596 546552 3602
rect 546500 3538 546552 3544
rect 546604 3482 546632 65486
rect 547696 3596 547748 3602
rect 547696 3538 547748 3544
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 3454 546632 3482
rect 546512 480 546540 3454
rect 547708 480 547736 3538
rect 547892 3482 547920 146882
rect 552020 145580 552072 145586
rect 552020 145522 552072 145528
rect 549260 84856 549312 84862
rect 549260 84798 549312 84804
rect 549272 3482 549300 84798
rect 550640 25560 550692 25566
rect 550640 25502 550692 25508
rect 550652 3482 550680 25502
rect 552032 3482 552060 145522
rect 553400 66904 553452 66910
rect 553400 66846 553452 66852
rect 553412 3482 553440 66846
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 173130
rect 557540 171828 557592 171834
rect 557540 171770 557592 171776
rect 556160 126268 556212 126274
rect 556160 126210 556212 126216
rect 554872 37936 554924 37942
rect 554872 37878 554924 37884
rect 554884 3482 554912 37878
rect 556172 3482 556200 126210
rect 557552 3482 557580 171770
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 564440 169040 564492 169046
rect 564440 168982 564492 168988
rect 563060 144220 563112 144226
rect 563060 144162 563112 144168
rect 560300 124908 560352 124914
rect 560300 124850 560352 124856
rect 558920 50380 558972 50386
rect 558920 50322 558972 50328
rect 558932 3482 558960 50322
rect 560312 3482 560340 124850
rect 561680 14476 561732 14482
rect 561680 14418 561732 14424
rect 561692 3482 561720 14418
rect 563072 3482 563100 144162
rect 563152 69692 563204 69698
rect 563152 69634 563204 69640
rect 563164 3602 563192 69634
rect 563152 3596 563204 3602
rect 563152 3538 563204 3544
rect 564348 3596 564400 3602
rect 564348 3538 564400 3544
rect 554884 3454 556016 3482
rect 556172 3454 557212 3482
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 560312 3454 560800 3482
rect 561692 3454 561996 3482
rect 563072 3454 563192 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3454
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3454
rect 561968 480 561996 3454
rect 563164 480 563192 3454
rect 564360 480 564388 3538
rect 564452 3482 564480 168982
rect 571340 167680 571392 167686
rect 571340 167622 571392 167628
rect 565820 142860 565872 142866
rect 565820 142802 565872 142808
rect 565832 3482 565860 142802
rect 569960 141432 570012 141438
rect 569960 141374 570012 141380
rect 567200 71052 567252 71058
rect 567200 70994 567252 71000
rect 567212 3482 567240 70994
rect 568580 31068 568632 31074
rect 568580 31010 568632 31016
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 567212 3454 567884 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3454
rect 568592 1306 568620 31010
rect 569972 3482 570000 141374
rect 569972 3454 570276 3482
rect 568592 1278 569080 1306
rect 569052 480 569080 1278
rect 570248 480 570276 3454
rect 571352 3330 571380 167622
rect 575480 166320 575532 166326
rect 575480 166262 575532 166268
rect 574100 79348 574152 79354
rect 574100 79290 574152 79296
rect 571432 72480 571484 72486
rect 571432 72422 571484 72428
rect 571340 3324 571392 3330
rect 571340 3266 571392 3272
rect 571444 480 571472 72422
rect 572720 51740 572772 51746
rect 572720 51682 572772 51688
rect 572732 3482 572760 51682
rect 574112 3482 574140 79290
rect 575492 3482 575520 166262
rect 578884 164892 578936 164898
rect 578884 164834 578936 164840
rect 576860 33788 576912 33794
rect 576860 33730 576912 33736
rect 572732 3454 573864 3482
rect 574112 3454 575060 3482
rect 575492 3454 576256 3482
rect 572628 3324 572680 3330
rect 572628 3266 572680 3272
rect 572640 480 572668 3266
rect 573836 480 573864 3454
rect 575032 480 575060 3454
rect 576228 480 576256 3454
rect 576872 610 576900 33730
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 576860 604 576912 610
rect 576860 546 576912 552
rect 577412 604 577464 610
rect 577412 546 577464 552
rect 577424 480 577452 546
rect 578620 480 578648 3470
rect 578896 3330 578924 164834
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 578976 36576 579028 36582
rect 578976 36518 579028 36524
rect 578988 3534 579016 36518
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 578976 3528 579028 3534
rect 578976 3470 579028 3476
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 578884 3324 578936 3330
rect 578884 3266 578936 3272
rect 579804 3324 579856 3330
rect 579804 3266 579856 3272
rect 579816 480 579844 3266
rect 581012 480 581040 3470
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3330 682216 3386 682272
rect 3422 667936 3478 667992
rect 3054 653520 3110 653576
rect 3238 624824 3294 624880
rect 3330 595992 3386 596048
rect 3238 509904 3294 509960
rect 3514 610408 3570 610464
rect 3422 495488 3478 495544
rect 4066 567316 4122 567352
rect 4066 567296 4068 567316
rect 4068 567296 4120 567316
rect 4120 567296 4122 567316
rect 3606 553016 3662 553072
rect 3698 538600 3754 538656
rect 3514 452376 3570 452432
rect 3422 423680 3478 423736
rect 8206 540912 8262 540968
rect 8390 540912 8446 540968
rect 8114 531256 8170 531312
rect 8298 531256 8354 531312
rect 3790 481072 3846 481128
rect 3606 437960 3662 438016
rect 72974 608504 73030 608560
rect 73158 608504 73214 608560
rect 128358 508544 128414 508600
rect 128358 500928 128414 500984
rect 154210 540912 154266 540968
rect 154486 540912 154542 540968
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 284206 540912 284262 540968
rect 284390 540912 284446 540968
rect 284114 531256 284170 531312
rect 284298 531256 284354 531312
rect 347870 560224 347926 560280
rect 348054 560224 348110 560280
rect 364430 560224 364486 560280
rect 364614 560224 364670 560280
rect 347870 540912 347926 540968
rect 348054 540912 348110 540968
rect 364430 540912 364486 540968
rect 364614 540912 364670 540968
rect 453210 508816 453266 508872
rect 453394 501744 453450 501800
rect 453946 494536 454002 494592
rect 129002 493312 129058 493368
rect 453762 487464 453818 487520
rect 128358 485732 128360 485752
rect 128360 485732 128412 485752
rect 128412 485732 128414 485752
rect 128358 485696 128414 485732
rect 453762 480392 453818 480448
rect 128358 478080 128414 478136
rect 453946 473184 454002 473240
rect 128358 470500 128360 470520
rect 128360 470500 128412 470520
rect 128412 470500 128414 470520
rect 128358 470464 128414 470500
rect 452750 466112 452806 466168
rect 128358 462848 128414 462904
rect 453394 459040 453450 459096
rect 128358 455232 128414 455288
rect 453946 451832 454002 451888
rect 128358 447616 128414 447672
rect 453670 444760 453726 444816
rect 128358 440000 128414 440056
rect 128358 432248 128414 432304
rect 128358 424632 128414 424688
rect 128358 417016 128414 417072
rect 128358 409400 128414 409456
rect 128358 401784 128414 401840
rect 3422 394984 3478 395040
rect 128358 394168 128414 394224
rect 453762 437688 453818 437744
rect 453946 430516 453948 430536
rect 453948 430516 454000 430536
rect 454000 430516 454002 430536
rect 453946 430480 454002 430516
rect 453946 423408 454002 423464
rect 453946 416372 453948 416392
rect 453948 416372 454000 416392
rect 454000 416372 454002 416392
rect 453946 416336 454002 416372
rect 477590 560224 477646 560280
rect 477774 560224 477830 560280
rect 477590 540912 477646 540968
rect 477774 540912 477830 540968
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 494150 560224 494206 560280
rect 494334 560224 494390 560280
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 580170 697992 580226 698048
rect 580262 686296 580318 686352
rect 542358 683168 542414 683224
rect 542726 683168 542782 683224
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 579894 592456 579950 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 579894 545536 579950 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580354 639376 580410 639432
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 453394 409128 453450 409184
rect 580262 451696 580318 451752
rect 579894 439864 579950 439920
rect 578882 416472 578938 416528
rect 453946 402056 454002 402112
rect 453762 394848 453818 394904
rect 453302 387776 453358 387832
rect 129002 386552 129058 386608
rect 453946 380704 454002 380760
rect 3238 380568 3294 380624
rect 129002 378936 129058 378992
rect 453394 373496 453450 373552
rect 129278 371320 129334 371376
rect 3146 366152 3202 366208
rect 129002 363704 129058 363760
rect 128358 348336 128414 348392
rect 3330 308760 3386 308816
rect 3514 337456 3570 337512
rect 128358 333104 128414 333160
rect 3514 323040 3570 323096
rect 3422 294344 3478 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3146 222536 3202 222592
rect 3146 208156 3148 208176
rect 3148 208156 3200 208176
rect 3200 208156 3202 208176
rect 3146 208120 3202 208156
rect 2870 193840 2926 193896
rect 3238 179424 3294 179480
rect 3514 265648 3570 265704
rect 3514 251232 3570 251288
rect 3514 236952 3570 237008
rect 128358 325488 128414 325544
rect 129186 356088 129242 356144
rect 129094 340720 129150 340776
rect 129002 317872 129058 317928
rect 128358 310256 128414 310312
rect 3422 165008 3478 165064
rect 3146 150728 3202 150784
rect 3422 136312 3478 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3422 78920 3478 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 128358 302640 128414 302696
rect 128358 287408 128414 287464
rect 128266 279792 128322 279848
rect 128358 264424 128414 264480
rect 128358 256808 128414 256864
rect 128358 241576 128414 241632
rect 580354 404776 580410 404832
rect 580170 392944 580226 393000
rect 580262 369552 580318 369608
rect 453946 366424 454002 366480
rect 453946 359352 454002 359408
rect 580262 357856 580318 357912
rect 453762 352144 453818 352200
rect 580170 346024 580226 346080
rect 453946 345072 454002 345128
rect 453486 338000 453542 338056
rect 453394 330792 453450 330848
rect 453302 323720 453358 323776
rect 580170 322632 580226 322688
rect 453578 316648 453634 316704
rect 453486 309440 453542 309496
rect 453394 295160 453450 295216
rect 129370 295024 129426 295080
rect 129278 272040 129334 272096
rect 129186 249192 129242 249248
rect 128358 233960 128414 234016
rect 129094 226344 129150 226400
rect 128358 218728 128414 218784
rect 128358 211148 128360 211168
rect 128360 211148 128412 211168
rect 128412 211148 128414 211168
rect 128358 211112 128414 211148
rect 129002 203496 129058 203552
rect 128634 195880 128690 195936
rect 453302 288088 453358 288144
rect 453026 252456 453082 252512
rect 453118 231104 453174 231160
rect 580170 310800 580226 310856
rect 453670 302388 453726 302424
rect 453670 302368 453672 302388
rect 453672 302368 453724 302388
rect 453724 302368 453726 302388
rect 453946 281016 454002 281072
rect 453670 273808 453726 273864
rect 453578 266736 453634 266792
rect 453486 245384 453542 245440
rect 453394 224032 453450 224088
rect 453302 202680 453358 202736
rect 2778 7112 2834 7168
rect 143998 183504 144054 183560
rect 144182 183504 144238 183560
rect 143630 154536 143686 154592
rect 143906 154536 143962 154592
rect 143630 115912 143686 115968
rect 143906 115912 143962 115968
rect 143630 96600 143686 96656
rect 143906 96600 143962 96656
rect 453946 259664 454002 259720
rect 579802 299104 579858 299160
rect 453946 238312 454002 238368
rect 453762 216960 453818 217016
rect 453946 209788 453948 209808
rect 453948 209788 454000 209808
rect 454000 209788 454002 209808
rect 453946 209752 454002 209788
rect 453946 195608 454002 195664
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 542353 683226 542419 683229
rect 542721 683226 542787 683229
rect 542353 683224 542787 683226
rect 542353 683168 542358 683224
rect 542414 683168 542726 683224
rect 542782 683168 542787 683224
rect 542353 683166 542787 683168
rect 542353 683163 542419 683166
rect 542721 683163 542787 683166
rect -960 682274 480 682364
rect 3325 682274 3391 682277
rect -960 682272 3391 682274
rect -960 682216 3330 682272
rect 3386 682216 3391 682272
rect -960 682214 3391 682216
rect -960 682124 480 682214
rect 3325 682211 3391 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3233 624882 3299 624885
rect -960 624880 3299 624882
rect -960 624824 3238 624880
rect 3294 624824 3299 624880
rect -960 624822 3299 624824
rect -960 624732 480 624822
rect 3233 624819 3299 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3509 610466 3575 610469
rect -960 610464 3575 610466
rect -960 610408 3514 610464
rect 3570 610408 3575 610464
rect -960 610406 3575 610408
rect -960 610316 480 610406
rect 3509 610403 3575 610406
rect 72969 608562 73035 608565
rect 73153 608562 73219 608565
rect 72969 608560 73219 608562
rect 72969 608504 72974 608560
rect 73030 608504 73158 608560
rect 73214 608504 73219 608560
rect 72969 608502 73219 608504
rect 72969 608499 73035 608502
rect 73153 608499 73219 608502
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 579889 592514 579955 592517
rect 583520 592514 584960 592604
rect 579889 592512 584960 592514
rect 579889 592456 579894 592512
rect 579950 592456 584960 592512
rect 579889 592454 584960 592456
rect 579889 592451 579955 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 347865 560282 347931 560285
rect 348049 560282 348115 560285
rect 347865 560280 348115 560282
rect 347865 560224 347870 560280
rect 347926 560224 348054 560280
rect 348110 560224 348115 560280
rect 347865 560222 348115 560224
rect 347865 560219 347931 560222
rect 348049 560219 348115 560222
rect 364425 560282 364491 560285
rect 364609 560282 364675 560285
rect 364425 560280 364675 560282
rect 364425 560224 364430 560280
rect 364486 560224 364614 560280
rect 364670 560224 364675 560280
rect 364425 560222 364675 560224
rect 364425 560219 364491 560222
rect 364609 560219 364675 560222
rect 477585 560282 477651 560285
rect 477769 560282 477835 560285
rect 477585 560280 477835 560282
rect 477585 560224 477590 560280
rect 477646 560224 477774 560280
rect 477830 560224 477835 560280
rect 477585 560222 477835 560224
rect 477585 560219 477651 560222
rect 477769 560219 477835 560222
rect 494145 560282 494211 560285
rect 494329 560282 494395 560285
rect 494145 560280 494395 560282
rect 494145 560224 494150 560280
rect 494206 560224 494334 560280
rect 494390 560224 494395 560280
rect 494145 560222 494395 560224
rect 494145 560219 494211 560222
rect 494329 560219 494395 560222
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3601 553074 3667 553077
rect -960 553072 3667 553074
rect -960 553016 3606 553072
rect 3662 553016 3667 553072
rect -960 553014 3667 553016
rect -960 552924 480 553014
rect 3601 553011 3667 553014
rect 579889 545594 579955 545597
rect 583520 545594 584960 545684
rect 579889 545592 584960 545594
rect 579889 545536 579894 545592
rect 579950 545536 584960 545592
rect 579889 545534 584960 545536
rect 579889 545531 579955 545534
rect 583520 545444 584960 545534
rect 8201 540970 8267 540973
rect 8385 540970 8451 540973
rect 8201 540968 8451 540970
rect 8201 540912 8206 540968
rect 8262 540912 8390 540968
rect 8446 540912 8451 540968
rect 8201 540910 8451 540912
rect 8201 540907 8267 540910
rect 8385 540907 8451 540910
rect 154205 540970 154271 540973
rect 154481 540970 154547 540973
rect 154205 540968 154547 540970
rect 154205 540912 154210 540968
rect 154266 540912 154486 540968
rect 154542 540912 154547 540968
rect 154205 540910 154547 540912
rect 154205 540907 154271 540910
rect 154481 540907 154547 540910
rect 284201 540970 284267 540973
rect 284385 540970 284451 540973
rect 284201 540968 284451 540970
rect 284201 540912 284206 540968
rect 284262 540912 284390 540968
rect 284446 540912 284451 540968
rect 284201 540910 284451 540912
rect 284201 540907 284267 540910
rect 284385 540907 284451 540910
rect 347865 540970 347931 540973
rect 348049 540970 348115 540973
rect 347865 540968 348115 540970
rect 347865 540912 347870 540968
rect 347926 540912 348054 540968
rect 348110 540912 348115 540968
rect 347865 540910 348115 540912
rect 347865 540907 347931 540910
rect 348049 540907 348115 540910
rect 364425 540970 364491 540973
rect 364609 540970 364675 540973
rect 364425 540968 364675 540970
rect 364425 540912 364430 540968
rect 364486 540912 364614 540968
rect 364670 540912 364675 540968
rect 364425 540910 364675 540912
rect 364425 540907 364491 540910
rect 364609 540907 364675 540910
rect 477585 540970 477651 540973
rect 477769 540970 477835 540973
rect 477585 540968 477835 540970
rect 477585 540912 477590 540968
rect 477646 540912 477774 540968
rect 477830 540912 477835 540968
rect 477585 540910 477835 540912
rect 477585 540907 477651 540910
rect 477769 540907 477835 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -960 538658 480 538748
rect 3693 538658 3759 538661
rect -960 538656 3759 538658
rect -960 538600 3698 538656
rect 3754 538600 3759 538656
rect -960 538598 3759 538600
rect -960 538508 480 538598
rect 3693 538595 3759 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 8109 531314 8175 531317
rect 8293 531314 8359 531317
rect 8109 531312 8359 531314
rect 8109 531256 8114 531312
rect 8170 531256 8298 531312
rect 8354 531256 8359 531312
rect 8109 531254 8359 531256
rect 8109 531251 8175 531254
rect 8293 531251 8359 531254
rect 284109 531314 284175 531317
rect 284293 531314 284359 531317
rect 284109 531312 284359 531314
rect 284109 531256 284114 531312
rect 284170 531256 284298 531312
rect 284354 531256 284359 531312
rect 284109 531254 284359 531256
rect 284109 531251 284175 531254
rect 284293 531251 284359 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3233 509962 3299 509965
rect -960 509960 3299 509962
rect -960 509904 3238 509960
rect 3294 509904 3299 509960
rect -960 509902 3299 509904
rect -960 509812 480 509902
rect 3233 509899 3299 509902
rect 453205 508874 453271 508877
rect 450156 508872 453271 508874
rect 450156 508816 453210 508872
rect 453266 508816 453271 508872
rect 450156 508814 453271 508816
rect 453205 508811 453271 508814
rect 128353 508602 128419 508605
rect 128353 508600 132020 508602
rect 128353 508544 128358 508600
rect 128414 508544 132020 508600
rect 128353 508542 132020 508544
rect 128353 508539 128419 508542
rect 453389 501802 453455 501805
rect 450156 501800 453455 501802
rect 450156 501744 453394 501800
rect 453450 501744 453455 501800
rect 450156 501742 453455 501744
rect 453389 501739 453455 501742
rect 128353 500986 128419 500989
rect 128353 500984 132020 500986
rect 128353 500928 128358 500984
rect 128414 500928 132020 500984
rect 128353 500926 132020 500928
rect 128353 500923 128419 500926
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 453941 494594 454007 494597
rect 450156 494592 454007 494594
rect 450156 494536 453946 494592
rect 454002 494536 454007 494592
rect 450156 494534 454007 494536
rect 453941 494531 454007 494534
rect 128997 493370 129063 493373
rect 128997 493368 132020 493370
rect 128997 493312 129002 493368
rect 129058 493312 132020 493368
rect 128997 493310 132020 493312
rect 128997 493307 129063 493310
rect 453757 487522 453823 487525
rect 450156 487520 453823 487522
rect 450156 487464 453762 487520
rect 453818 487464 453823 487520
rect 450156 487462 453823 487464
rect 453757 487459 453823 487462
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 128353 485754 128419 485757
rect 128353 485752 132020 485754
rect 128353 485696 128358 485752
rect 128414 485696 132020 485752
rect 128353 485694 132020 485696
rect 128353 485691 128419 485694
rect -960 481130 480 481220
rect 3785 481130 3851 481133
rect -960 481128 3851 481130
rect -960 481072 3790 481128
rect 3846 481072 3851 481128
rect -960 481070 3851 481072
rect -960 480980 480 481070
rect 3785 481067 3851 481070
rect 453757 480450 453823 480453
rect 450156 480448 453823 480450
rect 450156 480392 453762 480448
rect 453818 480392 453823 480448
rect 450156 480390 453823 480392
rect 453757 480387 453823 480390
rect 128353 478138 128419 478141
rect 128353 478136 132020 478138
rect 128353 478080 128358 478136
rect 128414 478080 132020 478136
rect 128353 478078 132020 478080
rect 128353 478075 128419 478078
rect 583520 474996 584960 475236
rect 453941 473242 454007 473245
rect 450156 473240 454007 473242
rect 450156 473184 453946 473240
rect 454002 473184 454007 473240
rect 450156 473182 454007 473184
rect 453941 473179 454007 473182
rect 128353 470522 128419 470525
rect 128353 470520 132020 470522
rect 128353 470464 128358 470520
rect 128414 470464 132020 470520
rect 128353 470462 132020 470464
rect 128353 470459 128419 470462
rect -960 466700 480 466940
rect 452745 466170 452811 466173
rect 450156 466168 452811 466170
rect 450156 466112 452750 466168
rect 452806 466112 452811 466168
rect 450156 466110 452811 466112
rect 452745 466107 452811 466110
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 128353 462906 128419 462909
rect 128353 462904 132020 462906
rect 128353 462848 128358 462904
rect 128414 462848 132020 462904
rect 128353 462846 132020 462848
rect 128353 462843 128419 462846
rect 453389 459098 453455 459101
rect 450156 459096 453455 459098
rect 450156 459040 453394 459096
rect 453450 459040 453455 459096
rect 450156 459038 453455 459040
rect 453389 459035 453455 459038
rect 128353 455290 128419 455293
rect 128353 455288 132020 455290
rect 128353 455232 128358 455288
rect 128414 455232 132020 455288
rect 128353 455230 132020 455232
rect 128353 455227 128419 455230
rect -960 452434 480 452524
rect 3509 452434 3575 452437
rect -960 452432 3575 452434
rect -960 452376 3514 452432
rect 3570 452376 3575 452432
rect -960 452374 3575 452376
rect -960 452284 480 452374
rect 3509 452371 3575 452374
rect 453941 451890 454007 451893
rect 450156 451888 454007 451890
rect 450156 451832 453946 451888
rect 454002 451832 454007 451888
rect 450156 451830 454007 451832
rect 453941 451827 454007 451830
rect 580257 451754 580323 451757
rect 583520 451754 584960 451844
rect 580257 451752 584960 451754
rect 580257 451696 580262 451752
rect 580318 451696 584960 451752
rect 580257 451694 584960 451696
rect 580257 451691 580323 451694
rect 583520 451604 584960 451694
rect 128353 447674 128419 447677
rect 128353 447672 132020 447674
rect 128353 447616 128358 447672
rect 128414 447616 132020 447672
rect 128353 447614 132020 447616
rect 128353 447611 128419 447614
rect 453665 444818 453731 444821
rect 450156 444816 453731 444818
rect 450156 444760 453670 444816
rect 453726 444760 453731 444816
rect 450156 444758 453731 444760
rect 453665 444755 453731 444758
rect 128353 440058 128419 440061
rect 128353 440056 132020 440058
rect 128353 440000 128358 440056
rect 128414 440000 132020 440056
rect 128353 439998 132020 440000
rect 128353 439995 128419 439998
rect 579889 439922 579955 439925
rect 583520 439922 584960 440012
rect 579889 439920 584960 439922
rect 579889 439864 579894 439920
rect 579950 439864 584960 439920
rect 579889 439862 584960 439864
rect 579889 439859 579955 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3601 438018 3667 438021
rect -960 438016 3667 438018
rect -960 437960 3606 438016
rect 3662 437960 3667 438016
rect -960 437958 3667 437960
rect -960 437868 480 437958
rect 3601 437955 3667 437958
rect 453757 437746 453823 437749
rect 450156 437744 453823 437746
rect 450156 437688 453762 437744
rect 453818 437688 453823 437744
rect 450156 437686 453823 437688
rect 453757 437683 453823 437686
rect 128353 432306 128419 432309
rect 128353 432304 132020 432306
rect 128353 432248 128358 432304
rect 128414 432248 132020 432304
rect 128353 432246 132020 432248
rect 128353 432243 128419 432246
rect 453941 430538 454007 430541
rect 450156 430536 454007 430538
rect 450156 430480 453946 430536
rect 454002 430480 454007 430536
rect 450156 430478 454007 430480
rect 453941 430475 454007 430478
rect 583520 428076 584960 428316
rect 128353 424690 128419 424693
rect 128353 424688 132020 424690
rect 128353 424632 128358 424688
rect 128414 424632 132020 424688
rect 128353 424630 132020 424632
rect 128353 424627 128419 424630
rect -960 423738 480 423828
rect 3417 423738 3483 423741
rect -960 423736 3483 423738
rect -960 423680 3422 423736
rect 3478 423680 3483 423736
rect -960 423678 3483 423680
rect -960 423588 480 423678
rect 3417 423675 3483 423678
rect 453941 423466 454007 423469
rect 450156 423464 454007 423466
rect 450156 423408 453946 423464
rect 454002 423408 454007 423464
rect 450156 423406 454007 423408
rect 453941 423403 454007 423406
rect 128353 417074 128419 417077
rect 128353 417072 132020 417074
rect 128353 417016 128358 417072
rect 128414 417016 132020 417072
rect 128353 417014 132020 417016
rect 128353 417011 128419 417014
rect 578877 416530 578943 416533
rect 583520 416530 584960 416620
rect 578877 416528 584960 416530
rect 578877 416472 578882 416528
rect 578938 416472 584960 416528
rect 578877 416470 584960 416472
rect 578877 416467 578943 416470
rect 453941 416394 454007 416397
rect 450156 416392 454007 416394
rect 450156 416336 453946 416392
rect 454002 416336 454007 416392
rect 583520 416380 584960 416470
rect 450156 416334 454007 416336
rect 453941 416331 454007 416334
rect 128353 409458 128419 409461
rect 128353 409456 132020 409458
rect -960 409172 480 409412
rect 128353 409400 128358 409456
rect 128414 409400 132020 409456
rect 128353 409398 132020 409400
rect 128353 409395 128419 409398
rect 453389 409186 453455 409189
rect 450156 409184 453455 409186
rect 450156 409128 453394 409184
rect 453450 409128 453455 409184
rect 450156 409126 453455 409128
rect 453389 409123 453455 409126
rect 580349 404834 580415 404837
rect 583520 404834 584960 404924
rect 580349 404832 584960 404834
rect 580349 404776 580354 404832
rect 580410 404776 584960 404832
rect 580349 404774 584960 404776
rect 580349 404771 580415 404774
rect 583520 404684 584960 404774
rect 453941 402114 454007 402117
rect 450156 402112 454007 402114
rect 450156 402056 453946 402112
rect 454002 402056 454007 402112
rect 450156 402054 454007 402056
rect 453941 402051 454007 402054
rect 128353 401842 128419 401845
rect 128353 401840 132020 401842
rect 128353 401784 128358 401840
rect 128414 401784 132020 401840
rect 128353 401782 132020 401784
rect 128353 401779 128419 401782
rect -960 395042 480 395132
rect 3417 395042 3483 395045
rect -960 395040 3483 395042
rect -960 394984 3422 395040
rect 3478 394984 3483 395040
rect -960 394982 3483 394984
rect -960 394892 480 394982
rect 3417 394979 3483 394982
rect 453757 394906 453823 394909
rect 450156 394904 453823 394906
rect 450156 394848 453762 394904
rect 453818 394848 453823 394904
rect 450156 394846 453823 394848
rect 453757 394843 453823 394846
rect 128353 394226 128419 394229
rect 128353 394224 132020 394226
rect 128353 394168 128358 394224
rect 128414 394168 132020 394224
rect 128353 394166 132020 394168
rect 128353 394163 128419 394166
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 453297 387834 453363 387837
rect 450156 387832 453363 387834
rect 450156 387776 453302 387832
rect 453358 387776 453363 387832
rect 450156 387774 453363 387776
rect 453297 387771 453363 387774
rect 128997 386610 129063 386613
rect 128997 386608 132020 386610
rect 128997 386552 129002 386608
rect 129058 386552 132020 386608
rect 128997 386550 132020 386552
rect 128997 386547 129063 386550
rect 583520 381156 584960 381396
rect 453941 380762 454007 380765
rect 450156 380760 454007 380762
rect -960 380626 480 380716
rect 450156 380704 453946 380760
rect 454002 380704 454007 380760
rect 450156 380702 454007 380704
rect 453941 380699 454007 380702
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 128997 378994 129063 378997
rect 128997 378992 132020 378994
rect 128997 378936 129002 378992
rect 129058 378936 132020 378992
rect 128997 378934 132020 378936
rect 128997 378931 129063 378934
rect 453389 373554 453455 373557
rect 450156 373552 453455 373554
rect 450156 373496 453394 373552
rect 453450 373496 453455 373552
rect 450156 373494 453455 373496
rect 453389 373491 453455 373494
rect 129273 371378 129339 371381
rect 129273 371376 132020 371378
rect 129273 371320 129278 371376
rect 129334 371320 132020 371376
rect 129273 371318 132020 371320
rect 129273 371315 129339 371318
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 583520 369460 584960 369550
rect 453941 366482 454007 366485
rect 450156 366480 454007 366482
rect 450156 366424 453946 366480
rect 454002 366424 454007 366480
rect 450156 366422 454007 366424
rect 453941 366419 454007 366422
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 128997 363762 129063 363765
rect 128997 363760 132020 363762
rect 128997 363704 129002 363760
rect 129058 363704 132020 363760
rect 128997 363702 132020 363704
rect 128997 363699 129063 363702
rect 453941 359410 454007 359413
rect 450156 359408 454007 359410
rect 450156 359352 453946 359408
rect 454002 359352 454007 359408
rect 450156 359350 454007 359352
rect 453941 359347 454007 359350
rect 580257 357914 580323 357917
rect 583520 357914 584960 358004
rect 580257 357912 584960 357914
rect 580257 357856 580262 357912
rect 580318 357856 584960 357912
rect 580257 357854 584960 357856
rect 580257 357851 580323 357854
rect 583520 357764 584960 357854
rect 129181 356146 129247 356149
rect 129181 356144 132020 356146
rect 129181 356088 129186 356144
rect 129242 356088 132020 356144
rect 129181 356086 132020 356088
rect 129181 356083 129247 356086
rect 453757 352202 453823 352205
rect 450156 352200 453823 352202
rect 450156 352144 453762 352200
rect 453818 352144 453823 352200
rect 450156 352142 453823 352144
rect 453757 352139 453823 352142
rect -960 351780 480 352020
rect 128353 348394 128419 348397
rect 128353 348392 132020 348394
rect 128353 348336 128358 348392
rect 128414 348336 132020 348392
rect 128353 348334 132020 348336
rect 128353 348331 128419 348334
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 453941 345130 454007 345133
rect 450156 345128 454007 345130
rect 450156 345072 453946 345128
rect 454002 345072 454007 345128
rect 450156 345070 454007 345072
rect 453941 345067 454007 345070
rect 129089 340778 129155 340781
rect 129089 340776 132020 340778
rect 129089 340720 129094 340776
rect 129150 340720 132020 340776
rect 129089 340718 132020 340720
rect 129089 340715 129155 340718
rect 453481 338058 453547 338061
rect 450156 338056 453547 338058
rect 450156 338000 453486 338056
rect 453542 338000 453547 338056
rect 450156 337998 453547 338000
rect 453481 337995 453547 337998
rect -960 337514 480 337604
rect 3509 337514 3575 337517
rect -960 337512 3575 337514
rect -960 337456 3514 337512
rect 3570 337456 3575 337512
rect -960 337454 3575 337456
rect -960 337364 480 337454
rect 3509 337451 3575 337454
rect 583520 334236 584960 334476
rect 128353 333162 128419 333165
rect 128353 333160 132020 333162
rect 128353 333104 128358 333160
rect 128414 333104 132020 333160
rect 128353 333102 132020 333104
rect 128353 333099 128419 333102
rect 453389 330850 453455 330853
rect 450156 330848 453455 330850
rect 450156 330792 453394 330848
rect 453450 330792 453455 330848
rect 450156 330790 453455 330792
rect 453389 330787 453455 330790
rect 128353 325546 128419 325549
rect 128353 325544 132020 325546
rect 128353 325488 128358 325544
rect 128414 325488 132020 325544
rect 128353 325486 132020 325488
rect 128353 325483 128419 325486
rect 453297 323778 453363 323781
rect 450156 323776 453363 323778
rect 450156 323720 453302 323776
rect 453358 323720 453363 323776
rect 450156 323718 453363 323720
rect 453297 323715 453363 323718
rect -960 323098 480 323188
rect 3509 323098 3575 323101
rect -960 323096 3575 323098
rect -960 323040 3514 323096
rect 3570 323040 3575 323096
rect -960 323038 3575 323040
rect -960 322948 480 323038
rect 3509 323035 3575 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 128997 317930 129063 317933
rect 128997 317928 132020 317930
rect 128997 317872 129002 317928
rect 129058 317872 132020 317928
rect 128997 317870 132020 317872
rect 128997 317867 129063 317870
rect 453573 316706 453639 316709
rect 450156 316704 453639 316706
rect 450156 316648 453578 316704
rect 453634 316648 453639 316704
rect 450156 316646 453639 316648
rect 453573 316643 453639 316646
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 128353 310314 128419 310317
rect 128353 310312 132020 310314
rect 128353 310256 128358 310312
rect 128414 310256 132020 310312
rect 128353 310254 132020 310256
rect 128353 310251 128419 310254
rect 453481 309498 453547 309501
rect 450156 309496 453547 309498
rect 450156 309440 453486 309496
rect 453542 309440 453547 309496
rect 450156 309438 453547 309440
rect 453481 309435 453547 309438
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 128353 302698 128419 302701
rect 128353 302696 132020 302698
rect 128353 302640 128358 302696
rect 128414 302640 132020 302696
rect 128353 302638 132020 302640
rect 128353 302635 128419 302638
rect 453665 302426 453731 302429
rect 450156 302424 453731 302426
rect 450156 302368 453670 302424
rect 453726 302368 453731 302424
rect 450156 302366 453731 302368
rect 453665 302363 453731 302366
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 453389 295218 453455 295221
rect 450156 295216 453455 295218
rect 450156 295160 453394 295216
rect 453450 295160 453455 295216
rect 450156 295158 453455 295160
rect 453389 295155 453455 295158
rect 129365 295082 129431 295085
rect 129365 295080 132020 295082
rect 129365 295024 129370 295080
rect 129426 295024 132020 295080
rect 129365 295022 132020 295024
rect 129365 295019 129431 295022
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 453297 288146 453363 288149
rect 450156 288144 453363 288146
rect 450156 288088 453302 288144
rect 453358 288088 453363 288144
rect 450156 288086 453363 288088
rect 453297 288083 453363 288086
rect 128353 287466 128419 287469
rect 128353 287464 132020 287466
rect 128353 287408 128358 287464
rect 128414 287408 132020 287464
rect 128353 287406 132020 287408
rect 128353 287403 128419 287406
rect 583520 287316 584960 287556
rect 453941 281074 454007 281077
rect 450156 281072 454007 281074
rect 450156 281016 453946 281072
rect 454002 281016 454007 281072
rect 450156 281014 454007 281016
rect 453941 281011 454007 281014
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 128261 279850 128327 279853
rect 128261 279848 132020 279850
rect 128261 279792 128266 279848
rect 128322 279792 132020 279848
rect 128261 279790 132020 279792
rect 128261 279787 128327 279790
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 453665 273866 453731 273869
rect 450156 273864 453731 273866
rect 450156 273808 453670 273864
rect 453726 273808 453731 273864
rect 450156 273806 453731 273808
rect 453665 273803 453731 273806
rect 129273 272098 129339 272101
rect 129273 272096 132020 272098
rect 129273 272040 129278 272096
rect 129334 272040 132020 272096
rect 129273 272038 132020 272040
rect 129273 272035 129339 272038
rect 453573 266794 453639 266797
rect 450156 266792 453639 266794
rect 450156 266736 453578 266792
rect 453634 266736 453639 266792
rect 450156 266734 453639 266736
rect 453573 266731 453639 266734
rect -960 265706 480 265796
rect 3509 265706 3575 265709
rect -960 265704 3575 265706
rect -960 265648 3514 265704
rect 3570 265648 3575 265704
rect -960 265646 3575 265648
rect -960 265556 480 265646
rect 3509 265643 3575 265646
rect 128353 264482 128419 264485
rect 128353 264480 132020 264482
rect 128353 264424 128358 264480
rect 128414 264424 132020 264480
rect 128353 264422 132020 264424
rect 128353 264419 128419 264422
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 453941 259722 454007 259725
rect 450156 259720 454007 259722
rect 450156 259664 453946 259720
rect 454002 259664 454007 259720
rect 450156 259662 454007 259664
rect 453941 259659 454007 259662
rect 128353 256866 128419 256869
rect 128353 256864 132020 256866
rect 128353 256808 128358 256864
rect 128414 256808 132020 256864
rect 128353 256806 132020 256808
rect 128353 256803 128419 256806
rect 453021 252514 453087 252517
rect 450156 252512 453087 252514
rect 450156 252456 453026 252512
rect 453082 252456 453087 252512
rect 450156 252454 453087 252456
rect 453021 252451 453087 252454
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3509 251290 3575 251293
rect -960 251288 3575 251290
rect -960 251232 3514 251288
rect 3570 251232 3575 251288
rect -960 251230 3575 251232
rect -960 251140 480 251230
rect 3509 251227 3575 251230
rect 129181 249250 129247 249253
rect 129181 249248 132020 249250
rect 129181 249192 129186 249248
rect 129242 249192 132020 249248
rect 129181 249190 132020 249192
rect 129181 249187 129247 249190
rect 453481 245442 453547 245445
rect 450156 245440 453547 245442
rect 450156 245384 453486 245440
rect 453542 245384 453547 245440
rect 450156 245382 453547 245384
rect 453481 245379 453547 245382
rect 128353 241634 128419 241637
rect 128353 241632 132020 241634
rect 128353 241576 128358 241632
rect 128414 241576 132020 241632
rect 128353 241574 132020 241576
rect 128353 241571 128419 241574
rect 583520 240396 584960 240636
rect 453941 238370 454007 238373
rect 450156 238368 454007 238370
rect 450156 238312 453946 238368
rect 454002 238312 454007 238368
rect 450156 238310 454007 238312
rect 453941 238307 454007 238310
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 128353 234018 128419 234021
rect 128353 234016 132020 234018
rect 128353 233960 128358 234016
rect 128414 233960 132020 234016
rect 128353 233958 132020 233960
rect 128353 233955 128419 233958
rect 453113 231162 453179 231165
rect 450156 231160 453179 231162
rect 450156 231104 453118 231160
rect 453174 231104 453179 231160
rect 450156 231102 453179 231104
rect 453113 231099 453179 231102
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 129089 226402 129155 226405
rect 129089 226400 132020 226402
rect 129089 226344 129094 226400
rect 129150 226344 132020 226400
rect 129089 226342 132020 226344
rect 129089 226339 129155 226342
rect 453389 224090 453455 224093
rect 450156 224088 453455 224090
rect 450156 224032 453394 224088
rect 453450 224032 453455 224088
rect 450156 224030 453455 224032
rect 453389 224027 453455 224030
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 128353 218786 128419 218789
rect 128353 218784 132020 218786
rect 128353 218728 128358 218784
rect 128414 218728 132020 218784
rect 128353 218726 132020 218728
rect 128353 218723 128419 218726
rect 453757 217018 453823 217021
rect 450156 217016 453823 217018
rect 450156 216960 453762 217016
rect 453818 216960 453823 217016
rect 450156 216958 453823 216960
rect 453757 216955 453823 216958
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 128353 211170 128419 211173
rect 128353 211168 132020 211170
rect 128353 211112 128358 211168
rect 128414 211112 132020 211168
rect 128353 211110 132020 211112
rect 128353 211107 128419 211110
rect 453941 209810 454007 209813
rect 450156 209808 454007 209810
rect 450156 209752 453946 209808
rect 454002 209752 454007 209808
rect 450156 209750 454007 209752
rect 453941 209747 454007 209750
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 128997 203554 129063 203557
rect 128997 203552 132020 203554
rect 128997 203496 129002 203552
rect 129058 203496 132020 203552
rect 128997 203494 132020 203496
rect 128997 203491 129063 203494
rect 453297 202738 453363 202741
rect 450156 202736 453363 202738
rect 450156 202680 453302 202736
rect 453358 202680 453363 202736
rect 450156 202678 453363 202680
rect 453297 202675 453363 202678
rect 128629 195938 128695 195941
rect 128629 195936 132020 195938
rect 128629 195880 128634 195936
rect 128690 195880 132020 195936
rect 128629 195878 132020 195880
rect 128629 195875 128695 195878
rect 453941 195666 454007 195669
rect 450156 195664 454007 195666
rect 450156 195608 453946 195664
rect 454002 195608 454007 195664
rect 450156 195606 454007 195608
rect 453941 195603 454007 195606
rect -960 193898 480 193988
rect 2865 193898 2931 193901
rect -960 193896 2931 193898
rect -960 193840 2870 193896
rect 2926 193840 2931 193896
rect -960 193838 2931 193840
rect -960 193748 480 193838
rect 2865 193835 2931 193838
rect 583520 193476 584960 193716
rect 143993 183562 144059 183565
rect 144177 183562 144243 183565
rect 143993 183560 144243 183562
rect 143993 183504 143998 183560
rect 144054 183504 144182 183560
rect 144238 183504 144243 183560
rect 143993 183502 144243 183504
rect 143993 183499 144059 183502
rect 144177 183499 144243 183502
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3417 165066 3483 165069
rect -960 165064 3483 165066
rect -960 165008 3422 165064
rect 3478 165008 3483 165064
rect -960 165006 3483 165008
rect -960 164916 480 165006
rect 3417 165003 3483 165006
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 143625 154594 143691 154597
rect 143901 154594 143967 154597
rect 143625 154592 143967 154594
rect 143625 154536 143630 154592
rect 143686 154536 143906 154592
rect 143962 154536 143967 154592
rect 143625 154534 143967 154536
rect 143625 154531 143691 154534
rect 143901 154531 143967 154534
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3417 136370 3483 136373
rect -960 136368 3483 136370
rect -960 136312 3422 136368
rect 3478 136312 3483 136368
rect -960 136310 3483 136312
rect -960 136220 480 136310
rect 3417 136307 3483 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 143625 115970 143691 115973
rect 143901 115970 143967 115973
rect 143625 115968 143967 115970
rect 143625 115912 143630 115968
rect 143686 115912 143906 115968
rect 143962 115912 143967 115968
rect 143625 115910 143967 115912
rect 143625 115907 143691 115910
rect 143901 115907 143967 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect 143625 96658 143691 96661
rect 143901 96658 143967 96661
rect 143625 96656 143967 96658
rect 143625 96600 143630 96656
rect 143686 96600 143906 96656
rect 143962 96600 143967 96656
rect 143625 96598 143967 96600
rect 143625 96595 143691 96598
rect 143901 96595 143967 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 2773 7170 2839 7173
rect -960 7168 2839 7170
rect -960 7112 2778 7168
rect 2834 7112 2839 7168
rect -960 7110 2839 7112
rect -960 7020 480 7110
rect 2773 7107 2839 7110
rect 583520 5796 584960 6036
<< metal4 >>
rect -4876 707718 -4276 707740
rect -4876 707482 -4694 707718
rect -4458 707482 -4276 707718
rect -4876 707398 -4276 707482
rect -4876 707162 -4694 707398
rect -4458 707162 -4276 707398
rect -4876 672054 -4276 707162
rect -4876 671818 -4694 672054
rect -4458 671818 -4276 672054
rect -4876 671734 -4276 671818
rect -4876 671498 -4694 671734
rect -4458 671498 -4276 671734
rect -4876 636054 -4276 671498
rect -4876 635818 -4694 636054
rect -4458 635818 -4276 636054
rect -4876 635734 -4276 635818
rect -4876 635498 -4694 635734
rect -4458 635498 -4276 635734
rect -4876 600054 -4276 635498
rect -4876 599818 -4694 600054
rect -4458 599818 -4276 600054
rect -4876 599734 -4276 599818
rect -4876 599498 -4694 599734
rect -4458 599498 -4276 599734
rect -4876 564054 -4276 599498
rect -4876 563818 -4694 564054
rect -4458 563818 -4276 564054
rect -4876 563734 -4276 563818
rect -4876 563498 -4694 563734
rect -4458 563498 -4276 563734
rect -4876 528054 -4276 563498
rect -4876 527818 -4694 528054
rect -4458 527818 -4276 528054
rect -4876 527734 -4276 527818
rect -4876 527498 -4694 527734
rect -4458 527498 -4276 527734
rect -4876 492054 -4276 527498
rect -4876 491818 -4694 492054
rect -4458 491818 -4276 492054
rect -4876 491734 -4276 491818
rect -4876 491498 -4694 491734
rect -4458 491498 -4276 491734
rect -4876 456054 -4276 491498
rect -4876 455818 -4694 456054
rect -4458 455818 -4276 456054
rect -4876 455734 -4276 455818
rect -4876 455498 -4694 455734
rect -4458 455498 -4276 455734
rect -4876 420054 -4276 455498
rect -4876 419818 -4694 420054
rect -4458 419818 -4276 420054
rect -4876 419734 -4276 419818
rect -4876 419498 -4694 419734
rect -4458 419498 -4276 419734
rect -4876 384054 -4276 419498
rect -4876 383818 -4694 384054
rect -4458 383818 -4276 384054
rect -4876 383734 -4276 383818
rect -4876 383498 -4694 383734
rect -4458 383498 -4276 383734
rect -4876 348054 -4276 383498
rect -4876 347818 -4694 348054
rect -4458 347818 -4276 348054
rect -4876 347734 -4276 347818
rect -4876 347498 -4694 347734
rect -4458 347498 -4276 347734
rect -4876 312054 -4276 347498
rect -4876 311818 -4694 312054
rect -4458 311818 -4276 312054
rect -4876 311734 -4276 311818
rect -4876 311498 -4694 311734
rect -4458 311498 -4276 311734
rect -4876 276054 -4276 311498
rect -4876 275818 -4694 276054
rect -4458 275818 -4276 276054
rect -4876 275734 -4276 275818
rect -4876 275498 -4694 275734
rect -4458 275498 -4276 275734
rect -4876 240054 -4276 275498
rect -4876 239818 -4694 240054
rect -4458 239818 -4276 240054
rect -4876 239734 -4276 239818
rect -4876 239498 -4694 239734
rect -4458 239498 -4276 239734
rect -4876 204054 -4276 239498
rect -4876 203818 -4694 204054
rect -4458 203818 -4276 204054
rect -4876 203734 -4276 203818
rect -4876 203498 -4694 203734
rect -4458 203498 -4276 203734
rect -4876 168054 -4276 203498
rect -4876 167818 -4694 168054
rect -4458 167818 -4276 168054
rect -4876 167734 -4276 167818
rect -4876 167498 -4694 167734
rect -4458 167498 -4276 167734
rect -4876 132054 -4276 167498
rect -4876 131818 -4694 132054
rect -4458 131818 -4276 132054
rect -4876 131734 -4276 131818
rect -4876 131498 -4694 131734
rect -4458 131498 -4276 131734
rect -4876 96054 -4276 131498
rect -4876 95818 -4694 96054
rect -4458 95818 -4276 96054
rect -4876 95734 -4276 95818
rect -4876 95498 -4694 95734
rect -4458 95498 -4276 95734
rect -4876 60054 -4276 95498
rect -4876 59818 -4694 60054
rect -4458 59818 -4276 60054
rect -4876 59734 -4276 59818
rect -4876 59498 -4694 59734
rect -4458 59498 -4276 59734
rect -4876 24054 -4276 59498
rect -4876 23818 -4694 24054
rect -4458 23818 -4276 24054
rect -4876 23734 -4276 23818
rect -4876 23498 -4694 23734
rect -4458 23498 -4276 23734
rect -4876 -3226 -4276 23498
rect -3916 706758 -3316 706780
rect -3916 706522 -3734 706758
rect -3498 706522 -3316 706758
rect -3916 706438 -3316 706522
rect -3916 706202 -3734 706438
rect -3498 706202 -3316 706438
rect -3916 690054 -3316 706202
rect 4404 706758 5004 707740
rect 4404 706522 4586 706758
rect 4822 706522 5004 706758
rect 4404 706438 5004 706522
rect 4404 706202 4586 706438
rect 4822 706202 5004 706438
rect -3916 689818 -3734 690054
rect -3498 689818 -3316 690054
rect -3916 689734 -3316 689818
rect -3916 689498 -3734 689734
rect -3498 689498 -3316 689734
rect -3916 654054 -3316 689498
rect -3916 653818 -3734 654054
rect -3498 653818 -3316 654054
rect -3916 653734 -3316 653818
rect -3916 653498 -3734 653734
rect -3498 653498 -3316 653734
rect -3916 618054 -3316 653498
rect -3916 617818 -3734 618054
rect -3498 617818 -3316 618054
rect -3916 617734 -3316 617818
rect -3916 617498 -3734 617734
rect -3498 617498 -3316 617734
rect -3916 582054 -3316 617498
rect -3916 581818 -3734 582054
rect -3498 581818 -3316 582054
rect -3916 581734 -3316 581818
rect -3916 581498 -3734 581734
rect -3498 581498 -3316 581734
rect -3916 546054 -3316 581498
rect -3916 545818 -3734 546054
rect -3498 545818 -3316 546054
rect -3916 545734 -3316 545818
rect -3916 545498 -3734 545734
rect -3498 545498 -3316 545734
rect -3916 510054 -3316 545498
rect -3916 509818 -3734 510054
rect -3498 509818 -3316 510054
rect -3916 509734 -3316 509818
rect -3916 509498 -3734 509734
rect -3498 509498 -3316 509734
rect -3916 474054 -3316 509498
rect -3916 473818 -3734 474054
rect -3498 473818 -3316 474054
rect -3916 473734 -3316 473818
rect -3916 473498 -3734 473734
rect -3498 473498 -3316 473734
rect -3916 438054 -3316 473498
rect -3916 437818 -3734 438054
rect -3498 437818 -3316 438054
rect -3916 437734 -3316 437818
rect -3916 437498 -3734 437734
rect -3498 437498 -3316 437734
rect -3916 402054 -3316 437498
rect -3916 401818 -3734 402054
rect -3498 401818 -3316 402054
rect -3916 401734 -3316 401818
rect -3916 401498 -3734 401734
rect -3498 401498 -3316 401734
rect -3916 366054 -3316 401498
rect -3916 365818 -3734 366054
rect -3498 365818 -3316 366054
rect -3916 365734 -3316 365818
rect -3916 365498 -3734 365734
rect -3498 365498 -3316 365734
rect -3916 330054 -3316 365498
rect -3916 329818 -3734 330054
rect -3498 329818 -3316 330054
rect -3916 329734 -3316 329818
rect -3916 329498 -3734 329734
rect -3498 329498 -3316 329734
rect -3916 294054 -3316 329498
rect -3916 293818 -3734 294054
rect -3498 293818 -3316 294054
rect -3916 293734 -3316 293818
rect -3916 293498 -3734 293734
rect -3498 293498 -3316 293734
rect -3916 258054 -3316 293498
rect -3916 257818 -3734 258054
rect -3498 257818 -3316 258054
rect -3916 257734 -3316 257818
rect -3916 257498 -3734 257734
rect -3498 257498 -3316 257734
rect -3916 222054 -3316 257498
rect -3916 221818 -3734 222054
rect -3498 221818 -3316 222054
rect -3916 221734 -3316 221818
rect -3916 221498 -3734 221734
rect -3498 221498 -3316 221734
rect -3916 186054 -3316 221498
rect -3916 185818 -3734 186054
rect -3498 185818 -3316 186054
rect -3916 185734 -3316 185818
rect -3916 185498 -3734 185734
rect -3498 185498 -3316 185734
rect -3916 150054 -3316 185498
rect -3916 149818 -3734 150054
rect -3498 149818 -3316 150054
rect -3916 149734 -3316 149818
rect -3916 149498 -3734 149734
rect -3498 149498 -3316 149734
rect -3916 114054 -3316 149498
rect -3916 113818 -3734 114054
rect -3498 113818 -3316 114054
rect -3916 113734 -3316 113818
rect -3916 113498 -3734 113734
rect -3498 113498 -3316 113734
rect -3916 78054 -3316 113498
rect -3916 77818 -3734 78054
rect -3498 77818 -3316 78054
rect -3916 77734 -3316 77818
rect -3916 77498 -3734 77734
rect -3498 77498 -3316 77734
rect -3916 42054 -3316 77498
rect -3916 41818 -3734 42054
rect -3498 41818 -3316 42054
rect -3916 41734 -3316 41818
rect -3916 41498 -3734 41734
rect -3498 41498 -3316 41734
rect -3916 6054 -3316 41498
rect -3916 5818 -3734 6054
rect -3498 5818 -3316 6054
rect -3916 5734 -3316 5818
rect -3916 5498 -3734 5734
rect -3498 5498 -3316 5734
rect -3916 -2266 -3316 5498
rect -2956 705798 -2356 705820
rect -2956 705562 -2774 705798
rect -2538 705562 -2356 705798
rect -2956 705478 -2356 705562
rect -2956 705242 -2774 705478
rect -2538 705242 -2356 705478
rect -2956 668454 -2356 705242
rect -2956 668218 -2774 668454
rect -2538 668218 -2356 668454
rect -2956 668134 -2356 668218
rect -2956 667898 -2774 668134
rect -2538 667898 -2356 668134
rect -2956 632454 -2356 667898
rect -2956 632218 -2774 632454
rect -2538 632218 -2356 632454
rect -2956 632134 -2356 632218
rect -2956 631898 -2774 632134
rect -2538 631898 -2356 632134
rect -2956 596454 -2356 631898
rect -2956 596218 -2774 596454
rect -2538 596218 -2356 596454
rect -2956 596134 -2356 596218
rect -2956 595898 -2774 596134
rect -2538 595898 -2356 596134
rect -2956 560454 -2356 595898
rect -2956 560218 -2774 560454
rect -2538 560218 -2356 560454
rect -2956 560134 -2356 560218
rect -2956 559898 -2774 560134
rect -2538 559898 -2356 560134
rect -2956 524454 -2356 559898
rect -2956 524218 -2774 524454
rect -2538 524218 -2356 524454
rect -2956 524134 -2356 524218
rect -2956 523898 -2774 524134
rect -2538 523898 -2356 524134
rect -2956 488454 -2356 523898
rect -2956 488218 -2774 488454
rect -2538 488218 -2356 488454
rect -2956 488134 -2356 488218
rect -2956 487898 -2774 488134
rect -2538 487898 -2356 488134
rect -2956 452454 -2356 487898
rect -2956 452218 -2774 452454
rect -2538 452218 -2356 452454
rect -2956 452134 -2356 452218
rect -2956 451898 -2774 452134
rect -2538 451898 -2356 452134
rect -2956 416454 -2356 451898
rect -2956 416218 -2774 416454
rect -2538 416218 -2356 416454
rect -2956 416134 -2356 416218
rect -2956 415898 -2774 416134
rect -2538 415898 -2356 416134
rect -2956 380454 -2356 415898
rect -2956 380218 -2774 380454
rect -2538 380218 -2356 380454
rect -2956 380134 -2356 380218
rect -2956 379898 -2774 380134
rect -2538 379898 -2356 380134
rect -2956 344454 -2356 379898
rect -2956 344218 -2774 344454
rect -2538 344218 -2356 344454
rect -2956 344134 -2356 344218
rect -2956 343898 -2774 344134
rect -2538 343898 -2356 344134
rect -2956 308454 -2356 343898
rect -2956 308218 -2774 308454
rect -2538 308218 -2356 308454
rect -2956 308134 -2356 308218
rect -2956 307898 -2774 308134
rect -2538 307898 -2356 308134
rect -2956 272454 -2356 307898
rect -2956 272218 -2774 272454
rect -2538 272218 -2356 272454
rect -2956 272134 -2356 272218
rect -2956 271898 -2774 272134
rect -2538 271898 -2356 272134
rect -2956 236454 -2356 271898
rect -2956 236218 -2774 236454
rect -2538 236218 -2356 236454
rect -2956 236134 -2356 236218
rect -2956 235898 -2774 236134
rect -2538 235898 -2356 236134
rect -2956 200454 -2356 235898
rect -2956 200218 -2774 200454
rect -2538 200218 -2356 200454
rect -2956 200134 -2356 200218
rect -2956 199898 -2774 200134
rect -2538 199898 -2356 200134
rect -2956 164454 -2356 199898
rect -2956 164218 -2774 164454
rect -2538 164218 -2356 164454
rect -2956 164134 -2356 164218
rect -2956 163898 -2774 164134
rect -2538 163898 -2356 164134
rect -2956 128454 -2356 163898
rect -2956 128218 -2774 128454
rect -2538 128218 -2356 128454
rect -2956 128134 -2356 128218
rect -2956 127898 -2774 128134
rect -2538 127898 -2356 128134
rect -2956 92454 -2356 127898
rect -2956 92218 -2774 92454
rect -2538 92218 -2356 92454
rect -2956 92134 -2356 92218
rect -2956 91898 -2774 92134
rect -2538 91898 -2356 92134
rect -2956 56454 -2356 91898
rect -2956 56218 -2774 56454
rect -2538 56218 -2356 56454
rect -2956 56134 -2356 56218
rect -2956 55898 -2774 56134
rect -2538 55898 -2356 56134
rect -2956 20454 -2356 55898
rect -2956 20218 -2774 20454
rect -2538 20218 -2356 20454
rect -2956 20134 -2356 20218
rect -2956 19898 -2774 20134
rect -2538 19898 -2356 20134
rect -2956 -1306 -2356 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705820
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2956 -1542 -2774 -1306
rect -2538 -1542 -2356 -1306
rect -2956 -1626 -2356 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 -2356 -1626
rect -2956 -1884 -2356 -1862
rect 804 -1884 1404 -902
rect 4404 690054 5004 706202
rect 22404 707718 23004 707740
rect 22404 707482 22586 707718
rect 22822 707482 23004 707718
rect 22404 707398 23004 707482
rect 22404 707162 22586 707398
rect 22822 707162 23004 707398
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3916 -2502 -3734 -2266
rect -3498 -2502 -3316 -2266
rect -3916 -2586 -3316 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 -3316 -2586
rect -3916 -2844 -3316 -2822
rect 4404 -2266 5004 5498
rect 18804 705798 19404 705820
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668454 19404 705242
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1306 19404 19898
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1884 19404 -1862
rect 22404 672054 23004 707162
rect 40404 706758 41004 707740
rect 40404 706522 40586 706758
rect 40822 706522 41004 706758
rect 40404 706438 41004 706522
rect 40404 706202 40586 706438
rect 40822 706202 41004 706438
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 4404 -2502 4586 -2266
rect 4822 -2502 5004 -2266
rect 4404 -2586 5004 -2502
rect 4404 -2822 4586 -2586
rect 4822 -2822 5004 -2586
rect -4876 -3462 -4694 -3226
rect -4458 -3462 -4276 -3226
rect -4876 -3546 -4276 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 -4276 -3546
rect -4876 -3804 -4276 -3782
rect 4404 -3804 5004 -2822
rect 22404 -3226 23004 23498
rect 36804 704838 37404 705820
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1884 37404 -902
rect 40404 690054 41004 706202
rect 58404 707718 59004 707740
rect 58404 707482 58586 707718
rect 58822 707482 59004 707718
rect 58404 707398 59004 707482
rect 58404 707162 58586 707398
rect 58822 707162 59004 707398
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 22404 -3462 22586 -3226
rect 22822 -3462 23004 -3226
rect 22404 -3546 23004 -3462
rect 22404 -3782 22586 -3546
rect 22822 -3782 23004 -3546
rect 22404 -3804 23004 -3782
rect 40404 -2266 41004 5498
rect 54804 705798 55404 705820
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668454 55404 705242
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1306 55404 19898
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1884 55404 -1862
rect 58404 672054 59004 707162
rect 76404 706758 77004 707740
rect 76404 706522 76586 706758
rect 76822 706522 77004 706758
rect 76404 706438 77004 706522
rect 76404 706202 76586 706438
rect 76822 706202 77004 706438
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 40404 -2502 40586 -2266
rect 40822 -2502 41004 -2266
rect 40404 -2586 41004 -2502
rect 40404 -2822 40586 -2586
rect 40822 -2822 41004 -2586
rect 40404 -3804 41004 -2822
rect 58404 -3226 59004 23498
rect 72804 704838 73404 705820
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1884 73404 -902
rect 76404 690054 77004 706202
rect 94404 707718 95004 707740
rect 94404 707482 94586 707718
rect 94822 707482 95004 707718
rect 94404 707398 95004 707482
rect 94404 707162 94586 707398
rect 94822 707162 95004 707398
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 58404 -3462 58586 -3226
rect 58822 -3462 59004 -3226
rect 58404 -3546 59004 -3462
rect 58404 -3782 58586 -3546
rect 58822 -3782 59004 -3546
rect 58404 -3804 59004 -3782
rect 76404 -2266 77004 5498
rect 90804 705798 91404 705820
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668454 91404 705242
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1306 91404 19898
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1884 91404 -1862
rect 94404 672054 95004 707162
rect 112404 706758 113004 707740
rect 112404 706522 112586 706758
rect 112822 706522 113004 706758
rect 112404 706438 113004 706522
rect 112404 706202 112586 706438
rect 112822 706202 113004 706438
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 76404 -2502 76586 -2266
rect 76822 -2502 77004 -2266
rect 76404 -2586 77004 -2502
rect 76404 -2822 76586 -2586
rect 76822 -2822 77004 -2586
rect 76404 -3804 77004 -2822
rect 94404 -3226 95004 23498
rect 108804 704838 109404 705820
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1884 109404 -902
rect 112404 690054 113004 706202
rect 130404 707718 131004 707740
rect 130404 707482 130586 707718
rect 130822 707482 131004 707718
rect 130404 707398 131004 707482
rect 130404 707162 130586 707398
rect 130822 707162 131004 707398
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 94404 -3462 94586 -3226
rect 94822 -3462 95004 -3226
rect 94404 -3546 95004 -3462
rect 94404 -3782 94586 -3546
rect 94822 -3782 95004 -3546
rect 94404 -3804 95004 -3782
rect 112404 -2266 113004 5498
rect 126804 705798 127404 705820
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668454 127404 705242
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1306 127404 19898
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1884 127404 -1862
rect 130404 672054 131004 707162
rect 148404 706758 149004 707740
rect 148404 706522 148586 706758
rect 148822 706522 149004 706758
rect 148404 706438 149004 706522
rect 148404 706202 148586 706438
rect 148822 706202 149004 706438
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 144804 704838 145404 705820
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 512437 145404 541898
rect 148404 690054 149004 706202
rect 166404 707718 167004 707740
rect 166404 707482 166586 707718
rect 166822 707482 167004 707718
rect 166404 707398 167004 707482
rect 166404 707162 166586 707398
rect 166822 707162 167004 707398
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 512437 149004 545498
rect 162804 705798 163404 705820
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668454 163404 705242
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 512437 163404 523898
rect 166404 672054 167004 707162
rect 184404 706758 185004 707740
rect 184404 706522 184586 706758
rect 184822 706522 185004 706758
rect 184404 706438 185004 706522
rect 184404 706202 184586 706438
rect 184822 706202 185004 706438
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 512437 167004 527498
rect 180804 704838 181404 705820
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 512437 181404 541898
rect 184404 690054 185004 706202
rect 202404 707718 203004 707740
rect 202404 707482 202586 707718
rect 202822 707482 203004 707718
rect 202404 707398 203004 707482
rect 202404 707162 202586 707398
rect 202822 707162 203004 707398
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 512437 185004 545498
rect 198804 705798 199404 705820
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668454 199404 705242
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 512437 199404 523898
rect 202404 672054 203004 707162
rect 220404 706758 221004 707740
rect 220404 706522 220586 706758
rect 220822 706522 221004 706758
rect 220404 706438 221004 706522
rect 220404 706202 220586 706438
rect 220822 706202 221004 706438
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 512437 203004 527498
rect 216804 704838 217404 705820
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 512437 217404 541898
rect 220404 690054 221004 706202
rect 238404 707718 239004 707740
rect 238404 707482 238586 707718
rect 238822 707482 239004 707718
rect 238404 707398 239004 707482
rect 238404 707162 238586 707398
rect 238822 707162 239004 707398
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 512437 221004 545498
rect 234804 705798 235404 705820
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668454 235404 705242
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 512437 235404 523898
rect 238404 672054 239004 707162
rect 256404 706758 257004 707740
rect 256404 706522 256586 706758
rect 256822 706522 257004 706758
rect 256404 706438 257004 706522
rect 256404 706202 256586 706438
rect 256822 706202 257004 706438
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 512437 239004 527498
rect 252804 704838 253404 705820
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 512437 253404 541898
rect 256404 690054 257004 706202
rect 274404 707718 275004 707740
rect 274404 707482 274586 707718
rect 274822 707482 275004 707718
rect 274404 707398 275004 707482
rect 274404 707162 274586 707398
rect 274822 707162 275004 707398
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 512437 257004 545498
rect 270804 705798 271404 705820
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668454 271404 705242
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 512437 271404 523898
rect 274404 672054 275004 707162
rect 292404 706758 293004 707740
rect 292404 706522 292586 706758
rect 292822 706522 293004 706758
rect 292404 706438 293004 706522
rect 292404 706202 292586 706438
rect 292822 706202 293004 706438
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 512437 275004 527498
rect 288804 704838 289404 705820
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 512437 289404 541898
rect 292404 690054 293004 706202
rect 310404 707718 311004 707740
rect 310404 707482 310586 707718
rect 310822 707482 311004 707718
rect 310404 707398 311004 707482
rect 310404 707162 310586 707398
rect 310822 707162 311004 707398
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 512437 293004 545498
rect 306804 705798 307404 705820
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668454 307404 705242
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 512437 307404 523898
rect 310404 672054 311004 707162
rect 328404 706758 329004 707740
rect 328404 706522 328586 706758
rect 328822 706522 329004 706758
rect 328404 706438 329004 706522
rect 328404 706202 328586 706438
rect 328822 706202 329004 706438
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 512437 311004 527498
rect 324804 704838 325404 705820
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 512437 325404 541898
rect 328404 690054 329004 706202
rect 346404 707718 347004 707740
rect 346404 707482 346586 707718
rect 346822 707482 347004 707718
rect 346404 707398 347004 707482
rect 346404 707162 346586 707398
rect 346822 707162 347004 707398
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 512437 329004 545498
rect 342804 705798 343404 705820
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668454 343404 705242
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 512437 343404 523898
rect 346404 672054 347004 707162
rect 364404 706758 365004 707740
rect 364404 706522 364586 706758
rect 364822 706522 365004 706758
rect 364404 706438 365004 706522
rect 364404 706202 364586 706438
rect 364822 706202 365004 706438
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 512437 347004 527498
rect 360804 704838 361404 705820
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 512437 361404 541898
rect 364404 690054 365004 706202
rect 382404 707718 383004 707740
rect 382404 707482 382586 707718
rect 382822 707482 383004 707718
rect 382404 707398 383004 707482
rect 382404 707162 382586 707398
rect 382822 707162 383004 707398
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 512437 365004 545498
rect 378804 705798 379404 705820
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668454 379404 705242
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 512437 379404 523898
rect 382404 672054 383004 707162
rect 400404 706758 401004 707740
rect 400404 706522 400586 706758
rect 400822 706522 401004 706758
rect 400404 706438 401004 706522
rect 400404 706202 400586 706438
rect 400822 706202 401004 706438
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 512437 383004 527498
rect 396804 704838 397404 705820
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 512437 397404 541898
rect 400404 690054 401004 706202
rect 418404 707718 419004 707740
rect 418404 707482 418586 707718
rect 418822 707482 419004 707718
rect 418404 707398 419004 707482
rect 418404 707162 418586 707398
rect 418822 707162 419004 707398
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 512437 401004 545498
rect 414804 705798 415404 705820
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668454 415404 705242
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 512437 415404 523898
rect 418404 672054 419004 707162
rect 436404 706758 437004 707740
rect 436404 706522 436586 706758
rect 436822 706522 437004 706758
rect 436404 706438 437004 706522
rect 436404 706202 436586 706438
rect 436822 706202 437004 706438
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 512437 419004 527498
rect 432804 704838 433404 705820
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 512437 433404 541898
rect 436404 690054 437004 706202
rect 454404 707718 455004 707740
rect 454404 707482 454586 707718
rect 454822 707482 455004 707718
rect 454404 707398 455004 707482
rect 454404 707162 454586 707398
rect 454822 707162 455004 707398
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 512437 437004 545498
rect 450804 705798 451404 705820
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668454 451404 705242
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 136208 510054 136528 510076
rect 136208 509818 136250 510054
rect 136486 509818 136528 510054
rect 136208 509734 136528 509818
rect 136208 509498 136250 509734
rect 136486 509498 136528 509734
rect 136208 509476 136528 509498
rect 136208 506454 136528 506476
rect 136208 506218 136250 506454
rect 136486 506218 136528 506454
rect 136208 506134 136528 506218
rect 136208 505898 136250 506134
rect 136486 505898 136528 506134
rect 136208 505876 136528 505898
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 151568 492054 151888 492076
rect 151568 491818 151610 492054
rect 151846 491818 151888 492054
rect 151568 491734 151888 491818
rect 151568 491498 151610 491734
rect 151846 491498 151888 491734
rect 151568 491476 151888 491498
rect 151568 488454 151888 488476
rect 151568 488218 151610 488454
rect 151846 488218 151888 488454
rect 151568 488134 151888 488218
rect 151568 487898 151610 488134
rect 151846 487898 151888 488134
rect 151568 487876 151888 487898
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 136208 474054 136528 474076
rect 136208 473818 136250 474054
rect 136486 473818 136528 474054
rect 136208 473734 136528 473818
rect 136208 473498 136250 473734
rect 136486 473498 136528 473734
rect 136208 473476 136528 473498
rect 136208 470454 136528 470476
rect 136208 470218 136250 470454
rect 136486 470218 136528 470454
rect 136208 470134 136528 470218
rect 136208 469898 136250 470134
rect 136486 469898 136528 470134
rect 136208 469876 136528 469898
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 151568 456054 151888 456076
rect 151568 455818 151610 456054
rect 151846 455818 151888 456054
rect 151568 455734 151888 455818
rect 151568 455498 151610 455734
rect 151846 455498 151888 455734
rect 151568 455476 151888 455498
rect 151568 452454 151888 452476
rect 151568 452218 151610 452454
rect 151846 452218 151888 452454
rect 151568 452134 151888 452218
rect 151568 451898 151610 452134
rect 151846 451898 151888 452134
rect 151568 451876 151888 451898
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 136208 438054 136528 438076
rect 136208 437818 136250 438054
rect 136486 437818 136528 438054
rect 136208 437734 136528 437818
rect 136208 437498 136250 437734
rect 136486 437498 136528 437734
rect 136208 437476 136528 437498
rect 136208 434454 136528 434476
rect 136208 434218 136250 434454
rect 136486 434218 136528 434454
rect 136208 434134 136528 434218
rect 136208 433898 136250 434134
rect 136486 433898 136528 434134
rect 136208 433876 136528 433898
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 151568 420054 151888 420076
rect 151568 419818 151610 420054
rect 151846 419818 151888 420054
rect 151568 419734 151888 419818
rect 151568 419498 151610 419734
rect 151846 419498 151888 419734
rect 151568 419476 151888 419498
rect 151568 416454 151888 416476
rect 151568 416218 151610 416454
rect 151846 416218 151888 416454
rect 151568 416134 151888 416218
rect 151568 415898 151610 416134
rect 151846 415898 151888 416134
rect 151568 415876 151888 415898
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 136208 402054 136528 402076
rect 136208 401818 136250 402054
rect 136486 401818 136528 402054
rect 136208 401734 136528 401818
rect 136208 401498 136250 401734
rect 136486 401498 136528 401734
rect 136208 401476 136528 401498
rect 136208 398454 136528 398476
rect 136208 398218 136250 398454
rect 136486 398218 136528 398454
rect 136208 398134 136528 398218
rect 136208 397898 136250 398134
rect 136486 397898 136528 398134
rect 136208 397876 136528 397898
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 151568 384054 151888 384076
rect 151568 383818 151610 384054
rect 151846 383818 151888 384054
rect 151568 383734 151888 383818
rect 151568 383498 151610 383734
rect 151846 383498 151888 383734
rect 151568 383476 151888 383498
rect 151568 380454 151888 380476
rect 151568 380218 151610 380454
rect 151846 380218 151888 380454
rect 151568 380134 151888 380218
rect 151568 379898 151610 380134
rect 151846 379898 151888 380134
rect 151568 379876 151888 379898
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 136208 366054 136528 366076
rect 136208 365818 136250 366054
rect 136486 365818 136528 366054
rect 136208 365734 136528 365818
rect 136208 365498 136250 365734
rect 136486 365498 136528 365734
rect 136208 365476 136528 365498
rect 136208 362454 136528 362476
rect 136208 362218 136250 362454
rect 136486 362218 136528 362454
rect 136208 362134 136528 362218
rect 136208 361898 136250 362134
rect 136486 361898 136528 362134
rect 136208 361876 136528 361898
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 151568 348054 151888 348076
rect 151568 347818 151610 348054
rect 151846 347818 151888 348054
rect 151568 347734 151888 347818
rect 151568 347498 151610 347734
rect 151846 347498 151888 347734
rect 151568 347476 151888 347498
rect 151568 344454 151888 344476
rect 151568 344218 151610 344454
rect 151846 344218 151888 344454
rect 151568 344134 151888 344218
rect 151568 343898 151610 344134
rect 151846 343898 151888 344134
rect 151568 343876 151888 343898
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 136208 330054 136528 330076
rect 136208 329818 136250 330054
rect 136486 329818 136528 330054
rect 136208 329734 136528 329818
rect 136208 329498 136250 329734
rect 136486 329498 136528 329734
rect 136208 329476 136528 329498
rect 136208 326454 136528 326476
rect 136208 326218 136250 326454
rect 136486 326218 136528 326454
rect 136208 326134 136528 326218
rect 136208 325898 136250 326134
rect 136486 325898 136528 326134
rect 136208 325876 136528 325898
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 151568 312054 151888 312076
rect 151568 311818 151610 312054
rect 151846 311818 151888 312054
rect 151568 311734 151888 311818
rect 151568 311498 151610 311734
rect 151846 311498 151888 311734
rect 151568 311476 151888 311498
rect 151568 308454 151888 308476
rect 151568 308218 151610 308454
rect 151846 308218 151888 308454
rect 151568 308134 151888 308218
rect 151568 307898 151610 308134
rect 151846 307898 151888 308134
rect 151568 307876 151888 307898
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 136208 294054 136528 294076
rect 136208 293818 136250 294054
rect 136486 293818 136528 294054
rect 136208 293734 136528 293818
rect 136208 293498 136250 293734
rect 136486 293498 136528 293734
rect 136208 293476 136528 293498
rect 136208 290454 136528 290476
rect 136208 290218 136250 290454
rect 136486 290218 136528 290454
rect 136208 290134 136528 290218
rect 136208 289898 136250 290134
rect 136486 289898 136528 290134
rect 136208 289876 136528 289898
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 151568 276054 151888 276076
rect 151568 275818 151610 276054
rect 151846 275818 151888 276054
rect 151568 275734 151888 275818
rect 151568 275498 151610 275734
rect 151846 275498 151888 275734
rect 151568 275476 151888 275498
rect 151568 272454 151888 272476
rect 151568 272218 151610 272454
rect 151846 272218 151888 272454
rect 151568 272134 151888 272218
rect 151568 271898 151610 272134
rect 151846 271898 151888 272134
rect 151568 271876 151888 271898
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 136208 258054 136528 258076
rect 136208 257818 136250 258054
rect 136486 257818 136528 258054
rect 136208 257734 136528 257818
rect 136208 257498 136250 257734
rect 136486 257498 136528 257734
rect 136208 257476 136528 257498
rect 136208 254454 136528 254476
rect 136208 254218 136250 254454
rect 136486 254218 136528 254454
rect 136208 254134 136528 254218
rect 136208 253898 136250 254134
rect 136486 253898 136528 254134
rect 136208 253876 136528 253898
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 151568 240054 151888 240076
rect 151568 239818 151610 240054
rect 151846 239818 151888 240054
rect 151568 239734 151888 239818
rect 151568 239498 151610 239734
rect 151846 239498 151888 239734
rect 151568 239476 151888 239498
rect 151568 236454 151888 236476
rect 151568 236218 151610 236454
rect 151846 236218 151888 236454
rect 151568 236134 151888 236218
rect 151568 235898 151610 236134
rect 151846 235898 151888 236134
rect 151568 235876 151888 235898
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 136208 222054 136528 222076
rect 136208 221818 136250 222054
rect 136486 221818 136528 222054
rect 136208 221734 136528 221818
rect 136208 221498 136250 221734
rect 136486 221498 136528 221734
rect 136208 221476 136528 221498
rect 136208 218454 136528 218476
rect 136208 218218 136250 218454
rect 136486 218218 136528 218454
rect 136208 218134 136528 218218
rect 136208 217898 136250 218134
rect 136486 217898 136528 218134
rect 136208 217876 136528 217898
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 151568 204054 151888 204076
rect 151568 203818 151610 204054
rect 151846 203818 151888 204054
rect 151568 203734 151888 203818
rect 151568 203498 151610 203734
rect 151846 203498 151888 203734
rect 151568 203476 151888 203498
rect 151568 200454 151888 200476
rect 151568 200218 151610 200454
rect 151846 200218 151888 200454
rect 151568 200134 151888 200218
rect 151568 199898 151610 200134
rect 151846 199898 151888 200134
rect 151568 199876 151888 199898
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 112404 -2502 112586 -2266
rect 112822 -2502 113004 -2266
rect 112404 -2586 113004 -2502
rect 112404 -2822 112586 -2586
rect 112822 -2822 113004 -2586
rect 112404 -3804 113004 -2822
rect 130404 -3226 131004 23498
rect 144804 182454 145404 192000
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1884 145404 -902
rect 148404 186054 149004 192000
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 130404 -3462 130586 -3226
rect 130822 -3462 131004 -3226
rect 130404 -3546 131004 -3462
rect 130404 -3782 130586 -3546
rect 130822 -3782 131004 -3546
rect 130404 -3804 131004 -3782
rect 148404 -2266 149004 5498
rect 162804 164454 163404 192000
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1306 163404 19898
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1884 163404 -1862
rect 166404 168054 167004 192000
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 148404 -2502 148586 -2266
rect 148822 -2502 149004 -2266
rect 148404 -2586 149004 -2502
rect 148404 -2822 148586 -2586
rect 148822 -2822 149004 -2586
rect 148404 -3804 149004 -2822
rect 166404 -3226 167004 23498
rect 180804 182454 181404 192000
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1884 181404 -902
rect 184404 186054 185004 192000
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 166404 -3462 166586 -3226
rect 166822 -3462 167004 -3226
rect 166404 -3546 167004 -3462
rect 166404 -3782 166586 -3546
rect 166822 -3782 167004 -3546
rect 166404 -3804 167004 -3782
rect 184404 -2266 185004 5498
rect 198804 164454 199404 192000
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1306 199404 19898
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1884 199404 -1862
rect 202404 168054 203004 192000
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 184404 -2502 184586 -2266
rect 184822 -2502 185004 -2266
rect 184404 -2586 185004 -2502
rect 184404 -2822 184586 -2586
rect 184822 -2822 185004 -2586
rect 184404 -3804 185004 -2822
rect 202404 -3226 203004 23498
rect 216804 182454 217404 192000
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1884 217404 -902
rect 220404 186054 221004 192000
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 202404 -3462 202586 -3226
rect 202822 -3462 203004 -3226
rect 202404 -3546 203004 -3462
rect 202404 -3782 202586 -3546
rect 202822 -3782 203004 -3546
rect 202404 -3804 203004 -3782
rect 220404 -2266 221004 5498
rect 234804 164454 235404 192000
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1306 235404 19898
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1884 235404 -1862
rect 238404 168054 239004 192000
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 220404 -2502 220586 -2266
rect 220822 -2502 221004 -2266
rect 220404 -2586 221004 -2502
rect 220404 -2822 220586 -2586
rect 220822 -2822 221004 -2586
rect 220404 -3804 221004 -2822
rect 238404 -3226 239004 23498
rect 252804 182454 253404 192000
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1884 253404 -902
rect 256404 186054 257004 192000
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 238404 -3462 238586 -3226
rect 238822 -3462 239004 -3226
rect 238404 -3546 239004 -3462
rect 238404 -3782 238586 -3546
rect 238822 -3782 239004 -3546
rect 238404 -3804 239004 -3782
rect 256404 -2266 257004 5498
rect 270804 164454 271404 192000
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1306 271404 19898
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1884 271404 -1862
rect 274404 168054 275004 192000
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 256404 -2502 256586 -2266
rect 256822 -2502 257004 -2266
rect 256404 -2586 257004 -2502
rect 256404 -2822 256586 -2586
rect 256822 -2822 257004 -2586
rect 256404 -3804 257004 -2822
rect 274404 -3226 275004 23498
rect 288804 182454 289404 192000
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1884 289404 -902
rect 292404 186054 293004 192000
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 274404 -3462 274586 -3226
rect 274822 -3462 275004 -3226
rect 274404 -3546 275004 -3462
rect 274404 -3782 274586 -3546
rect 274822 -3782 275004 -3546
rect 274404 -3804 275004 -3782
rect 292404 -2266 293004 5498
rect 306804 164454 307404 192000
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1306 307404 19898
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1884 307404 -1862
rect 310404 168054 311004 192000
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 292404 -2502 292586 -2266
rect 292822 -2502 293004 -2266
rect 292404 -2586 293004 -2502
rect 292404 -2822 292586 -2586
rect 292822 -2822 293004 -2586
rect 292404 -3804 293004 -2822
rect 310404 -3226 311004 23498
rect 324804 182454 325404 192000
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1884 325404 -902
rect 328404 186054 329004 192000
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 310404 -3462 310586 -3226
rect 310822 -3462 311004 -3226
rect 310404 -3546 311004 -3462
rect 310404 -3782 310586 -3546
rect 310822 -3782 311004 -3546
rect 310404 -3804 311004 -3782
rect 328404 -2266 329004 5498
rect 342804 164454 343404 192000
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1306 343404 19898
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1884 343404 -1862
rect 346404 168054 347004 192000
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 328404 -2502 328586 -2266
rect 328822 -2502 329004 -2266
rect 328404 -2586 329004 -2502
rect 328404 -2822 328586 -2586
rect 328822 -2822 329004 -2586
rect 328404 -3804 329004 -2822
rect 346404 -3226 347004 23498
rect 360804 182454 361404 192000
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1884 361404 -902
rect 364404 186054 365004 192000
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 346404 -3462 346586 -3226
rect 346822 -3462 347004 -3226
rect 346404 -3546 347004 -3462
rect 346404 -3782 346586 -3546
rect 346822 -3782 347004 -3546
rect 346404 -3804 347004 -3782
rect 364404 -2266 365004 5498
rect 378804 164454 379404 192000
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1306 379404 19898
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1884 379404 -1862
rect 382404 168054 383004 192000
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 364404 -2502 364586 -2266
rect 364822 -2502 365004 -2266
rect 364404 -2586 365004 -2502
rect 364404 -2822 364586 -2586
rect 364822 -2822 365004 -2586
rect 364404 -3804 365004 -2822
rect 382404 -3226 383004 23498
rect 396804 182454 397404 192000
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1884 397404 -902
rect 400404 186054 401004 192000
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 382404 -3462 382586 -3226
rect 382822 -3462 383004 -3226
rect 382404 -3546 383004 -3462
rect 382404 -3782 382586 -3546
rect 382822 -3782 383004 -3546
rect 382404 -3804 383004 -3782
rect 400404 -2266 401004 5498
rect 414804 164454 415404 192000
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1306 415404 19898
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1884 415404 -1862
rect 418404 168054 419004 192000
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 400404 -2502 400586 -2266
rect 400822 -2502 401004 -2266
rect 400404 -2586 401004 -2502
rect 400404 -2822 400586 -2586
rect 400822 -2822 401004 -2586
rect 400404 -3804 401004 -2822
rect 418404 -3226 419004 23498
rect 432804 182454 433404 192000
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1884 433404 -902
rect 436404 186054 437004 192000
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 418404 -3462 418586 -3226
rect 418822 -3462 419004 -3226
rect 418404 -3546 419004 -3462
rect 418404 -3782 418586 -3546
rect 418822 -3782 419004 -3546
rect 418404 -3804 419004 -3782
rect 436404 -2266 437004 5498
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1306 451404 19898
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1884 451404 -1862
rect 454404 672054 455004 707162
rect 472404 706758 473004 707740
rect 472404 706522 472586 706758
rect 472822 706522 473004 706758
rect 472404 706438 473004 706522
rect 472404 706202 472586 706438
rect 472822 706202 473004 706438
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 436404 -2502 436586 -2266
rect 436822 -2502 437004 -2266
rect 436404 -2586 437004 -2502
rect 436404 -2822 436586 -2586
rect 436822 -2822 437004 -2586
rect 436404 -3804 437004 -2822
rect 454404 -3226 455004 23498
rect 468804 704838 469404 705820
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1884 469404 -902
rect 472404 690054 473004 706202
rect 490404 707718 491004 707740
rect 490404 707482 490586 707718
rect 490822 707482 491004 707718
rect 490404 707398 491004 707482
rect 490404 707162 490586 707398
rect 490822 707162 491004 707398
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 454404 -3462 454586 -3226
rect 454822 -3462 455004 -3226
rect 454404 -3546 455004 -3462
rect 454404 -3782 454586 -3546
rect 454822 -3782 455004 -3546
rect 454404 -3804 455004 -3782
rect 472404 -2266 473004 5498
rect 486804 705798 487404 705820
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668454 487404 705242
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1306 487404 19898
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1884 487404 -1862
rect 490404 672054 491004 707162
rect 508404 706758 509004 707740
rect 508404 706522 508586 706758
rect 508822 706522 509004 706758
rect 508404 706438 509004 706522
rect 508404 706202 508586 706438
rect 508822 706202 509004 706438
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 472404 -2502 472586 -2266
rect 472822 -2502 473004 -2266
rect 472404 -2586 473004 -2502
rect 472404 -2822 472586 -2586
rect 472822 -2822 473004 -2586
rect 472404 -3804 473004 -2822
rect 490404 -3226 491004 23498
rect 504804 704838 505404 705820
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1884 505404 -902
rect 508404 690054 509004 706202
rect 526404 707718 527004 707740
rect 526404 707482 526586 707718
rect 526822 707482 527004 707718
rect 526404 707398 527004 707482
rect 526404 707162 526586 707398
rect 526822 707162 527004 707398
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 490404 -3462 490586 -3226
rect 490822 -3462 491004 -3226
rect 490404 -3546 491004 -3462
rect 490404 -3782 490586 -3546
rect 490822 -3782 491004 -3546
rect 490404 -3804 491004 -3782
rect 508404 -2266 509004 5498
rect 522804 705798 523404 705820
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668454 523404 705242
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1306 523404 19898
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1884 523404 -1862
rect 526404 672054 527004 707162
rect 544404 706758 545004 707740
rect 544404 706522 544586 706758
rect 544822 706522 545004 706758
rect 544404 706438 545004 706522
rect 544404 706202 544586 706438
rect 544822 706202 545004 706438
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 508404 -2502 508586 -2266
rect 508822 -2502 509004 -2266
rect 508404 -2586 509004 -2502
rect 508404 -2822 508586 -2586
rect 508822 -2822 509004 -2586
rect 508404 -3804 509004 -2822
rect 526404 -3226 527004 23498
rect 540804 704838 541404 705820
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1884 541404 -902
rect 544404 690054 545004 706202
rect 562404 707718 563004 707740
rect 562404 707482 562586 707718
rect 562822 707482 563004 707718
rect 562404 707398 563004 707482
rect 562404 707162 562586 707398
rect 562822 707162 563004 707398
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 526404 -3462 526586 -3226
rect 526822 -3462 527004 -3226
rect 526404 -3546 527004 -3462
rect 526404 -3782 526586 -3546
rect 526822 -3782 527004 -3546
rect 526404 -3804 527004 -3782
rect 544404 -2266 545004 5498
rect 558804 705798 559404 705820
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668454 559404 705242
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1306 559404 19898
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1884 559404 -1862
rect 562404 672054 563004 707162
rect 580404 706758 581004 707740
rect 588200 707718 588800 707740
rect 588200 707482 588382 707718
rect 588618 707482 588800 707718
rect 588200 707398 588800 707482
rect 588200 707162 588382 707398
rect 588618 707162 588800 707398
rect 580404 706522 580586 706758
rect 580822 706522 581004 706758
rect 580404 706438 581004 706522
rect 580404 706202 580586 706438
rect 580822 706202 581004 706438
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 544404 -2502 544586 -2266
rect 544822 -2502 545004 -2266
rect 544404 -2586 545004 -2502
rect 544404 -2822 544586 -2586
rect 544822 -2822 545004 -2586
rect 544404 -3804 545004 -2822
rect 562404 -3226 563004 23498
rect 576804 704838 577404 705820
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1884 577404 -902
rect 580404 690054 581004 706202
rect 587240 706758 587840 706780
rect 587240 706522 587422 706758
rect 587658 706522 587840 706758
rect 587240 706438 587840 706522
rect 587240 706202 587422 706438
rect 587658 706202 587840 706438
rect 586280 705798 586880 705820
rect 586280 705562 586462 705798
rect 586698 705562 586880 705798
rect 586280 705478 586880 705562
rect 586280 705242 586462 705478
rect 586698 705242 586880 705478
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 562404 -3462 562586 -3226
rect 562822 -3462 563004 -3226
rect 562404 -3546 563004 -3462
rect 562404 -3782 562586 -3546
rect 562822 -3782 563004 -3546
rect 562404 -3804 563004 -3782
rect 580404 -2266 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586280 668454 586880 705242
rect 586280 668218 586462 668454
rect 586698 668218 586880 668454
rect 586280 668134 586880 668218
rect 586280 667898 586462 668134
rect 586698 667898 586880 668134
rect 586280 632454 586880 667898
rect 586280 632218 586462 632454
rect 586698 632218 586880 632454
rect 586280 632134 586880 632218
rect 586280 631898 586462 632134
rect 586698 631898 586880 632134
rect 586280 596454 586880 631898
rect 586280 596218 586462 596454
rect 586698 596218 586880 596454
rect 586280 596134 586880 596218
rect 586280 595898 586462 596134
rect 586698 595898 586880 596134
rect 586280 560454 586880 595898
rect 586280 560218 586462 560454
rect 586698 560218 586880 560454
rect 586280 560134 586880 560218
rect 586280 559898 586462 560134
rect 586698 559898 586880 560134
rect 586280 524454 586880 559898
rect 586280 524218 586462 524454
rect 586698 524218 586880 524454
rect 586280 524134 586880 524218
rect 586280 523898 586462 524134
rect 586698 523898 586880 524134
rect 586280 488454 586880 523898
rect 586280 488218 586462 488454
rect 586698 488218 586880 488454
rect 586280 488134 586880 488218
rect 586280 487898 586462 488134
rect 586698 487898 586880 488134
rect 586280 452454 586880 487898
rect 586280 452218 586462 452454
rect 586698 452218 586880 452454
rect 586280 452134 586880 452218
rect 586280 451898 586462 452134
rect 586698 451898 586880 452134
rect 586280 416454 586880 451898
rect 586280 416218 586462 416454
rect 586698 416218 586880 416454
rect 586280 416134 586880 416218
rect 586280 415898 586462 416134
rect 586698 415898 586880 416134
rect 586280 380454 586880 415898
rect 586280 380218 586462 380454
rect 586698 380218 586880 380454
rect 586280 380134 586880 380218
rect 586280 379898 586462 380134
rect 586698 379898 586880 380134
rect 586280 344454 586880 379898
rect 586280 344218 586462 344454
rect 586698 344218 586880 344454
rect 586280 344134 586880 344218
rect 586280 343898 586462 344134
rect 586698 343898 586880 344134
rect 586280 308454 586880 343898
rect 586280 308218 586462 308454
rect 586698 308218 586880 308454
rect 586280 308134 586880 308218
rect 586280 307898 586462 308134
rect 586698 307898 586880 308134
rect 586280 272454 586880 307898
rect 586280 272218 586462 272454
rect 586698 272218 586880 272454
rect 586280 272134 586880 272218
rect 586280 271898 586462 272134
rect 586698 271898 586880 272134
rect 586280 236454 586880 271898
rect 586280 236218 586462 236454
rect 586698 236218 586880 236454
rect 586280 236134 586880 236218
rect 586280 235898 586462 236134
rect 586698 235898 586880 236134
rect 586280 200454 586880 235898
rect 586280 200218 586462 200454
rect 586698 200218 586880 200454
rect 586280 200134 586880 200218
rect 586280 199898 586462 200134
rect 586698 199898 586880 200134
rect 586280 164454 586880 199898
rect 586280 164218 586462 164454
rect 586698 164218 586880 164454
rect 586280 164134 586880 164218
rect 586280 163898 586462 164134
rect 586698 163898 586880 164134
rect 586280 128454 586880 163898
rect 586280 128218 586462 128454
rect 586698 128218 586880 128454
rect 586280 128134 586880 128218
rect 586280 127898 586462 128134
rect 586698 127898 586880 128134
rect 586280 92454 586880 127898
rect 586280 92218 586462 92454
rect 586698 92218 586880 92454
rect 586280 92134 586880 92218
rect 586280 91898 586462 92134
rect 586698 91898 586880 92134
rect 586280 56454 586880 91898
rect 586280 56218 586462 56454
rect 586698 56218 586880 56454
rect 586280 56134 586880 56218
rect 586280 55898 586462 56134
rect 586698 55898 586880 56134
rect 586280 20454 586880 55898
rect 586280 20218 586462 20454
rect 586698 20218 586880 20454
rect 586280 20134 586880 20218
rect 586280 19898 586462 20134
rect 586698 19898 586880 20134
rect 586280 -1306 586880 19898
rect 586280 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect 586280 -1626 586880 -1542
rect 586280 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect 586280 -1884 586880 -1862
rect 587240 690054 587840 706202
rect 587240 689818 587422 690054
rect 587658 689818 587840 690054
rect 587240 689734 587840 689818
rect 587240 689498 587422 689734
rect 587658 689498 587840 689734
rect 587240 654054 587840 689498
rect 587240 653818 587422 654054
rect 587658 653818 587840 654054
rect 587240 653734 587840 653818
rect 587240 653498 587422 653734
rect 587658 653498 587840 653734
rect 587240 618054 587840 653498
rect 587240 617818 587422 618054
rect 587658 617818 587840 618054
rect 587240 617734 587840 617818
rect 587240 617498 587422 617734
rect 587658 617498 587840 617734
rect 587240 582054 587840 617498
rect 587240 581818 587422 582054
rect 587658 581818 587840 582054
rect 587240 581734 587840 581818
rect 587240 581498 587422 581734
rect 587658 581498 587840 581734
rect 587240 546054 587840 581498
rect 587240 545818 587422 546054
rect 587658 545818 587840 546054
rect 587240 545734 587840 545818
rect 587240 545498 587422 545734
rect 587658 545498 587840 545734
rect 587240 510054 587840 545498
rect 587240 509818 587422 510054
rect 587658 509818 587840 510054
rect 587240 509734 587840 509818
rect 587240 509498 587422 509734
rect 587658 509498 587840 509734
rect 587240 474054 587840 509498
rect 587240 473818 587422 474054
rect 587658 473818 587840 474054
rect 587240 473734 587840 473818
rect 587240 473498 587422 473734
rect 587658 473498 587840 473734
rect 587240 438054 587840 473498
rect 587240 437818 587422 438054
rect 587658 437818 587840 438054
rect 587240 437734 587840 437818
rect 587240 437498 587422 437734
rect 587658 437498 587840 437734
rect 587240 402054 587840 437498
rect 587240 401818 587422 402054
rect 587658 401818 587840 402054
rect 587240 401734 587840 401818
rect 587240 401498 587422 401734
rect 587658 401498 587840 401734
rect 587240 366054 587840 401498
rect 587240 365818 587422 366054
rect 587658 365818 587840 366054
rect 587240 365734 587840 365818
rect 587240 365498 587422 365734
rect 587658 365498 587840 365734
rect 587240 330054 587840 365498
rect 587240 329818 587422 330054
rect 587658 329818 587840 330054
rect 587240 329734 587840 329818
rect 587240 329498 587422 329734
rect 587658 329498 587840 329734
rect 587240 294054 587840 329498
rect 587240 293818 587422 294054
rect 587658 293818 587840 294054
rect 587240 293734 587840 293818
rect 587240 293498 587422 293734
rect 587658 293498 587840 293734
rect 587240 258054 587840 293498
rect 587240 257818 587422 258054
rect 587658 257818 587840 258054
rect 587240 257734 587840 257818
rect 587240 257498 587422 257734
rect 587658 257498 587840 257734
rect 587240 222054 587840 257498
rect 587240 221818 587422 222054
rect 587658 221818 587840 222054
rect 587240 221734 587840 221818
rect 587240 221498 587422 221734
rect 587658 221498 587840 221734
rect 587240 186054 587840 221498
rect 587240 185818 587422 186054
rect 587658 185818 587840 186054
rect 587240 185734 587840 185818
rect 587240 185498 587422 185734
rect 587658 185498 587840 185734
rect 587240 150054 587840 185498
rect 587240 149818 587422 150054
rect 587658 149818 587840 150054
rect 587240 149734 587840 149818
rect 587240 149498 587422 149734
rect 587658 149498 587840 149734
rect 587240 114054 587840 149498
rect 587240 113818 587422 114054
rect 587658 113818 587840 114054
rect 587240 113734 587840 113818
rect 587240 113498 587422 113734
rect 587658 113498 587840 113734
rect 587240 78054 587840 113498
rect 587240 77818 587422 78054
rect 587658 77818 587840 78054
rect 587240 77734 587840 77818
rect 587240 77498 587422 77734
rect 587658 77498 587840 77734
rect 587240 42054 587840 77498
rect 587240 41818 587422 42054
rect 587658 41818 587840 42054
rect 587240 41734 587840 41818
rect 587240 41498 587422 41734
rect 587658 41498 587840 41734
rect 587240 6054 587840 41498
rect 587240 5818 587422 6054
rect 587658 5818 587840 6054
rect 587240 5734 587840 5818
rect 587240 5498 587422 5734
rect 587658 5498 587840 5734
rect 580404 -2502 580586 -2266
rect 580822 -2502 581004 -2266
rect 580404 -2586 581004 -2502
rect 580404 -2822 580586 -2586
rect 580822 -2822 581004 -2586
rect 580404 -3804 581004 -2822
rect 587240 -2266 587840 5498
rect 587240 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect 587240 -2586 587840 -2502
rect 587240 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect 587240 -2844 587840 -2822
rect 588200 672054 588800 707162
rect 588200 671818 588382 672054
rect 588618 671818 588800 672054
rect 588200 671734 588800 671818
rect 588200 671498 588382 671734
rect 588618 671498 588800 671734
rect 588200 636054 588800 671498
rect 588200 635818 588382 636054
rect 588618 635818 588800 636054
rect 588200 635734 588800 635818
rect 588200 635498 588382 635734
rect 588618 635498 588800 635734
rect 588200 600054 588800 635498
rect 588200 599818 588382 600054
rect 588618 599818 588800 600054
rect 588200 599734 588800 599818
rect 588200 599498 588382 599734
rect 588618 599498 588800 599734
rect 588200 564054 588800 599498
rect 588200 563818 588382 564054
rect 588618 563818 588800 564054
rect 588200 563734 588800 563818
rect 588200 563498 588382 563734
rect 588618 563498 588800 563734
rect 588200 528054 588800 563498
rect 588200 527818 588382 528054
rect 588618 527818 588800 528054
rect 588200 527734 588800 527818
rect 588200 527498 588382 527734
rect 588618 527498 588800 527734
rect 588200 492054 588800 527498
rect 588200 491818 588382 492054
rect 588618 491818 588800 492054
rect 588200 491734 588800 491818
rect 588200 491498 588382 491734
rect 588618 491498 588800 491734
rect 588200 456054 588800 491498
rect 588200 455818 588382 456054
rect 588618 455818 588800 456054
rect 588200 455734 588800 455818
rect 588200 455498 588382 455734
rect 588618 455498 588800 455734
rect 588200 420054 588800 455498
rect 588200 419818 588382 420054
rect 588618 419818 588800 420054
rect 588200 419734 588800 419818
rect 588200 419498 588382 419734
rect 588618 419498 588800 419734
rect 588200 384054 588800 419498
rect 588200 383818 588382 384054
rect 588618 383818 588800 384054
rect 588200 383734 588800 383818
rect 588200 383498 588382 383734
rect 588618 383498 588800 383734
rect 588200 348054 588800 383498
rect 588200 347818 588382 348054
rect 588618 347818 588800 348054
rect 588200 347734 588800 347818
rect 588200 347498 588382 347734
rect 588618 347498 588800 347734
rect 588200 312054 588800 347498
rect 588200 311818 588382 312054
rect 588618 311818 588800 312054
rect 588200 311734 588800 311818
rect 588200 311498 588382 311734
rect 588618 311498 588800 311734
rect 588200 276054 588800 311498
rect 588200 275818 588382 276054
rect 588618 275818 588800 276054
rect 588200 275734 588800 275818
rect 588200 275498 588382 275734
rect 588618 275498 588800 275734
rect 588200 240054 588800 275498
rect 588200 239818 588382 240054
rect 588618 239818 588800 240054
rect 588200 239734 588800 239818
rect 588200 239498 588382 239734
rect 588618 239498 588800 239734
rect 588200 204054 588800 239498
rect 588200 203818 588382 204054
rect 588618 203818 588800 204054
rect 588200 203734 588800 203818
rect 588200 203498 588382 203734
rect 588618 203498 588800 203734
rect 588200 168054 588800 203498
rect 588200 167818 588382 168054
rect 588618 167818 588800 168054
rect 588200 167734 588800 167818
rect 588200 167498 588382 167734
rect 588618 167498 588800 167734
rect 588200 132054 588800 167498
rect 588200 131818 588382 132054
rect 588618 131818 588800 132054
rect 588200 131734 588800 131818
rect 588200 131498 588382 131734
rect 588618 131498 588800 131734
rect 588200 96054 588800 131498
rect 588200 95818 588382 96054
rect 588618 95818 588800 96054
rect 588200 95734 588800 95818
rect 588200 95498 588382 95734
rect 588618 95498 588800 95734
rect 588200 60054 588800 95498
rect 588200 59818 588382 60054
rect 588618 59818 588800 60054
rect 588200 59734 588800 59818
rect 588200 59498 588382 59734
rect 588618 59498 588800 59734
rect 588200 24054 588800 59498
rect 588200 23818 588382 24054
rect 588618 23818 588800 24054
rect 588200 23734 588800 23818
rect 588200 23498 588382 23734
rect 588618 23498 588800 23734
rect 588200 -3226 588800 23498
rect 588200 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect 588200 -3546 588800 -3462
rect 588200 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect 588200 -3804 588800 -3782
<< via4 >>
rect -4694 707482 -4458 707718
rect -4694 707162 -4458 707398
rect -4694 671818 -4458 672054
rect -4694 671498 -4458 671734
rect -4694 635818 -4458 636054
rect -4694 635498 -4458 635734
rect -4694 599818 -4458 600054
rect -4694 599498 -4458 599734
rect -4694 563818 -4458 564054
rect -4694 563498 -4458 563734
rect -4694 527818 -4458 528054
rect -4694 527498 -4458 527734
rect -4694 491818 -4458 492054
rect -4694 491498 -4458 491734
rect -4694 455818 -4458 456054
rect -4694 455498 -4458 455734
rect -4694 419818 -4458 420054
rect -4694 419498 -4458 419734
rect -4694 383818 -4458 384054
rect -4694 383498 -4458 383734
rect -4694 347818 -4458 348054
rect -4694 347498 -4458 347734
rect -4694 311818 -4458 312054
rect -4694 311498 -4458 311734
rect -4694 275818 -4458 276054
rect -4694 275498 -4458 275734
rect -4694 239818 -4458 240054
rect -4694 239498 -4458 239734
rect -4694 203818 -4458 204054
rect -4694 203498 -4458 203734
rect -4694 167818 -4458 168054
rect -4694 167498 -4458 167734
rect -4694 131818 -4458 132054
rect -4694 131498 -4458 131734
rect -4694 95818 -4458 96054
rect -4694 95498 -4458 95734
rect -4694 59818 -4458 60054
rect -4694 59498 -4458 59734
rect -4694 23818 -4458 24054
rect -4694 23498 -4458 23734
rect -3734 706522 -3498 706758
rect -3734 706202 -3498 706438
rect 4586 706522 4822 706758
rect 4586 706202 4822 706438
rect -3734 689818 -3498 690054
rect -3734 689498 -3498 689734
rect -3734 653818 -3498 654054
rect -3734 653498 -3498 653734
rect -3734 617818 -3498 618054
rect -3734 617498 -3498 617734
rect -3734 581818 -3498 582054
rect -3734 581498 -3498 581734
rect -3734 545818 -3498 546054
rect -3734 545498 -3498 545734
rect -3734 509818 -3498 510054
rect -3734 509498 -3498 509734
rect -3734 473818 -3498 474054
rect -3734 473498 -3498 473734
rect -3734 437818 -3498 438054
rect -3734 437498 -3498 437734
rect -3734 401818 -3498 402054
rect -3734 401498 -3498 401734
rect -3734 365818 -3498 366054
rect -3734 365498 -3498 365734
rect -3734 329818 -3498 330054
rect -3734 329498 -3498 329734
rect -3734 293818 -3498 294054
rect -3734 293498 -3498 293734
rect -3734 257818 -3498 258054
rect -3734 257498 -3498 257734
rect -3734 221818 -3498 222054
rect -3734 221498 -3498 221734
rect -3734 185818 -3498 186054
rect -3734 185498 -3498 185734
rect -3734 149818 -3498 150054
rect -3734 149498 -3498 149734
rect -3734 113818 -3498 114054
rect -3734 113498 -3498 113734
rect -3734 77818 -3498 78054
rect -3734 77498 -3498 77734
rect -3734 41818 -3498 42054
rect -3734 41498 -3498 41734
rect -3734 5818 -3498 6054
rect -3734 5498 -3498 5734
rect -2774 705562 -2538 705798
rect -2774 705242 -2538 705478
rect -2774 668218 -2538 668454
rect -2774 667898 -2538 668134
rect -2774 632218 -2538 632454
rect -2774 631898 -2538 632134
rect -2774 596218 -2538 596454
rect -2774 595898 -2538 596134
rect -2774 560218 -2538 560454
rect -2774 559898 -2538 560134
rect -2774 524218 -2538 524454
rect -2774 523898 -2538 524134
rect -2774 488218 -2538 488454
rect -2774 487898 -2538 488134
rect -2774 452218 -2538 452454
rect -2774 451898 -2538 452134
rect -2774 416218 -2538 416454
rect -2774 415898 -2538 416134
rect -2774 380218 -2538 380454
rect -2774 379898 -2538 380134
rect -2774 344218 -2538 344454
rect -2774 343898 -2538 344134
rect -2774 308218 -2538 308454
rect -2774 307898 -2538 308134
rect -2774 272218 -2538 272454
rect -2774 271898 -2538 272134
rect -2774 236218 -2538 236454
rect -2774 235898 -2538 236134
rect -2774 200218 -2538 200454
rect -2774 199898 -2538 200134
rect -2774 164218 -2538 164454
rect -2774 163898 -2538 164134
rect -2774 128218 -2538 128454
rect -2774 127898 -2538 128134
rect -2774 92218 -2538 92454
rect -2774 91898 -2538 92134
rect -2774 56218 -2538 56454
rect -2774 55898 -2538 56134
rect -2774 20218 -2538 20454
rect -2774 19898 -2538 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2774 -1542 -2538 -1306
rect -2774 -1862 -2538 -1626
rect 22586 707482 22822 707718
rect 22586 707162 22822 707398
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3734 -2502 -3498 -2266
rect -3734 -2822 -3498 -2586
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 40586 706522 40822 706758
rect 40586 706202 40822 706438
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 4586 -2502 4822 -2266
rect 4586 -2822 4822 -2586
rect -4694 -3462 -4458 -3226
rect -4694 -3782 -4458 -3546
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 58586 707482 58822 707718
rect 58586 707162 58822 707398
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 22586 -3462 22822 -3226
rect 22586 -3782 22822 -3546
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 76586 706522 76822 706758
rect 76586 706202 76822 706438
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 40586 -2502 40822 -2266
rect 40586 -2822 40822 -2586
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 94586 707482 94822 707718
rect 94586 707162 94822 707398
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 58586 -3462 58822 -3226
rect 58586 -3782 58822 -3546
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 112586 706522 112822 706758
rect 112586 706202 112822 706438
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 76586 -2502 76822 -2266
rect 76586 -2822 76822 -2586
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 130586 707482 130822 707718
rect 130586 707162 130822 707398
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 94586 -3462 94822 -3226
rect 94586 -3782 94822 -3546
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 148586 706522 148822 706758
rect 148586 706202 148822 706438
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 166586 707482 166822 707718
rect 166586 707162 166822 707398
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 184586 706522 184822 706758
rect 184586 706202 184822 706438
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 202586 707482 202822 707718
rect 202586 707162 202822 707398
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 220586 706522 220822 706758
rect 220586 706202 220822 706438
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 238586 707482 238822 707718
rect 238586 707162 238822 707398
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 256586 706522 256822 706758
rect 256586 706202 256822 706438
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 274586 707482 274822 707718
rect 274586 707162 274822 707398
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 292586 706522 292822 706758
rect 292586 706202 292822 706438
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 310586 707482 310822 707718
rect 310586 707162 310822 707398
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 328586 706522 328822 706758
rect 328586 706202 328822 706438
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 346586 707482 346822 707718
rect 346586 707162 346822 707398
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 364586 706522 364822 706758
rect 364586 706202 364822 706438
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 382586 707482 382822 707718
rect 382586 707162 382822 707398
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 400586 706522 400822 706758
rect 400586 706202 400822 706438
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 418586 707482 418822 707718
rect 418586 707162 418822 707398
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 436586 706522 436822 706758
rect 436586 706202 436822 706438
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 454586 707482 454822 707718
rect 454586 707162 454822 707398
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 136250 509818 136486 510054
rect 136250 509498 136486 509734
rect 136250 506218 136486 506454
rect 136250 505898 136486 506134
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 151610 491818 151846 492054
rect 151610 491498 151846 491734
rect 151610 488218 151846 488454
rect 151610 487898 151846 488134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 136250 473818 136486 474054
rect 136250 473498 136486 473734
rect 136250 470218 136486 470454
rect 136250 469898 136486 470134
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 151610 455818 151846 456054
rect 151610 455498 151846 455734
rect 151610 452218 151846 452454
rect 151610 451898 151846 452134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 136250 437818 136486 438054
rect 136250 437498 136486 437734
rect 136250 434218 136486 434454
rect 136250 433898 136486 434134
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 151610 419818 151846 420054
rect 151610 419498 151846 419734
rect 151610 416218 151846 416454
rect 151610 415898 151846 416134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 136250 401818 136486 402054
rect 136250 401498 136486 401734
rect 136250 398218 136486 398454
rect 136250 397898 136486 398134
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 151610 383818 151846 384054
rect 151610 383498 151846 383734
rect 151610 380218 151846 380454
rect 151610 379898 151846 380134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 136250 365818 136486 366054
rect 136250 365498 136486 365734
rect 136250 362218 136486 362454
rect 136250 361898 136486 362134
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 151610 347818 151846 348054
rect 151610 347498 151846 347734
rect 151610 344218 151846 344454
rect 151610 343898 151846 344134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 136250 329818 136486 330054
rect 136250 329498 136486 329734
rect 136250 326218 136486 326454
rect 136250 325898 136486 326134
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 151610 311818 151846 312054
rect 151610 311498 151846 311734
rect 151610 308218 151846 308454
rect 151610 307898 151846 308134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 136250 293818 136486 294054
rect 136250 293498 136486 293734
rect 136250 290218 136486 290454
rect 136250 289898 136486 290134
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 151610 275818 151846 276054
rect 151610 275498 151846 275734
rect 151610 272218 151846 272454
rect 151610 271898 151846 272134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 136250 257818 136486 258054
rect 136250 257498 136486 257734
rect 136250 254218 136486 254454
rect 136250 253898 136486 254134
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 151610 239818 151846 240054
rect 151610 239498 151846 239734
rect 151610 236218 151846 236454
rect 151610 235898 151846 236134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 136250 221818 136486 222054
rect 136250 221498 136486 221734
rect 136250 218218 136486 218454
rect 136250 217898 136486 218134
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 151610 203818 151846 204054
rect 151610 203498 151846 203734
rect 151610 200218 151846 200454
rect 151610 199898 151846 200134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 112586 -2502 112822 -2266
rect 112586 -2822 112822 -2586
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 130586 -3462 130822 -3226
rect 130586 -3782 130822 -3546
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 148586 -2502 148822 -2266
rect 148586 -2822 148822 -2586
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 166586 -3462 166822 -3226
rect 166586 -3782 166822 -3546
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 184586 -2502 184822 -2266
rect 184586 -2822 184822 -2586
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 202586 -3462 202822 -3226
rect 202586 -3782 202822 -3546
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 220586 -2502 220822 -2266
rect 220586 -2822 220822 -2586
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 238586 -3462 238822 -3226
rect 238586 -3782 238822 -3546
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 256586 -2502 256822 -2266
rect 256586 -2822 256822 -2586
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 274586 -3462 274822 -3226
rect 274586 -3782 274822 -3546
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 292586 -2502 292822 -2266
rect 292586 -2822 292822 -2586
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 310586 -3462 310822 -3226
rect 310586 -3782 310822 -3546
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 328586 -2502 328822 -2266
rect 328586 -2822 328822 -2586
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 346586 -3462 346822 -3226
rect 346586 -3782 346822 -3546
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 364586 -2502 364822 -2266
rect 364586 -2822 364822 -2586
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 382586 -3462 382822 -3226
rect 382586 -3782 382822 -3546
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 400586 -2502 400822 -2266
rect 400586 -2822 400822 -2586
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 418586 -3462 418822 -3226
rect 418586 -3782 418822 -3546
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 472586 706522 472822 706758
rect 472586 706202 472822 706438
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 436586 -2502 436822 -2266
rect 436586 -2822 436822 -2586
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 490586 707482 490822 707718
rect 490586 707162 490822 707398
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 454586 -3462 454822 -3226
rect 454586 -3782 454822 -3546
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 508586 706522 508822 706758
rect 508586 706202 508822 706438
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 472586 -2502 472822 -2266
rect 472586 -2822 472822 -2586
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 526586 707482 526822 707718
rect 526586 707162 526822 707398
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 490586 -3462 490822 -3226
rect 490586 -3782 490822 -3546
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 544586 706522 544822 706758
rect 544586 706202 544822 706438
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 508586 -2502 508822 -2266
rect 508586 -2822 508822 -2586
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 562586 707482 562822 707718
rect 562586 707162 562822 707398
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 526586 -3462 526822 -3226
rect 526586 -3782 526822 -3546
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 588382 707482 588618 707718
rect 588382 707162 588618 707398
rect 580586 706522 580822 706758
rect 580586 706202 580822 706438
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 544586 -2502 544822 -2266
rect 544586 -2822 544822 -2586
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587422 706522 587658 706758
rect 587422 706202 587658 706438
rect 586462 705562 586698 705798
rect 586462 705242 586698 705478
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 562586 -3462 562822 -3226
rect 562586 -3782 562822 -3546
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586462 668218 586698 668454
rect 586462 667898 586698 668134
rect 586462 632218 586698 632454
rect 586462 631898 586698 632134
rect 586462 596218 586698 596454
rect 586462 595898 586698 596134
rect 586462 560218 586698 560454
rect 586462 559898 586698 560134
rect 586462 524218 586698 524454
rect 586462 523898 586698 524134
rect 586462 488218 586698 488454
rect 586462 487898 586698 488134
rect 586462 452218 586698 452454
rect 586462 451898 586698 452134
rect 586462 416218 586698 416454
rect 586462 415898 586698 416134
rect 586462 380218 586698 380454
rect 586462 379898 586698 380134
rect 586462 344218 586698 344454
rect 586462 343898 586698 344134
rect 586462 308218 586698 308454
rect 586462 307898 586698 308134
rect 586462 272218 586698 272454
rect 586462 271898 586698 272134
rect 586462 236218 586698 236454
rect 586462 235898 586698 236134
rect 586462 200218 586698 200454
rect 586462 199898 586698 200134
rect 586462 164218 586698 164454
rect 586462 163898 586698 164134
rect 586462 128218 586698 128454
rect 586462 127898 586698 128134
rect 586462 92218 586698 92454
rect 586462 91898 586698 92134
rect 586462 56218 586698 56454
rect 586462 55898 586698 56134
rect 586462 20218 586698 20454
rect 586462 19898 586698 20134
rect 586462 -1542 586698 -1306
rect 586462 -1862 586698 -1626
rect 587422 689818 587658 690054
rect 587422 689498 587658 689734
rect 587422 653818 587658 654054
rect 587422 653498 587658 653734
rect 587422 617818 587658 618054
rect 587422 617498 587658 617734
rect 587422 581818 587658 582054
rect 587422 581498 587658 581734
rect 587422 545818 587658 546054
rect 587422 545498 587658 545734
rect 587422 509818 587658 510054
rect 587422 509498 587658 509734
rect 587422 473818 587658 474054
rect 587422 473498 587658 473734
rect 587422 437818 587658 438054
rect 587422 437498 587658 437734
rect 587422 401818 587658 402054
rect 587422 401498 587658 401734
rect 587422 365818 587658 366054
rect 587422 365498 587658 365734
rect 587422 329818 587658 330054
rect 587422 329498 587658 329734
rect 587422 293818 587658 294054
rect 587422 293498 587658 293734
rect 587422 257818 587658 258054
rect 587422 257498 587658 257734
rect 587422 221818 587658 222054
rect 587422 221498 587658 221734
rect 587422 185818 587658 186054
rect 587422 185498 587658 185734
rect 587422 149818 587658 150054
rect 587422 149498 587658 149734
rect 587422 113818 587658 114054
rect 587422 113498 587658 113734
rect 587422 77818 587658 78054
rect 587422 77498 587658 77734
rect 587422 41818 587658 42054
rect 587422 41498 587658 41734
rect 587422 5818 587658 6054
rect 587422 5498 587658 5734
rect 580586 -2502 580822 -2266
rect 580586 -2822 580822 -2586
rect 587422 -2502 587658 -2266
rect 587422 -2822 587658 -2586
rect 588382 671818 588618 672054
rect 588382 671498 588618 671734
rect 588382 635818 588618 636054
rect 588382 635498 588618 635734
rect 588382 599818 588618 600054
rect 588382 599498 588618 599734
rect 588382 563818 588618 564054
rect 588382 563498 588618 563734
rect 588382 527818 588618 528054
rect 588382 527498 588618 527734
rect 588382 491818 588618 492054
rect 588382 491498 588618 491734
rect 588382 455818 588618 456054
rect 588382 455498 588618 455734
rect 588382 419818 588618 420054
rect 588382 419498 588618 419734
rect 588382 383818 588618 384054
rect 588382 383498 588618 383734
rect 588382 347818 588618 348054
rect 588382 347498 588618 347734
rect 588382 311818 588618 312054
rect 588382 311498 588618 311734
rect 588382 275818 588618 276054
rect 588382 275498 588618 275734
rect 588382 239818 588618 240054
rect 588382 239498 588618 239734
rect 588382 203818 588618 204054
rect 588382 203498 588618 203734
rect 588382 167818 588618 168054
rect 588382 167498 588618 167734
rect 588382 131818 588618 132054
rect 588382 131498 588618 131734
rect 588382 95818 588618 96054
rect 588382 95498 588618 95734
rect 588382 59818 588618 60054
rect 588382 59498 588618 59734
rect 588382 23818 588618 24054
rect 588382 23498 588618 23734
rect 588382 -3462 588618 -3226
rect 588382 -3782 588618 -3546
<< metal5 >>
rect -4876 707740 -4276 707742
rect 22404 707740 23004 707742
rect 58404 707740 59004 707742
rect 94404 707740 95004 707742
rect 130404 707740 131004 707742
rect 166404 707740 167004 707742
rect 202404 707740 203004 707742
rect 238404 707740 239004 707742
rect 274404 707740 275004 707742
rect 310404 707740 311004 707742
rect 346404 707740 347004 707742
rect 382404 707740 383004 707742
rect 418404 707740 419004 707742
rect 454404 707740 455004 707742
rect 490404 707740 491004 707742
rect 526404 707740 527004 707742
rect 562404 707740 563004 707742
rect 588200 707740 588800 707742
rect -4876 707718 588800 707740
rect -4876 707482 -4694 707718
rect -4458 707482 22586 707718
rect 22822 707482 58586 707718
rect 58822 707482 94586 707718
rect 94822 707482 130586 707718
rect 130822 707482 166586 707718
rect 166822 707482 202586 707718
rect 202822 707482 238586 707718
rect 238822 707482 274586 707718
rect 274822 707482 310586 707718
rect 310822 707482 346586 707718
rect 346822 707482 382586 707718
rect 382822 707482 418586 707718
rect 418822 707482 454586 707718
rect 454822 707482 490586 707718
rect 490822 707482 526586 707718
rect 526822 707482 562586 707718
rect 562822 707482 588382 707718
rect 588618 707482 588800 707718
rect -4876 707398 588800 707482
rect -4876 707162 -4694 707398
rect -4458 707162 22586 707398
rect 22822 707162 58586 707398
rect 58822 707162 94586 707398
rect 94822 707162 130586 707398
rect 130822 707162 166586 707398
rect 166822 707162 202586 707398
rect 202822 707162 238586 707398
rect 238822 707162 274586 707398
rect 274822 707162 310586 707398
rect 310822 707162 346586 707398
rect 346822 707162 382586 707398
rect 382822 707162 418586 707398
rect 418822 707162 454586 707398
rect 454822 707162 490586 707398
rect 490822 707162 526586 707398
rect 526822 707162 562586 707398
rect 562822 707162 588382 707398
rect 588618 707162 588800 707398
rect -4876 707140 588800 707162
rect -4876 707138 -4276 707140
rect 22404 707138 23004 707140
rect 58404 707138 59004 707140
rect 94404 707138 95004 707140
rect 130404 707138 131004 707140
rect 166404 707138 167004 707140
rect 202404 707138 203004 707140
rect 238404 707138 239004 707140
rect 274404 707138 275004 707140
rect 310404 707138 311004 707140
rect 346404 707138 347004 707140
rect 382404 707138 383004 707140
rect 418404 707138 419004 707140
rect 454404 707138 455004 707140
rect 490404 707138 491004 707140
rect 526404 707138 527004 707140
rect 562404 707138 563004 707140
rect 588200 707138 588800 707140
rect -3916 706780 -3316 706782
rect 4404 706780 5004 706782
rect 40404 706780 41004 706782
rect 76404 706780 77004 706782
rect 112404 706780 113004 706782
rect 148404 706780 149004 706782
rect 184404 706780 185004 706782
rect 220404 706780 221004 706782
rect 256404 706780 257004 706782
rect 292404 706780 293004 706782
rect 328404 706780 329004 706782
rect 364404 706780 365004 706782
rect 400404 706780 401004 706782
rect 436404 706780 437004 706782
rect 472404 706780 473004 706782
rect 508404 706780 509004 706782
rect 544404 706780 545004 706782
rect 580404 706780 581004 706782
rect 587240 706780 587840 706782
rect -3916 706758 587840 706780
rect -3916 706522 -3734 706758
rect -3498 706522 4586 706758
rect 4822 706522 40586 706758
rect 40822 706522 76586 706758
rect 76822 706522 112586 706758
rect 112822 706522 148586 706758
rect 148822 706522 184586 706758
rect 184822 706522 220586 706758
rect 220822 706522 256586 706758
rect 256822 706522 292586 706758
rect 292822 706522 328586 706758
rect 328822 706522 364586 706758
rect 364822 706522 400586 706758
rect 400822 706522 436586 706758
rect 436822 706522 472586 706758
rect 472822 706522 508586 706758
rect 508822 706522 544586 706758
rect 544822 706522 580586 706758
rect 580822 706522 587422 706758
rect 587658 706522 587840 706758
rect -3916 706438 587840 706522
rect -3916 706202 -3734 706438
rect -3498 706202 4586 706438
rect 4822 706202 40586 706438
rect 40822 706202 76586 706438
rect 76822 706202 112586 706438
rect 112822 706202 148586 706438
rect 148822 706202 184586 706438
rect 184822 706202 220586 706438
rect 220822 706202 256586 706438
rect 256822 706202 292586 706438
rect 292822 706202 328586 706438
rect 328822 706202 364586 706438
rect 364822 706202 400586 706438
rect 400822 706202 436586 706438
rect 436822 706202 472586 706438
rect 472822 706202 508586 706438
rect 508822 706202 544586 706438
rect 544822 706202 580586 706438
rect 580822 706202 587422 706438
rect 587658 706202 587840 706438
rect -3916 706180 587840 706202
rect -3916 706178 -3316 706180
rect 4404 706178 5004 706180
rect 40404 706178 41004 706180
rect 76404 706178 77004 706180
rect 112404 706178 113004 706180
rect 148404 706178 149004 706180
rect 184404 706178 185004 706180
rect 220404 706178 221004 706180
rect 256404 706178 257004 706180
rect 292404 706178 293004 706180
rect 328404 706178 329004 706180
rect 364404 706178 365004 706180
rect 400404 706178 401004 706180
rect 436404 706178 437004 706180
rect 472404 706178 473004 706180
rect 508404 706178 509004 706180
rect 544404 706178 545004 706180
rect 580404 706178 581004 706180
rect 587240 706178 587840 706180
rect -2956 705820 -2356 705822
rect 18804 705820 19404 705822
rect 54804 705820 55404 705822
rect 90804 705820 91404 705822
rect 126804 705820 127404 705822
rect 162804 705820 163404 705822
rect 198804 705820 199404 705822
rect 234804 705820 235404 705822
rect 270804 705820 271404 705822
rect 306804 705820 307404 705822
rect 342804 705820 343404 705822
rect 378804 705820 379404 705822
rect 414804 705820 415404 705822
rect 450804 705820 451404 705822
rect 486804 705820 487404 705822
rect 522804 705820 523404 705822
rect 558804 705820 559404 705822
rect 586280 705820 586880 705822
rect -2956 705798 586880 705820
rect -2956 705562 -2774 705798
rect -2538 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586462 705798
rect 586698 705562 586880 705798
rect -2956 705478 586880 705562
rect -2956 705242 -2774 705478
rect -2538 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586462 705478
rect 586698 705242 586880 705478
rect -2956 705220 586880 705242
rect -2956 705218 -2356 705220
rect 18804 705218 19404 705220
rect 54804 705218 55404 705220
rect 90804 705218 91404 705220
rect 126804 705218 127404 705220
rect 162804 705218 163404 705220
rect 198804 705218 199404 705220
rect 234804 705218 235404 705220
rect 270804 705218 271404 705220
rect 306804 705218 307404 705220
rect 342804 705218 343404 705220
rect 378804 705218 379404 705220
rect 414804 705218 415404 705220
rect 450804 705218 451404 705220
rect 486804 705218 487404 705220
rect 522804 705218 523404 705220
rect 558804 705218 559404 705220
rect 586280 705218 586880 705220
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -3916 690076 -3316 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587240 690076 587840 690078
rect -4876 690054 588800 690076
rect -4876 689818 -3734 690054
rect -3498 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587422 690054
rect 587658 689818 588800 690054
rect -4876 689734 588800 689818
rect -4876 689498 -3734 689734
rect -3498 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587422 689734
rect 587658 689498 588800 689734
rect -4876 689476 588800 689498
rect -3916 689474 -3316 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587240 689474 587840 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2956 686454 586880 686476
rect -2956 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586880 686454
rect -2956 686134 586880 686218
rect -2956 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586880 686134
rect -2956 685876 586880 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -4876 672076 -4276 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588200 672076 588800 672078
rect -4876 672054 588800 672076
rect -4876 671818 -4694 672054
rect -4458 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588382 672054
rect 588618 671818 588800 672054
rect -4876 671734 588800 671818
rect -4876 671498 -4694 671734
rect -4458 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588382 671734
rect 588618 671498 588800 671734
rect -4876 671476 588800 671498
rect -4876 671474 -4276 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588200 671474 588800 671476
rect -2956 668476 -2356 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586280 668476 586880 668478
rect -2956 668454 586880 668476
rect -2956 668218 -2774 668454
rect -2538 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586462 668454
rect 586698 668218 586880 668454
rect -2956 668134 586880 668218
rect -2956 667898 -2774 668134
rect -2538 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586462 668134
rect 586698 667898 586880 668134
rect -2956 667876 586880 667898
rect -2956 667874 -2356 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586280 667874 586880 667876
rect -3916 654076 -3316 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587240 654076 587840 654078
rect -4876 654054 588800 654076
rect -4876 653818 -3734 654054
rect -3498 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587422 654054
rect 587658 653818 588800 654054
rect -4876 653734 588800 653818
rect -4876 653498 -3734 653734
rect -3498 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587422 653734
rect 587658 653498 588800 653734
rect -4876 653476 588800 653498
rect -3916 653474 -3316 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587240 653474 587840 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2956 650454 586880 650476
rect -2956 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586880 650454
rect -2956 650134 586880 650218
rect -2956 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586880 650134
rect -2956 649876 586880 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -4876 636076 -4276 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588200 636076 588800 636078
rect -4876 636054 588800 636076
rect -4876 635818 -4694 636054
rect -4458 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588382 636054
rect 588618 635818 588800 636054
rect -4876 635734 588800 635818
rect -4876 635498 -4694 635734
rect -4458 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588382 635734
rect 588618 635498 588800 635734
rect -4876 635476 588800 635498
rect -4876 635474 -4276 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588200 635474 588800 635476
rect -2956 632476 -2356 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586280 632476 586880 632478
rect -2956 632454 586880 632476
rect -2956 632218 -2774 632454
rect -2538 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586462 632454
rect 586698 632218 586880 632454
rect -2956 632134 586880 632218
rect -2956 631898 -2774 632134
rect -2538 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586462 632134
rect 586698 631898 586880 632134
rect -2956 631876 586880 631898
rect -2956 631874 -2356 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586280 631874 586880 631876
rect -3916 618076 -3316 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587240 618076 587840 618078
rect -4876 618054 588800 618076
rect -4876 617818 -3734 618054
rect -3498 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587422 618054
rect 587658 617818 588800 618054
rect -4876 617734 588800 617818
rect -4876 617498 -3734 617734
rect -3498 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587422 617734
rect 587658 617498 588800 617734
rect -4876 617476 588800 617498
rect -3916 617474 -3316 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587240 617474 587840 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2956 614454 586880 614476
rect -2956 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586880 614454
rect -2956 614134 586880 614218
rect -2956 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586880 614134
rect -2956 613876 586880 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -4876 600076 -4276 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588200 600076 588800 600078
rect -4876 600054 588800 600076
rect -4876 599818 -4694 600054
rect -4458 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588382 600054
rect 588618 599818 588800 600054
rect -4876 599734 588800 599818
rect -4876 599498 -4694 599734
rect -4458 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588382 599734
rect 588618 599498 588800 599734
rect -4876 599476 588800 599498
rect -4876 599474 -4276 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588200 599474 588800 599476
rect -2956 596476 -2356 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586280 596476 586880 596478
rect -2956 596454 586880 596476
rect -2956 596218 -2774 596454
rect -2538 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586462 596454
rect 586698 596218 586880 596454
rect -2956 596134 586880 596218
rect -2956 595898 -2774 596134
rect -2538 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586462 596134
rect 586698 595898 586880 596134
rect -2956 595876 586880 595898
rect -2956 595874 -2356 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586280 595874 586880 595876
rect -3916 582076 -3316 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587240 582076 587840 582078
rect -4876 582054 588800 582076
rect -4876 581818 -3734 582054
rect -3498 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587422 582054
rect 587658 581818 588800 582054
rect -4876 581734 588800 581818
rect -4876 581498 -3734 581734
rect -3498 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587422 581734
rect 587658 581498 588800 581734
rect -4876 581476 588800 581498
rect -3916 581474 -3316 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587240 581474 587840 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2956 578454 586880 578476
rect -2956 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586880 578454
rect -2956 578134 586880 578218
rect -2956 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586880 578134
rect -2956 577876 586880 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -4876 564076 -4276 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588200 564076 588800 564078
rect -4876 564054 588800 564076
rect -4876 563818 -4694 564054
rect -4458 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588382 564054
rect 588618 563818 588800 564054
rect -4876 563734 588800 563818
rect -4876 563498 -4694 563734
rect -4458 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588382 563734
rect 588618 563498 588800 563734
rect -4876 563476 588800 563498
rect -4876 563474 -4276 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588200 563474 588800 563476
rect -2956 560476 -2356 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586280 560476 586880 560478
rect -2956 560454 586880 560476
rect -2956 560218 -2774 560454
rect -2538 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586462 560454
rect 586698 560218 586880 560454
rect -2956 560134 586880 560218
rect -2956 559898 -2774 560134
rect -2538 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586462 560134
rect 586698 559898 586880 560134
rect -2956 559876 586880 559898
rect -2956 559874 -2356 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586280 559874 586880 559876
rect -3916 546076 -3316 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587240 546076 587840 546078
rect -4876 546054 588800 546076
rect -4876 545818 -3734 546054
rect -3498 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587422 546054
rect 587658 545818 588800 546054
rect -4876 545734 588800 545818
rect -4876 545498 -3734 545734
rect -3498 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587422 545734
rect 587658 545498 588800 545734
rect -4876 545476 588800 545498
rect -3916 545474 -3316 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587240 545474 587840 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2956 542454 586880 542476
rect -2956 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586880 542454
rect -2956 542134 586880 542218
rect -2956 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586880 542134
rect -2956 541876 586880 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -4876 528076 -4276 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588200 528076 588800 528078
rect -4876 528054 588800 528076
rect -4876 527818 -4694 528054
rect -4458 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588382 528054
rect 588618 527818 588800 528054
rect -4876 527734 588800 527818
rect -4876 527498 -4694 527734
rect -4458 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588382 527734
rect 588618 527498 588800 527734
rect -4876 527476 588800 527498
rect -4876 527474 -4276 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588200 527474 588800 527476
rect -2956 524476 -2356 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586280 524476 586880 524478
rect -2956 524454 586880 524476
rect -2956 524218 -2774 524454
rect -2538 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586462 524454
rect 586698 524218 586880 524454
rect -2956 524134 586880 524218
rect -2956 523898 -2774 524134
rect -2538 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586462 524134
rect 586698 523898 586880 524134
rect -2956 523876 586880 523898
rect -2956 523874 -2356 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586280 523874 586880 523876
rect -3916 510076 -3316 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 136208 510076 136528 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587240 510076 587840 510078
rect -4876 510054 588800 510076
rect -4876 509818 -3734 510054
rect -3498 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 136250 510054
rect 136486 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587422 510054
rect 587658 509818 588800 510054
rect -4876 509734 588800 509818
rect -4876 509498 -3734 509734
rect -3498 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 136250 509734
rect 136486 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587422 509734
rect 587658 509498 588800 509734
rect -4876 509476 588800 509498
rect -3916 509474 -3316 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 136208 509474 136528 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587240 509474 587840 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 136208 506476 136528 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2956 506454 586880 506476
rect -2956 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 136250 506454
rect 136486 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586880 506454
rect -2956 506134 586880 506218
rect -2956 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 136250 506134
rect 136486 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586880 506134
rect -2956 505876 586880 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 136208 505874 136528 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -4876 492076 -4276 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 151568 492076 151888 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588200 492076 588800 492078
rect -4876 492054 588800 492076
rect -4876 491818 -4694 492054
rect -4458 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 151610 492054
rect 151846 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588382 492054
rect 588618 491818 588800 492054
rect -4876 491734 588800 491818
rect -4876 491498 -4694 491734
rect -4458 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 151610 491734
rect 151846 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588382 491734
rect 588618 491498 588800 491734
rect -4876 491476 588800 491498
rect -4876 491474 -4276 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 151568 491474 151888 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588200 491474 588800 491476
rect -2956 488476 -2356 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 151568 488476 151888 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586280 488476 586880 488478
rect -2956 488454 586880 488476
rect -2956 488218 -2774 488454
rect -2538 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 151610 488454
rect 151846 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586462 488454
rect 586698 488218 586880 488454
rect -2956 488134 586880 488218
rect -2956 487898 -2774 488134
rect -2538 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 151610 488134
rect 151846 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586462 488134
rect 586698 487898 586880 488134
rect -2956 487876 586880 487898
rect -2956 487874 -2356 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 151568 487874 151888 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586280 487874 586880 487876
rect -3916 474076 -3316 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 136208 474076 136528 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587240 474076 587840 474078
rect -4876 474054 588800 474076
rect -4876 473818 -3734 474054
rect -3498 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 136250 474054
rect 136486 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587422 474054
rect 587658 473818 588800 474054
rect -4876 473734 588800 473818
rect -4876 473498 -3734 473734
rect -3498 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 136250 473734
rect 136486 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587422 473734
rect 587658 473498 588800 473734
rect -4876 473476 588800 473498
rect -3916 473474 -3316 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 136208 473474 136528 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587240 473474 587840 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 136208 470476 136528 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2956 470454 586880 470476
rect -2956 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 136250 470454
rect 136486 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586880 470454
rect -2956 470134 586880 470218
rect -2956 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 136250 470134
rect 136486 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586880 470134
rect -2956 469876 586880 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 136208 469874 136528 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -4876 456076 -4276 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 151568 456076 151888 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588200 456076 588800 456078
rect -4876 456054 588800 456076
rect -4876 455818 -4694 456054
rect -4458 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 151610 456054
rect 151846 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588382 456054
rect 588618 455818 588800 456054
rect -4876 455734 588800 455818
rect -4876 455498 -4694 455734
rect -4458 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 151610 455734
rect 151846 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588382 455734
rect 588618 455498 588800 455734
rect -4876 455476 588800 455498
rect -4876 455474 -4276 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 151568 455474 151888 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588200 455474 588800 455476
rect -2956 452476 -2356 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 151568 452476 151888 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586280 452476 586880 452478
rect -2956 452454 586880 452476
rect -2956 452218 -2774 452454
rect -2538 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 151610 452454
rect 151846 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586462 452454
rect 586698 452218 586880 452454
rect -2956 452134 586880 452218
rect -2956 451898 -2774 452134
rect -2538 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 151610 452134
rect 151846 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586462 452134
rect 586698 451898 586880 452134
rect -2956 451876 586880 451898
rect -2956 451874 -2356 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 151568 451874 151888 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586280 451874 586880 451876
rect -3916 438076 -3316 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 136208 438076 136528 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587240 438076 587840 438078
rect -4876 438054 588800 438076
rect -4876 437818 -3734 438054
rect -3498 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 136250 438054
rect 136486 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587422 438054
rect 587658 437818 588800 438054
rect -4876 437734 588800 437818
rect -4876 437498 -3734 437734
rect -3498 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 136250 437734
rect 136486 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587422 437734
rect 587658 437498 588800 437734
rect -4876 437476 588800 437498
rect -3916 437474 -3316 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 136208 437474 136528 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587240 437474 587840 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 136208 434476 136528 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2956 434454 586880 434476
rect -2956 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 136250 434454
rect 136486 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586880 434454
rect -2956 434134 586880 434218
rect -2956 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 136250 434134
rect 136486 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586880 434134
rect -2956 433876 586880 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 136208 433874 136528 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -4876 420076 -4276 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 151568 420076 151888 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588200 420076 588800 420078
rect -4876 420054 588800 420076
rect -4876 419818 -4694 420054
rect -4458 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 151610 420054
rect 151846 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588382 420054
rect 588618 419818 588800 420054
rect -4876 419734 588800 419818
rect -4876 419498 -4694 419734
rect -4458 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 151610 419734
rect 151846 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588382 419734
rect 588618 419498 588800 419734
rect -4876 419476 588800 419498
rect -4876 419474 -4276 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 151568 419474 151888 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588200 419474 588800 419476
rect -2956 416476 -2356 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 151568 416476 151888 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586280 416476 586880 416478
rect -2956 416454 586880 416476
rect -2956 416218 -2774 416454
rect -2538 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 151610 416454
rect 151846 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586462 416454
rect 586698 416218 586880 416454
rect -2956 416134 586880 416218
rect -2956 415898 -2774 416134
rect -2538 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 151610 416134
rect 151846 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586462 416134
rect 586698 415898 586880 416134
rect -2956 415876 586880 415898
rect -2956 415874 -2356 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 151568 415874 151888 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586280 415874 586880 415876
rect -3916 402076 -3316 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 136208 402076 136528 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587240 402076 587840 402078
rect -4876 402054 588800 402076
rect -4876 401818 -3734 402054
rect -3498 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 136250 402054
rect 136486 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587422 402054
rect 587658 401818 588800 402054
rect -4876 401734 588800 401818
rect -4876 401498 -3734 401734
rect -3498 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 136250 401734
rect 136486 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587422 401734
rect 587658 401498 588800 401734
rect -4876 401476 588800 401498
rect -3916 401474 -3316 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 136208 401474 136528 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587240 401474 587840 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 136208 398476 136528 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2956 398454 586880 398476
rect -2956 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 136250 398454
rect 136486 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586880 398454
rect -2956 398134 586880 398218
rect -2956 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 136250 398134
rect 136486 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586880 398134
rect -2956 397876 586880 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 136208 397874 136528 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -4876 384076 -4276 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 151568 384076 151888 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588200 384076 588800 384078
rect -4876 384054 588800 384076
rect -4876 383818 -4694 384054
rect -4458 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 151610 384054
rect 151846 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588382 384054
rect 588618 383818 588800 384054
rect -4876 383734 588800 383818
rect -4876 383498 -4694 383734
rect -4458 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 151610 383734
rect 151846 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588382 383734
rect 588618 383498 588800 383734
rect -4876 383476 588800 383498
rect -4876 383474 -4276 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 151568 383474 151888 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588200 383474 588800 383476
rect -2956 380476 -2356 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 151568 380476 151888 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586280 380476 586880 380478
rect -2956 380454 586880 380476
rect -2956 380218 -2774 380454
rect -2538 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 151610 380454
rect 151846 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586462 380454
rect 586698 380218 586880 380454
rect -2956 380134 586880 380218
rect -2956 379898 -2774 380134
rect -2538 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 151610 380134
rect 151846 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586462 380134
rect 586698 379898 586880 380134
rect -2956 379876 586880 379898
rect -2956 379874 -2356 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 151568 379874 151888 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586280 379874 586880 379876
rect -3916 366076 -3316 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 136208 366076 136528 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587240 366076 587840 366078
rect -4876 366054 588800 366076
rect -4876 365818 -3734 366054
rect -3498 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 136250 366054
rect 136486 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587422 366054
rect 587658 365818 588800 366054
rect -4876 365734 588800 365818
rect -4876 365498 -3734 365734
rect -3498 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 136250 365734
rect 136486 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587422 365734
rect 587658 365498 588800 365734
rect -4876 365476 588800 365498
rect -3916 365474 -3316 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 136208 365474 136528 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587240 365474 587840 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 136208 362476 136528 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2956 362454 586880 362476
rect -2956 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 136250 362454
rect 136486 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586880 362454
rect -2956 362134 586880 362218
rect -2956 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 136250 362134
rect 136486 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586880 362134
rect -2956 361876 586880 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 136208 361874 136528 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -4876 348076 -4276 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 151568 348076 151888 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588200 348076 588800 348078
rect -4876 348054 588800 348076
rect -4876 347818 -4694 348054
rect -4458 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 151610 348054
rect 151846 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588382 348054
rect 588618 347818 588800 348054
rect -4876 347734 588800 347818
rect -4876 347498 -4694 347734
rect -4458 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 151610 347734
rect 151846 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588382 347734
rect 588618 347498 588800 347734
rect -4876 347476 588800 347498
rect -4876 347474 -4276 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 151568 347474 151888 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588200 347474 588800 347476
rect -2956 344476 -2356 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 151568 344476 151888 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586280 344476 586880 344478
rect -2956 344454 586880 344476
rect -2956 344218 -2774 344454
rect -2538 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 151610 344454
rect 151846 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586462 344454
rect 586698 344218 586880 344454
rect -2956 344134 586880 344218
rect -2956 343898 -2774 344134
rect -2538 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 151610 344134
rect 151846 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586462 344134
rect 586698 343898 586880 344134
rect -2956 343876 586880 343898
rect -2956 343874 -2356 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 151568 343874 151888 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586280 343874 586880 343876
rect -3916 330076 -3316 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 136208 330076 136528 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587240 330076 587840 330078
rect -4876 330054 588800 330076
rect -4876 329818 -3734 330054
rect -3498 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 136250 330054
rect 136486 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587422 330054
rect 587658 329818 588800 330054
rect -4876 329734 588800 329818
rect -4876 329498 -3734 329734
rect -3498 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 136250 329734
rect 136486 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587422 329734
rect 587658 329498 588800 329734
rect -4876 329476 588800 329498
rect -3916 329474 -3316 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 136208 329474 136528 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587240 329474 587840 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 136208 326476 136528 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2956 326454 586880 326476
rect -2956 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 136250 326454
rect 136486 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586880 326454
rect -2956 326134 586880 326218
rect -2956 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 136250 326134
rect 136486 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586880 326134
rect -2956 325876 586880 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 136208 325874 136528 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -4876 312076 -4276 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 151568 312076 151888 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588200 312076 588800 312078
rect -4876 312054 588800 312076
rect -4876 311818 -4694 312054
rect -4458 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 151610 312054
rect 151846 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588382 312054
rect 588618 311818 588800 312054
rect -4876 311734 588800 311818
rect -4876 311498 -4694 311734
rect -4458 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 151610 311734
rect 151846 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588382 311734
rect 588618 311498 588800 311734
rect -4876 311476 588800 311498
rect -4876 311474 -4276 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 151568 311474 151888 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588200 311474 588800 311476
rect -2956 308476 -2356 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 151568 308476 151888 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586280 308476 586880 308478
rect -2956 308454 586880 308476
rect -2956 308218 -2774 308454
rect -2538 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 151610 308454
rect 151846 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586462 308454
rect 586698 308218 586880 308454
rect -2956 308134 586880 308218
rect -2956 307898 -2774 308134
rect -2538 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 151610 308134
rect 151846 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586462 308134
rect 586698 307898 586880 308134
rect -2956 307876 586880 307898
rect -2956 307874 -2356 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 151568 307874 151888 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586280 307874 586880 307876
rect -3916 294076 -3316 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 136208 294076 136528 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587240 294076 587840 294078
rect -4876 294054 588800 294076
rect -4876 293818 -3734 294054
rect -3498 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 136250 294054
rect 136486 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587422 294054
rect 587658 293818 588800 294054
rect -4876 293734 588800 293818
rect -4876 293498 -3734 293734
rect -3498 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 136250 293734
rect 136486 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587422 293734
rect 587658 293498 588800 293734
rect -4876 293476 588800 293498
rect -3916 293474 -3316 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 136208 293474 136528 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587240 293474 587840 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 136208 290476 136528 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2956 290454 586880 290476
rect -2956 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 136250 290454
rect 136486 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586880 290454
rect -2956 290134 586880 290218
rect -2956 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 136250 290134
rect 136486 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586880 290134
rect -2956 289876 586880 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 136208 289874 136528 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -4876 276076 -4276 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 151568 276076 151888 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588200 276076 588800 276078
rect -4876 276054 588800 276076
rect -4876 275818 -4694 276054
rect -4458 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 151610 276054
rect 151846 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588382 276054
rect 588618 275818 588800 276054
rect -4876 275734 588800 275818
rect -4876 275498 -4694 275734
rect -4458 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 151610 275734
rect 151846 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588382 275734
rect 588618 275498 588800 275734
rect -4876 275476 588800 275498
rect -4876 275474 -4276 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 151568 275474 151888 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588200 275474 588800 275476
rect -2956 272476 -2356 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 151568 272476 151888 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586280 272476 586880 272478
rect -2956 272454 586880 272476
rect -2956 272218 -2774 272454
rect -2538 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 151610 272454
rect 151846 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586462 272454
rect 586698 272218 586880 272454
rect -2956 272134 586880 272218
rect -2956 271898 -2774 272134
rect -2538 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 151610 272134
rect 151846 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586462 272134
rect 586698 271898 586880 272134
rect -2956 271876 586880 271898
rect -2956 271874 -2356 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 151568 271874 151888 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586280 271874 586880 271876
rect -3916 258076 -3316 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 136208 258076 136528 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587240 258076 587840 258078
rect -4876 258054 588800 258076
rect -4876 257818 -3734 258054
rect -3498 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 136250 258054
rect 136486 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587422 258054
rect 587658 257818 588800 258054
rect -4876 257734 588800 257818
rect -4876 257498 -3734 257734
rect -3498 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 136250 257734
rect 136486 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587422 257734
rect 587658 257498 588800 257734
rect -4876 257476 588800 257498
rect -3916 257474 -3316 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 136208 257474 136528 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587240 257474 587840 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 136208 254476 136528 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2956 254454 586880 254476
rect -2956 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 136250 254454
rect 136486 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586880 254454
rect -2956 254134 586880 254218
rect -2956 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 136250 254134
rect 136486 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586880 254134
rect -2956 253876 586880 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 136208 253874 136528 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -4876 240076 -4276 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 151568 240076 151888 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588200 240076 588800 240078
rect -4876 240054 588800 240076
rect -4876 239818 -4694 240054
rect -4458 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 151610 240054
rect 151846 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588382 240054
rect 588618 239818 588800 240054
rect -4876 239734 588800 239818
rect -4876 239498 -4694 239734
rect -4458 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 151610 239734
rect 151846 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588382 239734
rect 588618 239498 588800 239734
rect -4876 239476 588800 239498
rect -4876 239474 -4276 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 151568 239474 151888 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588200 239474 588800 239476
rect -2956 236476 -2356 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 151568 236476 151888 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586280 236476 586880 236478
rect -2956 236454 586880 236476
rect -2956 236218 -2774 236454
rect -2538 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 151610 236454
rect 151846 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586462 236454
rect 586698 236218 586880 236454
rect -2956 236134 586880 236218
rect -2956 235898 -2774 236134
rect -2538 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 151610 236134
rect 151846 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586462 236134
rect 586698 235898 586880 236134
rect -2956 235876 586880 235898
rect -2956 235874 -2356 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 151568 235874 151888 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586280 235874 586880 235876
rect -3916 222076 -3316 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 136208 222076 136528 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587240 222076 587840 222078
rect -4876 222054 588800 222076
rect -4876 221818 -3734 222054
rect -3498 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 136250 222054
rect 136486 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587422 222054
rect 587658 221818 588800 222054
rect -4876 221734 588800 221818
rect -4876 221498 -3734 221734
rect -3498 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 136250 221734
rect 136486 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587422 221734
rect 587658 221498 588800 221734
rect -4876 221476 588800 221498
rect -3916 221474 -3316 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 136208 221474 136528 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587240 221474 587840 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 136208 218476 136528 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2956 218454 586880 218476
rect -2956 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 136250 218454
rect 136486 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586880 218454
rect -2956 218134 586880 218218
rect -2956 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 136250 218134
rect 136486 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586880 218134
rect -2956 217876 586880 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 136208 217874 136528 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -4876 204076 -4276 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 151568 204076 151888 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588200 204076 588800 204078
rect -4876 204054 588800 204076
rect -4876 203818 -4694 204054
rect -4458 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 151610 204054
rect 151846 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588382 204054
rect 588618 203818 588800 204054
rect -4876 203734 588800 203818
rect -4876 203498 -4694 203734
rect -4458 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 151610 203734
rect 151846 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588382 203734
rect 588618 203498 588800 203734
rect -4876 203476 588800 203498
rect -4876 203474 -4276 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 151568 203474 151888 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588200 203474 588800 203476
rect -2956 200476 -2356 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 151568 200476 151888 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586280 200476 586880 200478
rect -2956 200454 586880 200476
rect -2956 200218 -2774 200454
rect -2538 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 151610 200454
rect 151846 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586462 200454
rect 586698 200218 586880 200454
rect -2956 200134 586880 200218
rect -2956 199898 -2774 200134
rect -2538 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 151610 200134
rect 151846 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586462 200134
rect 586698 199898 586880 200134
rect -2956 199876 586880 199898
rect -2956 199874 -2356 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 151568 199874 151888 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586280 199874 586880 199876
rect -3916 186076 -3316 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587240 186076 587840 186078
rect -4876 186054 588800 186076
rect -4876 185818 -3734 186054
rect -3498 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587422 186054
rect 587658 185818 588800 186054
rect -4876 185734 588800 185818
rect -4876 185498 -3734 185734
rect -3498 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587422 185734
rect 587658 185498 588800 185734
rect -4876 185476 588800 185498
rect -3916 185474 -3316 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587240 185474 587840 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2956 182454 586880 182476
rect -2956 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586880 182454
rect -2956 182134 586880 182218
rect -2956 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586880 182134
rect -2956 181876 586880 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -4876 168076 -4276 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588200 168076 588800 168078
rect -4876 168054 588800 168076
rect -4876 167818 -4694 168054
rect -4458 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588382 168054
rect 588618 167818 588800 168054
rect -4876 167734 588800 167818
rect -4876 167498 -4694 167734
rect -4458 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588382 167734
rect 588618 167498 588800 167734
rect -4876 167476 588800 167498
rect -4876 167474 -4276 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588200 167474 588800 167476
rect -2956 164476 -2356 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586280 164476 586880 164478
rect -2956 164454 586880 164476
rect -2956 164218 -2774 164454
rect -2538 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586462 164454
rect 586698 164218 586880 164454
rect -2956 164134 586880 164218
rect -2956 163898 -2774 164134
rect -2538 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586462 164134
rect 586698 163898 586880 164134
rect -2956 163876 586880 163898
rect -2956 163874 -2356 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586280 163874 586880 163876
rect -3916 150076 -3316 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587240 150076 587840 150078
rect -4876 150054 588800 150076
rect -4876 149818 -3734 150054
rect -3498 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587422 150054
rect 587658 149818 588800 150054
rect -4876 149734 588800 149818
rect -4876 149498 -3734 149734
rect -3498 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587422 149734
rect 587658 149498 588800 149734
rect -4876 149476 588800 149498
rect -3916 149474 -3316 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587240 149474 587840 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2956 146454 586880 146476
rect -2956 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586880 146454
rect -2956 146134 586880 146218
rect -2956 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586880 146134
rect -2956 145876 586880 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -4876 132076 -4276 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588200 132076 588800 132078
rect -4876 132054 588800 132076
rect -4876 131818 -4694 132054
rect -4458 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588382 132054
rect 588618 131818 588800 132054
rect -4876 131734 588800 131818
rect -4876 131498 -4694 131734
rect -4458 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588382 131734
rect 588618 131498 588800 131734
rect -4876 131476 588800 131498
rect -4876 131474 -4276 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588200 131474 588800 131476
rect -2956 128476 -2356 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586280 128476 586880 128478
rect -2956 128454 586880 128476
rect -2956 128218 -2774 128454
rect -2538 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586462 128454
rect 586698 128218 586880 128454
rect -2956 128134 586880 128218
rect -2956 127898 -2774 128134
rect -2538 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586462 128134
rect 586698 127898 586880 128134
rect -2956 127876 586880 127898
rect -2956 127874 -2356 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586280 127874 586880 127876
rect -3916 114076 -3316 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587240 114076 587840 114078
rect -4876 114054 588800 114076
rect -4876 113818 -3734 114054
rect -3498 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587422 114054
rect 587658 113818 588800 114054
rect -4876 113734 588800 113818
rect -4876 113498 -3734 113734
rect -3498 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587422 113734
rect 587658 113498 588800 113734
rect -4876 113476 588800 113498
rect -3916 113474 -3316 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587240 113474 587840 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2956 110454 586880 110476
rect -2956 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586880 110454
rect -2956 110134 586880 110218
rect -2956 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586880 110134
rect -2956 109876 586880 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -4876 96076 -4276 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588200 96076 588800 96078
rect -4876 96054 588800 96076
rect -4876 95818 -4694 96054
rect -4458 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588382 96054
rect 588618 95818 588800 96054
rect -4876 95734 588800 95818
rect -4876 95498 -4694 95734
rect -4458 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588382 95734
rect 588618 95498 588800 95734
rect -4876 95476 588800 95498
rect -4876 95474 -4276 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588200 95474 588800 95476
rect -2956 92476 -2356 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586280 92476 586880 92478
rect -2956 92454 586880 92476
rect -2956 92218 -2774 92454
rect -2538 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586462 92454
rect 586698 92218 586880 92454
rect -2956 92134 586880 92218
rect -2956 91898 -2774 92134
rect -2538 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586462 92134
rect 586698 91898 586880 92134
rect -2956 91876 586880 91898
rect -2956 91874 -2356 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586280 91874 586880 91876
rect -3916 78076 -3316 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587240 78076 587840 78078
rect -4876 78054 588800 78076
rect -4876 77818 -3734 78054
rect -3498 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587422 78054
rect 587658 77818 588800 78054
rect -4876 77734 588800 77818
rect -4876 77498 -3734 77734
rect -3498 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587422 77734
rect 587658 77498 588800 77734
rect -4876 77476 588800 77498
rect -3916 77474 -3316 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587240 77474 587840 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2956 74454 586880 74476
rect -2956 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586880 74454
rect -2956 74134 586880 74218
rect -2956 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586880 74134
rect -2956 73876 586880 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -4876 60076 -4276 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588200 60076 588800 60078
rect -4876 60054 588800 60076
rect -4876 59818 -4694 60054
rect -4458 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588382 60054
rect 588618 59818 588800 60054
rect -4876 59734 588800 59818
rect -4876 59498 -4694 59734
rect -4458 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588382 59734
rect 588618 59498 588800 59734
rect -4876 59476 588800 59498
rect -4876 59474 -4276 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588200 59474 588800 59476
rect -2956 56476 -2356 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586280 56476 586880 56478
rect -2956 56454 586880 56476
rect -2956 56218 -2774 56454
rect -2538 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586462 56454
rect 586698 56218 586880 56454
rect -2956 56134 586880 56218
rect -2956 55898 -2774 56134
rect -2538 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586462 56134
rect 586698 55898 586880 56134
rect -2956 55876 586880 55898
rect -2956 55874 -2356 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586280 55874 586880 55876
rect -3916 42076 -3316 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587240 42076 587840 42078
rect -4876 42054 588800 42076
rect -4876 41818 -3734 42054
rect -3498 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587422 42054
rect 587658 41818 588800 42054
rect -4876 41734 588800 41818
rect -4876 41498 -3734 41734
rect -3498 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587422 41734
rect 587658 41498 588800 41734
rect -4876 41476 588800 41498
rect -3916 41474 -3316 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587240 41474 587840 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2956 38454 586880 38476
rect -2956 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586880 38454
rect -2956 38134 586880 38218
rect -2956 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586880 38134
rect -2956 37876 586880 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -4876 24076 -4276 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588200 24076 588800 24078
rect -4876 24054 588800 24076
rect -4876 23818 -4694 24054
rect -4458 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588382 24054
rect 588618 23818 588800 24054
rect -4876 23734 588800 23818
rect -4876 23498 -4694 23734
rect -4458 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588382 23734
rect 588618 23498 588800 23734
rect -4876 23476 588800 23498
rect -4876 23474 -4276 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588200 23474 588800 23476
rect -2956 20476 -2356 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586280 20476 586880 20478
rect -2956 20454 586880 20476
rect -2956 20218 -2774 20454
rect -2538 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586462 20454
rect 586698 20218 586880 20454
rect -2956 20134 586880 20218
rect -2956 19898 -2774 20134
rect -2538 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586462 20134
rect 586698 19898 586880 20134
rect -2956 19876 586880 19898
rect -2956 19874 -2356 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586280 19874 586880 19876
rect -3916 6076 -3316 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587240 6076 587840 6078
rect -4876 6054 588800 6076
rect -4876 5818 -3734 6054
rect -3498 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587422 6054
rect 587658 5818 588800 6054
rect -4876 5734 588800 5818
rect -4876 5498 -3734 5734
rect -3498 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587422 5734
rect 587658 5498 588800 5734
rect -4876 5476 588800 5498
rect -3916 5474 -3316 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587240 5474 587840 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2956 2454 586880 2476
rect -2956 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586880 2454
rect -2956 2134 586880 2218
rect -2956 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586880 2134
rect -2956 1876 586880 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2956 -1284 -2356 -1282
rect 18804 -1284 19404 -1282
rect 54804 -1284 55404 -1282
rect 90804 -1284 91404 -1282
rect 126804 -1284 127404 -1282
rect 162804 -1284 163404 -1282
rect 198804 -1284 199404 -1282
rect 234804 -1284 235404 -1282
rect 270804 -1284 271404 -1282
rect 306804 -1284 307404 -1282
rect 342804 -1284 343404 -1282
rect 378804 -1284 379404 -1282
rect 414804 -1284 415404 -1282
rect 450804 -1284 451404 -1282
rect 486804 -1284 487404 -1282
rect 522804 -1284 523404 -1282
rect 558804 -1284 559404 -1282
rect 586280 -1284 586880 -1282
rect -2956 -1306 586880 -1284
rect -2956 -1542 -2774 -1306
rect -2538 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect -2956 -1626 586880 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect -2956 -1884 586880 -1862
rect -2956 -1886 -2356 -1884
rect 18804 -1886 19404 -1884
rect 54804 -1886 55404 -1884
rect 90804 -1886 91404 -1884
rect 126804 -1886 127404 -1884
rect 162804 -1886 163404 -1884
rect 198804 -1886 199404 -1884
rect 234804 -1886 235404 -1884
rect 270804 -1886 271404 -1884
rect 306804 -1886 307404 -1884
rect 342804 -1886 343404 -1884
rect 378804 -1886 379404 -1884
rect 414804 -1886 415404 -1884
rect 450804 -1886 451404 -1884
rect 486804 -1886 487404 -1884
rect 522804 -1886 523404 -1884
rect 558804 -1886 559404 -1884
rect 586280 -1886 586880 -1884
rect -3916 -2244 -3316 -2242
rect 4404 -2244 5004 -2242
rect 40404 -2244 41004 -2242
rect 76404 -2244 77004 -2242
rect 112404 -2244 113004 -2242
rect 148404 -2244 149004 -2242
rect 184404 -2244 185004 -2242
rect 220404 -2244 221004 -2242
rect 256404 -2244 257004 -2242
rect 292404 -2244 293004 -2242
rect 328404 -2244 329004 -2242
rect 364404 -2244 365004 -2242
rect 400404 -2244 401004 -2242
rect 436404 -2244 437004 -2242
rect 472404 -2244 473004 -2242
rect 508404 -2244 509004 -2242
rect 544404 -2244 545004 -2242
rect 580404 -2244 581004 -2242
rect 587240 -2244 587840 -2242
rect -3916 -2266 587840 -2244
rect -3916 -2502 -3734 -2266
rect -3498 -2502 4586 -2266
rect 4822 -2502 40586 -2266
rect 40822 -2502 76586 -2266
rect 76822 -2502 112586 -2266
rect 112822 -2502 148586 -2266
rect 148822 -2502 184586 -2266
rect 184822 -2502 220586 -2266
rect 220822 -2502 256586 -2266
rect 256822 -2502 292586 -2266
rect 292822 -2502 328586 -2266
rect 328822 -2502 364586 -2266
rect 364822 -2502 400586 -2266
rect 400822 -2502 436586 -2266
rect 436822 -2502 472586 -2266
rect 472822 -2502 508586 -2266
rect 508822 -2502 544586 -2266
rect 544822 -2502 580586 -2266
rect 580822 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect -3916 -2586 587840 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 4586 -2586
rect 4822 -2822 40586 -2586
rect 40822 -2822 76586 -2586
rect 76822 -2822 112586 -2586
rect 112822 -2822 148586 -2586
rect 148822 -2822 184586 -2586
rect 184822 -2822 220586 -2586
rect 220822 -2822 256586 -2586
rect 256822 -2822 292586 -2586
rect 292822 -2822 328586 -2586
rect 328822 -2822 364586 -2586
rect 364822 -2822 400586 -2586
rect 400822 -2822 436586 -2586
rect 436822 -2822 472586 -2586
rect 472822 -2822 508586 -2586
rect 508822 -2822 544586 -2586
rect 544822 -2822 580586 -2586
rect 580822 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect -3916 -2844 587840 -2822
rect -3916 -2846 -3316 -2844
rect 4404 -2846 5004 -2844
rect 40404 -2846 41004 -2844
rect 76404 -2846 77004 -2844
rect 112404 -2846 113004 -2844
rect 148404 -2846 149004 -2844
rect 184404 -2846 185004 -2844
rect 220404 -2846 221004 -2844
rect 256404 -2846 257004 -2844
rect 292404 -2846 293004 -2844
rect 328404 -2846 329004 -2844
rect 364404 -2846 365004 -2844
rect 400404 -2846 401004 -2844
rect 436404 -2846 437004 -2844
rect 472404 -2846 473004 -2844
rect 508404 -2846 509004 -2844
rect 544404 -2846 545004 -2844
rect 580404 -2846 581004 -2844
rect 587240 -2846 587840 -2844
rect -4876 -3204 -4276 -3202
rect 22404 -3204 23004 -3202
rect 58404 -3204 59004 -3202
rect 94404 -3204 95004 -3202
rect 130404 -3204 131004 -3202
rect 166404 -3204 167004 -3202
rect 202404 -3204 203004 -3202
rect 238404 -3204 239004 -3202
rect 274404 -3204 275004 -3202
rect 310404 -3204 311004 -3202
rect 346404 -3204 347004 -3202
rect 382404 -3204 383004 -3202
rect 418404 -3204 419004 -3202
rect 454404 -3204 455004 -3202
rect 490404 -3204 491004 -3202
rect 526404 -3204 527004 -3202
rect 562404 -3204 563004 -3202
rect 588200 -3204 588800 -3202
rect -4876 -3226 588800 -3204
rect -4876 -3462 -4694 -3226
rect -4458 -3462 22586 -3226
rect 22822 -3462 58586 -3226
rect 58822 -3462 94586 -3226
rect 94822 -3462 130586 -3226
rect 130822 -3462 166586 -3226
rect 166822 -3462 202586 -3226
rect 202822 -3462 238586 -3226
rect 238822 -3462 274586 -3226
rect 274822 -3462 310586 -3226
rect 310822 -3462 346586 -3226
rect 346822 -3462 382586 -3226
rect 382822 -3462 418586 -3226
rect 418822 -3462 454586 -3226
rect 454822 -3462 490586 -3226
rect 490822 -3462 526586 -3226
rect 526822 -3462 562586 -3226
rect 562822 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect -4876 -3546 588800 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 22586 -3546
rect 22822 -3782 58586 -3546
rect 58822 -3782 94586 -3546
rect 94822 -3782 130586 -3546
rect 130822 -3782 166586 -3546
rect 166822 -3782 202586 -3546
rect 202822 -3782 238586 -3546
rect 238822 -3782 274586 -3546
rect 274822 -3782 310586 -3546
rect 310822 -3782 346586 -3546
rect 346822 -3782 382586 -3546
rect 382822 -3782 418586 -3546
rect 418822 -3782 454586 -3546
rect 454822 -3782 490586 -3546
rect 490822 -3782 526586 -3546
rect 526822 -3782 562586 -3546
rect 562822 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect -4876 -3804 588800 -3782
rect -4876 -3806 -4276 -3804
rect 22404 -3806 23004 -3804
rect 58404 -3806 59004 -3804
rect 94404 -3806 95004 -3804
rect 130404 -3806 131004 -3804
rect 166404 -3806 167004 -3804
rect 202404 -3806 203004 -3804
rect 238404 -3806 239004 -3804
rect 274404 -3806 275004 -3804
rect 310404 -3806 311004 -3804
rect 346404 -3806 347004 -3804
rect 382404 -3806 383004 -3804
rect 418404 -3806 419004 -3804
rect 454404 -3806 455004 -3804
rect 490404 -3806 491004 -3804
rect 526404 -3806 527004 -3804
rect 562404 -3806 563004 -3804
rect 588200 -3806 588800 -3804
use Ibtida_top_dffram_cv  mprj
timestamp 1608140683
transform 1 0 132000 0 1 192000
box 0 0 318293 320437
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2956 -1884 586880 -1284 8 vssd1
port 637 nsew default input
rlabel metal5 s -3916 -2844 587840 -2244 8 vccd2
port 638 nsew default input
rlabel metal5 s -4876 -3804 588800 -3204 8 vssd2
port 639 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
