VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.330 531.660 2521.650 531.720 ;
        RECT 2859.890 531.660 2860.210 531.720 ;
        RECT 2521.330 531.520 2860.210 531.660 ;
        RECT 2521.330 531.460 2521.650 531.520 ;
        RECT 2859.890 531.460 2860.210 531.520 ;
        RECT 2859.890 89.660 2860.210 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2859.890 89.520 2899.310 89.660 ;
        RECT 2859.890 89.460 2860.210 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2521.360 531.460 2521.620 531.720 ;
        RECT 2859.920 531.460 2860.180 531.720 ;
        RECT 2859.920 89.460 2860.180 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2521.350 537.355 2521.630 537.725 ;
        RECT 2521.420 531.750 2521.560 537.355 ;
        RECT 2521.360 531.430 2521.620 531.750 ;
        RECT 2859.920 531.430 2860.180 531.750 ;
        RECT 2859.980 89.750 2860.120 531.430 ;
        RECT 2859.920 89.430 2860.180 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2521.350 537.400 2521.630 537.680 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2506.000 537.690 2510.000 537.840 ;
        RECT 2521.325 537.690 2521.655 537.705 ;
        RECT 2506.000 537.390 2521.655 537.690 ;
        RECT 2506.000 537.240 2510.000 537.390 ;
        RECT 2521.325 537.375 2521.655 537.390 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 2429.200 2522.110 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2521.790 2429.060 2901.150 2429.200 ;
        RECT 2521.790 2429.000 2522.110 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
      LAYER via ;
        RECT 2521.820 2429.000 2522.080 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2521.820 2428.970 2522.080 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2521.880 2203.725 2522.020 2428.970 ;
        RECT 2521.810 2203.355 2522.090 2203.725 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2521.810 2203.400 2522.090 2203.680 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2506.000 2203.690 2510.000 2203.840 ;
        RECT 2521.785 2203.690 2522.115 2203.705 ;
        RECT 2506.000 2203.390 2522.115 2203.690 ;
        RECT 2506.000 2203.240 2510.000 2203.390 ;
        RECT 2521.785 2203.375 2522.115 2203.390 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2528.690 2663.800 2529.010 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2528.690 2663.660 2901.150 2663.800 ;
        RECT 2528.690 2663.600 2529.010 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2518.570 2371.740 2518.890 2371.800 ;
        RECT 2528.690 2371.740 2529.010 2371.800 ;
        RECT 2518.570 2371.600 2529.010 2371.740 ;
        RECT 2518.570 2371.540 2518.890 2371.600 ;
        RECT 2528.690 2371.540 2529.010 2371.600 ;
      LAYER via ;
        RECT 2528.720 2663.600 2528.980 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2518.600 2371.540 2518.860 2371.800 ;
        RECT 2528.720 2371.540 2528.980 2371.800 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2528.720 2663.570 2528.980 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2528.780 2371.830 2528.920 2663.570 ;
        RECT 2518.600 2371.510 2518.860 2371.830 ;
        RECT 2528.720 2371.510 2528.980 2371.830 ;
        RECT 2518.660 2370.325 2518.800 2371.510 ;
        RECT 2518.590 2369.955 2518.870 2370.325 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2518.590 2370.000 2518.870 2370.280 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2506.000 2370.290 2510.000 2370.440 ;
        RECT 2518.565 2370.290 2518.895 2370.305 ;
        RECT 2506.000 2369.990 2518.895 2370.290 ;
        RECT 2506.000 2369.840 2510.000 2369.990 ;
        RECT 2518.565 2369.975 2518.895 2369.990 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2556.290 2898.400 2556.610 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2556.290 2898.260 2901.150 2898.400 ;
        RECT 2556.290 2898.200 2556.610 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2525.010 2538.680 2525.330 2538.740 ;
        RECT 2556.290 2538.680 2556.610 2538.740 ;
        RECT 2525.010 2538.540 2556.610 2538.680 ;
        RECT 2525.010 2538.480 2525.330 2538.540 ;
        RECT 2556.290 2538.480 2556.610 2538.540 ;
      LAYER via ;
        RECT 2556.320 2898.200 2556.580 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2525.040 2538.480 2525.300 2538.740 ;
        RECT 2556.320 2538.480 2556.580 2538.740 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2556.320 2898.170 2556.580 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2556.380 2538.770 2556.520 2898.170 ;
        RECT 2525.040 2538.450 2525.300 2538.770 ;
        RECT 2556.320 2538.450 2556.580 2538.770 ;
        RECT 2525.100 2536.925 2525.240 2538.450 ;
        RECT 2525.030 2536.555 2525.310 2536.925 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2525.030 2536.600 2525.310 2536.880 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2506.000 2536.890 2510.000 2537.040 ;
        RECT 2525.005 2536.890 2525.335 2536.905 ;
        RECT 2506.000 2536.590 2525.335 2536.890 ;
        RECT 2506.000 2536.440 2510.000 2536.590 ;
        RECT 2525.005 2536.575 2525.335 2536.590 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2859.890 3133.000 2860.210 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2859.890 3132.860 2901.150 3133.000 ;
        RECT 2859.890 3132.800 2860.210 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2525.010 2704.600 2525.330 2704.660 ;
        RECT 2859.890 2704.600 2860.210 2704.660 ;
        RECT 2525.010 2704.460 2860.210 2704.600 ;
        RECT 2525.010 2704.400 2525.330 2704.460 ;
        RECT 2859.890 2704.400 2860.210 2704.460 ;
      LAYER via ;
        RECT 2859.920 3132.800 2860.180 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2525.040 2704.400 2525.300 2704.660 ;
        RECT 2859.920 2704.400 2860.180 2704.660 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2859.920 3132.770 2860.180 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2859.980 2704.690 2860.120 3132.770 ;
        RECT 2525.040 2704.370 2525.300 2704.690 ;
        RECT 2859.920 2704.370 2860.180 2704.690 ;
        RECT 2525.100 2703.525 2525.240 2704.370 ;
        RECT 2525.030 2703.155 2525.310 2703.525 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2525.030 2703.200 2525.310 2703.480 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2506.000 2703.490 2510.000 2703.640 ;
        RECT 2525.005 2703.490 2525.335 2703.505 ;
        RECT 2506.000 2703.190 2525.335 2703.490 ;
        RECT 2506.000 2703.040 2510.000 2703.190 ;
        RECT 2525.005 2703.175 2525.335 2703.190 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2680.490 3367.600 2680.810 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2680.490 3367.460 2901.150 3367.600 ;
        RECT 2680.490 3367.400 2680.810 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2525.010 2870.180 2525.330 2870.240 ;
        RECT 2680.490 2870.180 2680.810 2870.240 ;
        RECT 2525.010 2870.040 2680.810 2870.180 ;
        RECT 2525.010 2869.980 2525.330 2870.040 ;
        RECT 2680.490 2869.980 2680.810 2870.040 ;
      LAYER via ;
        RECT 2680.520 3367.400 2680.780 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2525.040 2869.980 2525.300 2870.240 ;
        RECT 2680.520 2869.980 2680.780 2870.240 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2680.520 3367.370 2680.780 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2680.580 2870.270 2680.720 3367.370 ;
        RECT 2525.040 2870.125 2525.300 2870.270 ;
        RECT 2525.030 2869.755 2525.310 2870.125 ;
        RECT 2680.520 2869.950 2680.780 2870.270 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2525.030 2869.800 2525.310 2870.080 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2506.000 2870.090 2510.000 2870.240 ;
        RECT 2525.005 2870.090 2525.335 2870.105 ;
        RECT 2506.000 2869.790 2525.335 2870.090 ;
        RECT 2506.000 2869.640 2510.000 2869.790 ;
        RECT 2525.005 2869.775 2525.335 2869.790 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3415.555 ;
      LAYER mcon ;
        RECT 2796.485 3415.385 2796.655 3415.555 ;
      LAYER met1 ;
        RECT 2794.570 3422.340 2794.890 3422.400 ;
        RECT 2798.250 3422.340 2798.570 3422.400 ;
        RECT 2794.570 3422.200 2798.570 3422.340 ;
        RECT 2794.570 3422.140 2794.890 3422.200 ;
        RECT 2798.250 3422.140 2798.570 3422.200 ;
        RECT 2794.570 3415.540 2794.890 3415.600 ;
        RECT 2796.425 3415.540 2796.715 3415.585 ;
        RECT 2794.570 3415.400 2796.715 3415.540 ;
        RECT 2794.570 3415.340 2794.890 3415.400 ;
        RECT 2796.425 3415.355 2796.715 3415.400 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2471.650 3019.440 2471.970 3019.500 ;
        RECT 2795.030 3019.440 2795.350 3019.500 ;
        RECT 2471.650 3019.300 2795.350 3019.440 ;
        RECT 2471.650 3019.240 2471.970 3019.300 ;
        RECT 2795.030 3019.240 2795.350 3019.300 ;
      LAYER via ;
        RECT 2794.600 3422.140 2794.860 3422.400 ;
        RECT 2798.280 3422.140 2798.540 3422.400 ;
        RECT 2794.600 3415.340 2794.860 3415.600 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2471.680 3019.240 2471.940 3019.500 ;
        RECT 2795.060 3019.240 2795.320 3019.500 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.430 2798.480 3517.600 ;
        RECT 2794.600 3422.110 2794.860 3422.430 ;
        RECT 2798.280 3422.110 2798.540 3422.430 ;
        RECT 2794.660 3415.630 2794.800 3422.110 ;
        RECT 2794.600 3415.310 2794.860 3415.630 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3019.530 2795.260 3056.610 ;
        RECT 2471.680 3019.210 2471.940 3019.530 ;
        RECT 2795.060 3019.210 2795.320 3019.530 ;
        RECT 2470.430 3009.410 2470.710 3010.000 ;
        RECT 2471.740 3009.410 2471.880 3019.210 ;
        RECT 2470.430 3009.270 2471.880 3009.410 ;
        RECT 2470.430 3006.000 2470.710 3009.270 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2470.270 3464.160 2470.590 3464.220 ;
        RECT 2474.410 3464.160 2474.730 3464.220 ;
        RECT 2470.270 3464.020 2474.730 3464.160 ;
        RECT 2470.270 3463.960 2470.590 3464.020 ;
        RECT 2474.410 3463.960 2474.730 3464.020 ;
        RECT 2470.270 3367.600 2470.590 3367.660 ;
        RECT 2471.190 3367.600 2471.510 3367.660 ;
        RECT 2470.270 3367.460 2471.510 3367.600 ;
        RECT 2470.270 3367.400 2470.590 3367.460 ;
        RECT 2471.190 3367.400 2471.510 3367.460 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2237.050 3019.440 2237.370 3019.500 ;
        RECT 2471.190 3019.440 2471.510 3019.500 ;
        RECT 2237.050 3019.300 2471.510 3019.440 ;
        RECT 2237.050 3019.240 2237.370 3019.300 ;
        RECT 2471.190 3019.240 2471.510 3019.300 ;
      LAYER via ;
        RECT 2470.300 3463.960 2470.560 3464.220 ;
        RECT 2474.440 3463.960 2474.700 3464.220 ;
        RECT 2470.300 3367.400 2470.560 3367.660 ;
        RECT 2471.220 3367.400 2471.480 3367.660 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2237.080 3019.240 2237.340 3019.500 ;
        RECT 2471.220 3019.240 2471.480 3019.500 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3464.250 2474.640 3517.230 ;
        RECT 2470.300 3463.930 2470.560 3464.250 ;
        RECT 2474.440 3463.930 2474.700 3464.250 ;
        RECT 2470.360 3415.370 2470.500 3463.930 ;
        RECT 2470.360 3415.230 2471.420 3415.370 ;
        RECT 2471.280 3367.690 2471.420 3415.230 ;
        RECT 2470.300 3367.370 2470.560 3367.690 ;
        RECT 2471.220 3367.370 2471.480 3367.690 ;
        RECT 2470.360 3318.810 2470.500 3367.370 ;
        RECT 2470.360 3318.670 2471.420 3318.810 ;
        RECT 2471.280 3270.790 2471.420 3318.670 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 3019.530 2471.420 3028.990 ;
        RECT 2237.080 3019.210 2237.340 3019.530 ;
        RECT 2471.220 3019.210 2471.480 3019.530 ;
        RECT 2237.140 3010.000 2237.280 3019.210 ;
        RECT 2237.140 3009.340 2237.490 3010.000 ;
        RECT 2237.210 3006.000 2237.490 3009.340 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3415.555 ;
      LAYER mcon ;
        RECT 2147.885 3415.385 2148.055 3415.555 ;
      LAYER met1 ;
        RECT 2145.970 3422.340 2146.290 3422.400 ;
        RECT 2149.190 3422.340 2149.510 3422.400 ;
        RECT 2145.970 3422.200 2149.510 3422.340 ;
        RECT 2145.970 3422.140 2146.290 3422.200 ;
        RECT 2149.190 3422.140 2149.510 3422.200 ;
        RECT 2145.970 3415.540 2146.290 3415.600 ;
        RECT 2147.825 3415.540 2148.115 3415.585 ;
        RECT 2145.970 3415.400 2148.115 3415.540 ;
        RECT 2145.970 3415.340 2146.290 3415.400 ;
        RECT 2147.825 3415.355 2148.115 3415.400 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2003.830 3019.100 2004.150 3019.160 ;
        RECT 2146.430 3019.100 2146.750 3019.160 ;
        RECT 2003.830 3018.960 2146.750 3019.100 ;
        RECT 2003.830 3018.900 2004.150 3018.960 ;
        RECT 2146.430 3018.900 2146.750 3018.960 ;
      LAYER via ;
        RECT 2146.000 3422.140 2146.260 3422.400 ;
        RECT 2149.220 3422.140 2149.480 3422.400 ;
        RECT 2146.000 3415.340 2146.260 3415.600 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2003.860 3018.900 2004.120 3019.160 ;
        RECT 2146.460 3018.900 2146.720 3019.160 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3422.430 2149.420 3517.600 ;
        RECT 2146.000 3422.110 2146.260 3422.430 ;
        RECT 2149.220 3422.110 2149.480 3422.430 ;
        RECT 2146.060 3415.630 2146.200 3422.110 ;
        RECT 2146.000 3415.310 2146.260 3415.630 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3019.190 2146.660 3056.610 ;
        RECT 2003.860 3018.870 2004.120 3019.190 ;
        RECT 2146.460 3018.870 2146.720 3019.190 ;
        RECT 2003.920 3010.000 2004.060 3018.870 ;
        RECT 2003.920 3009.340 2004.270 3010.000 ;
        RECT 2003.990 3006.000 2004.270 3009.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.670 3464.160 1821.990 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1821.670 3464.020 1825.670 3464.160 ;
        RECT 1821.670 3463.960 1821.990 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1821.670 3367.600 1821.990 3367.660 ;
        RECT 1822.590 3367.600 1822.910 3367.660 ;
        RECT 1821.670 3367.460 1822.910 3367.600 ;
        RECT 1821.670 3367.400 1821.990 3367.460 ;
        RECT 1822.590 3367.400 1822.910 3367.460 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1770.610 3018.760 1770.930 3018.820 ;
        RECT 1822.590 3018.760 1822.910 3018.820 ;
        RECT 1770.610 3018.620 1822.910 3018.760 ;
        RECT 1770.610 3018.560 1770.930 3018.620 ;
        RECT 1822.590 3018.560 1822.910 3018.620 ;
      LAYER via ;
        RECT 1821.700 3463.960 1821.960 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1821.700 3367.400 1821.960 3367.660 ;
        RECT 1822.620 3367.400 1822.880 3367.660 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1770.640 3018.560 1770.900 3018.820 ;
        RECT 1822.620 3018.560 1822.880 3018.820 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1821.700 3463.930 1821.960 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1821.760 3415.370 1821.900 3463.930 ;
        RECT 1821.760 3415.230 1822.820 3415.370 ;
        RECT 1822.680 3367.690 1822.820 3415.230 ;
        RECT 1821.700 3367.370 1821.960 3367.690 ;
        RECT 1822.620 3367.370 1822.880 3367.690 ;
        RECT 1821.760 3318.810 1821.900 3367.370 ;
        RECT 1821.760 3318.670 1822.820 3318.810 ;
        RECT 1822.680 3270.790 1822.820 3318.670 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 3018.850 1822.820 3028.990 ;
        RECT 1770.640 3018.530 1770.900 3018.850 ;
        RECT 1822.620 3018.530 1822.880 3018.850 ;
        RECT 1770.700 3010.000 1770.840 3018.530 ;
        RECT 1770.700 3009.340 1771.050 3010.000 ;
        RECT 1770.770 3006.000 1771.050 3009.340 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3022.160 1504.130 3022.220 ;
        RECT 1537.390 3022.160 1537.710 3022.220 ;
        RECT 1503.810 3022.020 1537.710 3022.160 ;
        RECT 1503.810 3021.960 1504.130 3022.020 ;
        RECT 1537.390 3021.960 1537.710 3022.020 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3021.960 1504.100 3022.220 ;
        RECT 1537.420 3021.960 1537.680 3022.220 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3022.250 1504.040 3498.270 ;
        RECT 1503.840 3021.930 1504.100 3022.250 ;
        RECT 1537.420 3021.930 1537.680 3022.250 ;
        RECT 1537.480 3010.000 1537.620 3021.930 ;
        RECT 1537.480 3009.340 1537.830 3010.000 ;
        RECT 1537.550 3006.000 1537.830 3009.340 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 704.040 2525.330 704.100 ;
        RECT 2639.090 704.040 2639.410 704.100 ;
        RECT 2525.010 703.900 2639.410 704.040 ;
        RECT 2525.010 703.840 2525.330 703.900 ;
        RECT 2639.090 703.840 2639.410 703.900 ;
        RECT 2639.090 324.260 2639.410 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2639.090 324.120 2899.310 324.260 ;
        RECT 2639.090 324.060 2639.410 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2525.040 703.840 2525.300 704.100 ;
        RECT 2639.120 703.840 2639.380 704.100 ;
        RECT 2639.120 324.060 2639.380 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2525.030 703.955 2525.310 704.325 ;
        RECT 2525.040 703.810 2525.300 703.955 ;
        RECT 2639.120 703.810 2639.380 704.130 ;
        RECT 2639.180 324.350 2639.320 703.810 ;
        RECT 2639.120 324.030 2639.380 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2525.030 704.000 2525.310 704.280 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2506.000 704.290 2510.000 704.440 ;
        RECT 2525.005 704.290 2525.335 704.305 ;
        RECT 2506.000 703.990 2525.335 704.290 ;
        RECT 2506.000 703.840 2510.000 703.990 ;
        RECT 2525.005 703.975 2525.335 703.990 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3019.100 1179.830 3019.160 ;
        RECT 1303.710 3019.100 1304.030 3019.160 ;
        RECT 1179.510 3018.960 1304.030 3019.100 ;
        RECT 1179.510 3018.900 1179.830 3018.960 ;
        RECT 1303.710 3018.900 1304.030 3018.960 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3018.900 1179.800 3019.160 ;
        RECT 1303.740 3018.900 1304.000 3019.160 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3019.190 1179.740 3498.270 ;
        RECT 1179.540 3018.870 1179.800 3019.190 ;
        RECT 1303.740 3018.870 1304.000 3019.190 ;
        RECT 1303.800 3010.000 1303.940 3018.870 ;
        RECT 1303.800 3009.340 1304.150 3010.000 ;
        RECT 1303.870 3006.000 1304.150 3009.340 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 3018.760 855.530 3018.820 ;
        RECT 1070.490 3018.760 1070.810 3018.820 ;
        RECT 855.210 3018.620 1070.810 3018.760 ;
        RECT 855.210 3018.560 855.530 3018.620 ;
        RECT 1070.490 3018.560 1070.810 3018.620 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 3018.560 855.500 3018.820 ;
        RECT 1070.520 3018.560 1070.780 3018.820 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 3018.850 855.440 3500.990 ;
        RECT 855.240 3018.530 855.500 3018.850 ;
        RECT 1070.520 3018.530 1070.780 3018.850 ;
        RECT 1070.580 3010.000 1070.720 3018.530 ;
        RECT 1070.580 3009.340 1070.930 3010.000 ;
        RECT 1070.650 3006.000 1070.930 3009.340 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 3018.760 531.230 3018.820 ;
        RECT 837.270 3018.760 837.590 3018.820 ;
        RECT 530.910 3018.620 837.590 3018.760 ;
        RECT 530.910 3018.560 531.230 3018.620 ;
        RECT 837.270 3018.560 837.590 3018.620 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 3018.560 531.200 3018.820 ;
        RECT 837.300 3018.560 837.560 3018.820 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3018.850 531.140 3498.270 ;
        RECT 530.940 3018.530 531.200 3018.850 ;
        RECT 837.300 3018.530 837.560 3018.850 ;
        RECT 837.360 3010.000 837.500 3018.530 ;
        RECT 837.360 3009.340 837.710 3010.000 ;
        RECT 837.430 3006.000 837.710 3009.340 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 3019.440 206.930 3019.500 ;
        RECT 604.050 3019.440 604.370 3019.500 ;
        RECT 206.610 3019.300 604.370 3019.440 ;
        RECT 206.610 3019.240 206.930 3019.300 ;
        RECT 604.050 3019.240 604.370 3019.300 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 3019.240 206.900 3019.500 ;
        RECT 604.080 3019.240 604.340 3019.500 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 3019.530 206.840 3501.670 ;
        RECT 206.640 3019.210 206.900 3019.530 ;
        RECT 604.080 3019.210 604.340 3019.530 ;
        RECT 604.140 3010.000 604.280 3019.210 ;
        RECT 604.140 3009.340 604.490 3010.000 ;
        RECT 604.210 3006.000 604.490 3009.340 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 3408.740 19.250 3408.800 ;
        RECT 161.990 3408.740 162.310 3408.800 ;
        RECT 18.930 3408.600 162.310 3408.740 ;
        RECT 18.930 3408.540 19.250 3408.600 ;
        RECT 161.990 3408.540 162.310 3408.600 ;
        RECT 161.990 2980.680 162.310 2980.740 ;
        RECT 393.370 2980.680 393.690 2980.740 ;
        RECT 161.990 2980.540 393.690 2980.680 ;
        RECT 161.990 2980.480 162.310 2980.540 ;
        RECT 393.370 2980.480 393.690 2980.540 ;
      LAYER via ;
        RECT 18.960 3408.540 19.220 3408.800 ;
        RECT 162.020 3408.540 162.280 3408.800 ;
        RECT 162.020 2980.480 162.280 2980.740 ;
        RECT 393.400 2980.480 393.660 2980.740 ;
      LAYER met2 ;
        RECT 18.950 3411.035 19.230 3411.405 ;
        RECT 19.020 3408.830 19.160 3411.035 ;
        RECT 18.960 3408.510 19.220 3408.830 ;
        RECT 162.020 3408.510 162.280 3408.830 ;
        RECT 162.080 2980.770 162.220 3408.510 ;
        RECT 162.020 2980.450 162.280 2980.770 ;
        RECT 393.400 2980.450 393.660 2980.770 ;
        RECT 393.460 2979.605 393.600 2980.450 ;
        RECT 393.390 2979.235 393.670 2979.605 ;
      LAYER via2 ;
        RECT 18.950 3411.080 19.230 3411.360 ;
        RECT 393.390 2979.280 393.670 2979.560 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 18.925 3411.370 19.255 3411.385 ;
        RECT -4.800 3411.070 19.255 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 18.925 3411.055 19.255 3411.070 ;
        RECT 393.365 2979.570 393.695 2979.585 ;
        RECT 410.000 2979.570 414.000 2979.720 ;
        RECT 393.365 2979.270 414.000 2979.570 ;
        RECT 393.365 2979.255 393.695 2979.270 ;
        RECT 410.000 2979.120 414.000 2979.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 44.690 3119.060 45.010 3119.120 ;
        RECT 16.170 3118.920 45.010 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 44.690 3118.860 45.010 3118.920 ;
        RECT 44.690 2801.160 45.010 2801.220 ;
        RECT 393.370 2801.160 393.690 2801.220 ;
        RECT 44.690 2801.020 393.690 2801.160 ;
        RECT 44.690 2800.960 45.010 2801.020 ;
        RECT 393.370 2800.960 393.690 2801.020 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 44.720 3118.860 44.980 3119.120 ;
        RECT 44.720 2800.960 44.980 2801.220 ;
        RECT 393.400 2800.960 393.660 2801.220 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 44.720 3118.830 44.980 3119.150 ;
        RECT 44.780 2801.250 44.920 3118.830 ;
        RECT 44.720 2800.930 44.980 2801.250 ;
        RECT 393.400 2800.930 393.660 2801.250 ;
        RECT 393.460 2800.765 393.600 2800.930 ;
        RECT 393.390 2800.395 393.670 2800.765 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
        RECT 393.390 2800.440 393.670 2800.720 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
        RECT 393.365 2800.730 393.695 2800.745 ;
        RECT 410.000 2800.730 414.000 2800.880 ;
        RECT 393.365 2800.430 414.000 2800.730 ;
        RECT 393.365 2800.415 393.695 2800.430 ;
        RECT 410.000 2800.280 414.000 2800.430 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 51.590 2836.180 51.910 2836.240 ;
        RECT 17.090 2836.040 51.910 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 51.590 2835.980 51.910 2836.040 ;
        RECT 51.590 2628.780 51.910 2628.840 ;
        RECT 393.370 2628.780 393.690 2628.840 ;
        RECT 51.590 2628.640 393.690 2628.780 ;
        RECT 51.590 2628.580 51.910 2628.640 ;
        RECT 393.370 2628.580 393.690 2628.640 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 51.620 2835.980 51.880 2836.240 ;
        RECT 51.620 2628.580 51.880 2628.840 ;
        RECT 393.400 2628.580 393.660 2628.840 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 51.620 2835.950 51.880 2836.270 ;
        RECT 51.680 2628.870 51.820 2835.950 ;
        RECT 51.620 2628.550 51.880 2628.870 ;
        RECT 393.400 2628.550 393.660 2628.870 ;
        RECT 393.460 2622.605 393.600 2628.550 ;
        RECT 393.390 2622.235 393.670 2622.605 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 393.390 2622.280 393.670 2622.560 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 393.365 2622.570 393.695 2622.585 ;
        RECT 410.000 2622.570 414.000 2622.720 ;
        RECT 393.365 2622.270 414.000 2622.570 ;
        RECT 393.365 2622.255 393.695 2622.270 ;
        RECT 410.000 2622.120 414.000 2622.270 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2449.260 17.410 2449.320 ;
        RECT 393.370 2449.260 393.690 2449.320 ;
        RECT 17.090 2449.120 393.690 2449.260 ;
        RECT 17.090 2449.060 17.410 2449.120 ;
        RECT 393.370 2449.060 393.690 2449.120 ;
      LAYER via ;
        RECT 17.120 2449.060 17.380 2449.320 ;
        RECT 393.400 2449.060 393.660 2449.320 ;
      LAYER met2 ;
        RECT 17.110 2549.475 17.390 2549.845 ;
        RECT 17.180 2449.350 17.320 2549.475 ;
        RECT 17.120 2449.030 17.380 2449.350 ;
        RECT 393.400 2449.030 393.660 2449.350 ;
        RECT 393.460 2443.765 393.600 2449.030 ;
        RECT 393.390 2443.395 393.670 2443.765 ;
      LAYER via2 ;
        RECT 17.110 2549.520 17.390 2549.800 ;
        RECT 393.390 2443.440 393.670 2443.720 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 17.085 2549.810 17.415 2549.825 ;
        RECT -4.800 2549.510 17.415 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 17.085 2549.495 17.415 2549.510 ;
        RECT 393.365 2443.730 393.695 2443.745 ;
        RECT 410.000 2443.730 414.000 2443.880 ;
        RECT 393.365 2443.430 414.000 2443.730 ;
        RECT 393.365 2443.415 393.695 2443.430 ;
        RECT 410.000 2443.280 414.000 2443.430 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 393.370 2262.940 393.690 2263.000 ;
        RECT 17.090 2262.800 393.690 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 393.370 2262.740 393.690 2262.800 ;
      LAYER via ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 393.400 2262.740 393.660 2263.000 ;
      LAYER met2 ;
        RECT 393.390 2265.235 393.670 2265.605 ;
        RECT 393.460 2263.030 393.600 2265.235 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 393.400 2262.710 393.660 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 393.390 2265.280 393.670 2265.560 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT 393.365 2265.570 393.695 2265.585 ;
        RECT 410.000 2265.570 414.000 2265.720 ;
        RECT 393.365 2265.270 414.000 2265.570 ;
        RECT 393.365 2265.255 393.695 2265.270 ;
        RECT 410.000 2265.120 414.000 2265.270 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 396.590 1980.060 396.910 1980.120 ;
        RECT 15.710 1979.920 396.910 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 396.590 1979.860 396.910 1979.920 ;
      LAYER via ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 396.620 1979.860 396.880 1980.120 ;
      LAYER met2 ;
        RECT 396.610 2086.395 396.890 2086.765 ;
        RECT 396.680 1980.150 396.820 2086.395 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 396.620 1979.830 396.880 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 396.610 2086.440 396.890 2086.720 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 396.585 2086.730 396.915 2086.745 ;
        RECT 410.000 2086.730 414.000 2086.880 ;
        RECT 396.585 2086.430 414.000 2086.730 ;
        RECT 396.585 2086.415 396.915 2086.430 ;
        RECT 410.000 2086.280 414.000 2086.430 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2523.630 558.860 2523.950 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2523.630 558.720 2899.310 558.860 ;
        RECT 2523.630 558.660 2523.950 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2523.660 558.660 2523.920 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2523.650 870.555 2523.930 870.925 ;
        RECT 2523.720 558.950 2523.860 870.555 ;
        RECT 2523.660 558.630 2523.920 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2523.650 870.600 2523.930 870.880 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2506.000 870.890 2510.000 871.040 ;
        RECT 2523.625 870.890 2523.955 870.905 ;
        RECT 2506.000 870.590 2523.955 870.890 ;
        RECT 2506.000 870.440 2510.000 870.590 ;
        RECT 2523.625 870.575 2523.955 870.590 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 397.970 1690.380 398.290 1690.440 ;
        RECT 17.090 1690.240 398.290 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 397.970 1690.180 398.290 1690.240 ;
      LAYER via ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 398.000 1690.180 398.260 1690.440 ;
      LAYER met2 ;
        RECT 397.990 1908.235 398.270 1908.605 ;
        RECT 398.060 1690.470 398.200 1908.235 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 398.000 1690.150 398.260 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 397.990 1908.280 398.270 1908.560 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 397.965 1908.570 398.295 1908.585 ;
        RECT 410.000 1908.570 414.000 1908.720 ;
        RECT 397.965 1908.270 414.000 1908.570 ;
        RECT 397.965 1908.255 398.295 1908.270 ;
        RECT 410.000 1908.120 414.000 1908.270 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 396.590 1476.520 396.910 1476.580 ;
        RECT 17.090 1476.380 396.910 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 396.590 1476.320 396.910 1476.380 ;
      LAYER via ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 396.620 1476.320 396.880 1476.580 ;
      LAYER met2 ;
        RECT 396.610 1729.395 396.890 1729.765 ;
        RECT 396.680 1476.610 396.820 1729.395 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 396.620 1476.290 396.880 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 396.610 1729.440 396.890 1729.720 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 396.585 1729.730 396.915 1729.745 ;
        RECT 410.000 1729.730 414.000 1729.880 ;
        RECT 396.585 1729.430 414.000 1729.730 ;
        RECT 396.585 1729.415 396.915 1729.430 ;
        RECT 410.000 1729.280 414.000 1729.430 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 397.510 1262.660 397.830 1262.720 ;
        RECT 17.090 1262.520 397.830 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 397.510 1262.460 397.830 1262.520 ;
      LAYER via ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 397.540 1262.460 397.800 1262.720 ;
      LAYER met2 ;
        RECT 397.530 1550.555 397.810 1550.925 ;
        RECT 397.600 1262.750 397.740 1550.555 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 397.540 1262.430 397.800 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 397.530 1550.600 397.810 1550.880 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 397.505 1550.890 397.835 1550.905 ;
        RECT 410.000 1550.890 414.000 1551.040 ;
        RECT 397.505 1550.590 414.000 1550.890 ;
        RECT 397.505 1550.575 397.835 1550.590 ;
        RECT 410.000 1550.440 414.000 1550.590 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 1366.360 51.910 1366.420 ;
        RECT 393.370 1366.360 393.690 1366.420 ;
        RECT 51.590 1366.220 393.690 1366.360 ;
        RECT 51.590 1366.160 51.910 1366.220 ;
        RECT 393.370 1366.160 393.690 1366.220 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 51.590 1041.660 51.910 1041.720 ;
        RECT 17.090 1041.520 51.910 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 51.590 1041.460 51.910 1041.520 ;
      LAYER via ;
        RECT 51.620 1366.160 51.880 1366.420 ;
        RECT 393.400 1366.160 393.660 1366.420 ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 51.620 1041.460 51.880 1041.720 ;
      LAYER met2 ;
        RECT 393.390 1372.395 393.670 1372.765 ;
        RECT 393.460 1366.450 393.600 1372.395 ;
        RECT 51.620 1366.130 51.880 1366.450 ;
        RECT 393.400 1366.130 393.660 1366.450 ;
        RECT 51.680 1041.750 51.820 1366.130 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 51.620 1041.430 51.880 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 393.390 1372.440 393.670 1372.720 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 393.365 1372.730 393.695 1372.745 ;
        RECT 410.000 1372.730 414.000 1372.880 ;
        RECT 393.365 1372.430 414.000 1372.730 ;
        RECT 393.365 1372.415 393.695 1372.430 ;
        RECT 410.000 1372.280 414.000 1372.430 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 1193.980 127.810 1194.040 ;
        RECT 393.370 1193.980 393.690 1194.040 ;
        RECT 127.490 1193.840 393.690 1193.980 ;
        RECT 127.490 1193.780 127.810 1193.840 ;
        RECT 393.370 1193.780 393.690 1193.840 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 127.490 827.800 127.810 827.860 ;
        RECT 17.550 827.660 127.810 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 127.490 827.600 127.810 827.660 ;
      LAYER via ;
        RECT 127.520 1193.780 127.780 1194.040 ;
        RECT 393.400 1193.780 393.660 1194.040 ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 127.520 827.600 127.780 827.860 ;
      LAYER met2 ;
        RECT 127.520 1193.750 127.780 1194.070 ;
        RECT 393.400 1193.925 393.660 1194.070 ;
        RECT 127.580 827.890 127.720 1193.750 ;
        RECT 393.390 1193.555 393.670 1193.925 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 127.520 827.570 127.780 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 393.390 1193.600 393.670 1193.880 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT 393.365 1193.890 393.695 1193.905 ;
        RECT 410.000 1193.890 414.000 1194.040 ;
        RECT 393.365 1193.590 414.000 1193.890 ;
        RECT 393.365 1193.575 393.695 1193.590 ;
        RECT 410.000 1193.440 414.000 1193.590 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 120.590 1014.460 120.910 1014.520 ;
        RECT 393.370 1014.460 393.690 1014.520 ;
        RECT 120.590 1014.320 393.690 1014.460 ;
        RECT 120.590 1014.260 120.910 1014.320 ;
        RECT 393.370 1014.260 393.690 1014.320 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 120.590 613.940 120.910 614.000 ;
        RECT 17.090 613.800 120.910 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 120.590 613.740 120.910 613.800 ;
      LAYER via ;
        RECT 120.620 1014.260 120.880 1014.520 ;
        RECT 393.400 1014.260 393.660 1014.520 ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 120.620 613.740 120.880 614.000 ;
      LAYER met2 ;
        RECT 393.390 1015.395 393.670 1015.765 ;
        RECT 393.460 1014.550 393.600 1015.395 ;
        RECT 120.620 1014.230 120.880 1014.550 ;
        RECT 393.400 1014.230 393.660 1014.550 ;
        RECT 120.680 614.030 120.820 1014.230 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 120.620 613.710 120.880 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 393.390 1015.440 393.670 1015.720 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 393.365 1015.730 393.695 1015.745 ;
        RECT 410.000 1015.730 414.000 1015.880 ;
        RECT 393.365 1015.430 414.000 1015.730 ;
        RECT 393.365 1015.415 393.695 1015.430 ;
        RECT 410.000 1015.280 414.000 1015.430 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 835.280 45.010 835.340 ;
        RECT 393.370 835.280 393.690 835.340 ;
        RECT 44.690 835.140 393.690 835.280 ;
        RECT 44.690 835.080 45.010 835.140 ;
        RECT 393.370 835.080 393.690 835.140 ;
        RECT 17.550 397.360 17.870 397.420 ;
        RECT 44.690 397.360 45.010 397.420 ;
        RECT 17.550 397.220 45.010 397.360 ;
        RECT 17.550 397.160 17.870 397.220 ;
        RECT 44.690 397.160 45.010 397.220 ;
      LAYER via ;
        RECT 44.720 835.080 44.980 835.340 ;
        RECT 393.400 835.080 393.660 835.340 ;
        RECT 17.580 397.160 17.840 397.420 ;
        RECT 44.720 397.160 44.980 397.420 ;
      LAYER met2 ;
        RECT 393.390 836.555 393.670 836.925 ;
        RECT 393.460 835.370 393.600 836.555 ;
        RECT 44.720 835.050 44.980 835.370 ;
        RECT 393.400 835.050 393.660 835.370 ;
        RECT 44.780 397.450 44.920 835.050 ;
        RECT 17.580 397.130 17.840 397.450 ;
        RECT 44.720 397.130 44.980 397.450 ;
        RECT 17.640 394.925 17.780 397.130 ;
        RECT 17.570 394.555 17.850 394.925 ;
      LAYER via2 ;
        RECT 393.390 836.600 393.670 836.880 ;
        RECT 17.570 394.600 17.850 394.880 ;
      LAYER met3 ;
        RECT 393.365 836.890 393.695 836.905 ;
        RECT 410.000 836.890 414.000 837.040 ;
        RECT 393.365 836.590 414.000 836.890 ;
        RECT 393.365 836.575 393.695 836.590 ;
        RECT 410.000 836.440 414.000 836.590 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.545 394.890 17.875 394.905 ;
        RECT -4.800 394.590 17.875 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.545 394.575 17.875 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 72.290 655.760 72.610 655.820 ;
        RECT 393.370 655.760 393.690 655.820 ;
        RECT 72.290 655.620 393.690 655.760 ;
        RECT 72.290 655.560 72.610 655.620 ;
        RECT 393.370 655.560 393.690 655.620 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 72.290 179.420 72.610 179.480 ;
        RECT 17.090 179.280 72.610 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 72.290 179.220 72.610 179.280 ;
      LAYER via ;
        RECT 72.320 655.560 72.580 655.820 ;
        RECT 393.400 655.560 393.660 655.820 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 72.320 179.220 72.580 179.480 ;
      LAYER met2 ;
        RECT 393.390 658.395 393.670 658.765 ;
        RECT 393.460 655.850 393.600 658.395 ;
        RECT 72.320 655.530 72.580 655.850 ;
        RECT 393.400 655.530 393.660 655.850 ;
        RECT 72.380 179.510 72.520 655.530 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 72.320 179.190 72.580 179.510 ;
      LAYER via2 ;
        RECT 393.390 658.440 393.670 658.720 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 393.365 658.730 393.695 658.745 ;
        RECT 410.000 658.730 414.000 658.880 ;
        RECT 393.365 658.430 414.000 658.730 ;
        RECT 393.365 658.415 393.695 658.430 ;
        RECT 410.000 658.280 414.000 658.430 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.250 793.460 2522.570 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2522.250 793.320 2899.310 793.460 ;
        RECT 2522.250 793.260 2522.570 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2522.280 793.260 2522.540 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2522.270 1037.155 2522.550 1037.525 ;
        RECT 2522.340 793.550 2522.480 1037.155 ;
        RECT 2522.280 793.230 2522.540 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2522.270 1037.200 2522.550 1037.480 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2506.000 1037.490 2510.000 1037.640 ;
        RECT 2522.245 1037.490 2522.575 1037.505 ;
        RECT 2506.000 1037.190 2522.575 1037.490 ;
        RECT 2506.000 1037.040 2510.000 1037.190 ;
        RECT 2522.245 1037.175 2522.575 1037.190 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1028.060 2522.110 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2521.790 1027.920 2899.310 1028.060 ;
        RECT 2521.790 1027.860 2522.110 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2521.820 1027.860 2522.080 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2521.810 1203.755 2522.090 1204.125 ;
        RECT 2521.880 1028.150 2522.020 1203.755 ;
        RECT 2521.820 1027.830 2522.080 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2521.810 1203.800 2522.090 1204.080 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2506.000 1204.090 2510.000 1204.240 ;
        RECT 2521.785 1204.090 2522.115 1204.105 ;
        RECT 2506.000 1203.790 2522.115 1204.090 ;
        RECT 2506.000 1203.640 2510.000 1203.790 ;
        RECT 2521.785 1203.775 2522.115 1203.790 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1262.660 2522.110 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2521.790 1262.520 2899.310 1262.660 ;
        RECT 2521.790 1262.460 2522.110 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2521.820 1262.460 2522.080 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2521.810 1370.355 2522.090 1370.725 ;
        RECT 2521.880 1262.750 2522.020 1370.355 ;
        RECT 2521.820 1262.430 2522.080 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2521.810 1370.400 2522.090 1370.680 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2506.000 1370.690 2510.000 1370.840 ;
        RECT 2521.785 1370.690 2522.115 1370.705 ;
        RECT 2506.000 1370.390 2522.115 1370.690 ;
        RECT 2506.000 1370.240 2510.000 1370.390 ;
        RECT 2521.785 1370.375 2522.115 1370.390 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1497.260 2522.110 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 2521.790 1497.120 2899.310 1497.260 ;
        RECT 2521.790 1497.060 2522.110 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 2521.820 1497.060 2522.080 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 2521.810 1536.955 2522.090 1537.325 ;
        RECT 2521.880 1497.350 2522.020 1536.955 ;
        RECT 2521.820 1497.030 2522.080 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2521.810 1537.000 2522.090 1537.280 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2506.000 1537.290 2510.000 1537.440 ;
        RECT 2521.785 1537.290 2522.115 1537.305 ;
        RECT 2506.000 1536.990 2522.115 1537.290 ;
        RECT 2506.000 1536.840 2510.000 1536.990 ;
        RECT 2521.785 1536.975 2522.115 1536.990 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1704.320 2525.330 1704.380 ;
        RECT 2904.510 1704.320 2904.830 1704.380 ;
        RECT 2525.010 1704.180 2904.830 1704.320 ;
        RECT 2525.010 1704.120 2525.330 1704.180 ;
        RECT 2904.510 1704.120 2904.830 1704.180 ;
      LAYER via ;
        RECT 2525.040 1704.120 2525.300 1704.380 ;
        RECT 2904.540 1704.120 2904.800 1704.380 ;
      LAYER met2 ;
        RECT 2904.530 1730.075 2904.810 1730.445 ;
        RECT 2904.600 1704.410 2904.740 1730.075 ;
        RECT 2525.040 1704.090 2525.300 1704.410 ;
        RECT 2904.540 1704.090 2904.800 1704.410 ;
        RECT 2525.100 1703.925 2525.240 1704.090 ;
        RECT 2525.030 1703.555 2525.310 1703.925 ;
      LAYER via2 ;
        RECT 2904.530 1730.120 2904.810 1730.400 ;
        RECT 2525.030 1703.600 2525.310 1703.880 ;
      LAYER met3 ;
        RECT 2904.505 1730.410 2904.835 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2904.505 1730.110 2924.800 1730.410 ;
        RECT 2904.505 1730.095 2904.835 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2506.000 1703.890 2510.000 1704.040 ;
        RECT 2525.005 1703.890 2525.335 1703.905 ;
        RECT 2506.000 1703.590 2525.335 1703.890 ;
        RECT 2506.000 1703.440 2510.000 1703.590 ;
        RECT 2525.005 1703.575 2525.335 1703.590 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1876.700 2525.330 1876.760 ;
        RECT 2901.750 1876.700 2902.070 1876.760 ;
        RECT 2525.010 1876.560 2902.070 1876.700 ;
        RECT 2525.010 1876.500 2525.330 1876.560 ;
        RECT 2901.750 1876.500 2902.070 1876.560 ;
      LAYER via ;
        RECT 2525.040 1876.500 2525.300 1876.760 ;
        RECT 2901.780 1876.500 2902.040 1876.760 ;
      LAYER met2 ;
        RECT 2901.770 1964.675 2902.050 1965.045 ;
        RECT 2901.840 1876.790 2901.980 1964.675 ;
        RECT 2525.040 1876.470 2525.300 1876.790 ;
        RECT 2901.780 1876.470 2902.040 1876.790 ;
        RECT 2525.100 1870.525 2525.240 1876.470 ;
        RECT 2525.030 1870.155 2525.310 1870.525 ;
      LAYER via2 ;
        RECT 2901.770 1964.720 2902.050 1965.000 ;
        RECT 2525.030 1870.200 2525.310 1870.480 ;
      LAYER met3 ;
        RECT 2901.745 1965.010 2902.075 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2901.745 1964.710 2924.800 1965.010 ;
        RECT 2901.745 1964.695 2902.075 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2506.000 1870.490 2510.000 1870.640 ;
        RECT 2525.005 1870.490 2525.335 1870.505 ;
        RECT 2506.000 1870.190 2525.335 1870.490 ;
        RECT 2506.000 1870.040 2510.000 1870.190 ;
        RECT 2525.005 1870.175 2525.335 1870.190 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 2194.600 2522.110 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2521.790 2194.460 2901.150 2194.600 ;
        RECT 2521.790 2194.400 2522.110 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2521.820 2194.400 2522.080 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2521.820 2194.370 2522.080 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2521.880 2037.125 2522.020 2194.370 ;
        RECT 2521.810 2036.755 2522.090 2037.125 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2521.810 2036.800 2522.090 2037.080 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2506.000 2037.090 2510.000 2037.240 ;
        RECT 2521.785 2037.090 2522.115 2037.105 ;
        RECT 2506.000 2036.790 2522.115 2037.090 ;
        RECT 2506.000 2036.640 2510.000 2036.790 ;
        RECT 2521.785 2036.775 2522.115 2036.790 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 206.960 2522.570 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2522.250 206.820 2901.150 206.960 ;
        RECT 2522.250 206.760 2522.570 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2522.280 206.760 2522.540 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2522.270 648.195 2522.550 648.565 ;
        RECT 2522.340 207.050 2522.480 648.195 ;
        RECT 2522.280 206.730 2522.540 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2522.270 648.240 2522.550 648.520 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2506.000 648.530 2510.000 648.680 ;
        RECT 2522.245 648.530 2522.575 648.545 ;
        RECT 2506.000 648.230 2522.575 648.530 ;
        RECT 2506.000 648.080 2510.000 648.230 ;
        RECT 2522.245 648.215 2522.575 648.230 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2535.590 2546.500 2535.910 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2535.590 2546.360 2901.150 2546.500 ;
        RECT 2535.590 2546.300 2535.910 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
        RECT 2519.030 2318.360 2519.350 2318.420 ;
        RECT 2535.590 2318.360 2535.910 2318.420 ;
        RECT 2519.030 2318.220 2535.910 2318.360 ;
        RECT 2519.030 2318.160 2519.350 2318.220 ;
        RECT 2535.590 2318.160 2535.910 2318.220 ;
      LAYER via ;
        RECT 2535.620 2546.300 2535.880 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
        RECT 2519.060 2318.160 2519.320 2318.420 ;
        RECT 2535.620 2318.160 2535.880 2318.420 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2535.620 2546.270 2535.880 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2535.680 2318.450 2535.820 2546.270 ;
        RECT 2519.060 2318.130 2519.320 2318.450 ;
        RECT 2535.620 2318.130 2535.880 2318.450 ;
        RECT 2519.120 2315.245 2519.260 2318.130 ;
        RECT 2519.050 2314.875 2519.330 2315.245 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2519.050 2314.920 2519.330 2315.200 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2506.000 2315.210 2510.000 2315.360 ;
        RECT 2519.025 2315.210 2519.355 2315.225 ;
        RECT 2506.000 2314.910 2519.355 2315.210 ;
        RECT 2506.000 2314.760 2510.000 2314.910 ;
        RECT 2519.025 2314.895 2519.355 2314.910 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 2781.100 2522.110 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2521.790 2780.960 2901.150 2781.100 ;
        RECT 2521.790 2780.900 2522.110 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2521.820 2780.900 2522.080 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2521.820 2780.870 2522.080 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2521.880 2481.845 2522.020 2780.870 ;
        RECT 2521.810 2481.475 2522.090 2481.845 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2521.810 2481.520 2522.090 2481.800 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2506.000 2481.810 2510.000 2481.960 ;
        RECT 2521.785 2481.810 2522.115 2481.825 ;
        RECT 2506.000 2481.510 2522.115 2481.810 ;
        RECT 2506.000 2481.360 2510.000 2481.510 ;
        RECT 2521.785 2481.495 2522.115 2481.510 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2825.390 3015.700 2825.710 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2825.390 3015.560 2901.150 3015.700 ;
        RECT 2825.390 3015.500 2825.710 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2525.010 2649.520 2525.330 2649.580 ;
        RECT 2825.390 2649.520 2825.710 2649.580 ;
        RECT 2525.010 2649.380 2825.710 2649.520 ;
        RECT 2525.010 2649.320 2525.330 2649.380 ;
        RECT 2825.390 2649.320 2825.710 2649.380 ;
      LAYER via ;
        RECT 2825.420 3015.500 2825.680 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2525.040 2649.320 2525.300 2649.580 ;
        RECT 2825.420 2649.320 2825.680 2649.580 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2825.420 3015.470 2825.680 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2825.480 2649.610 2825.620 3015.470 ;
        RECT 2525.040 2649.290 2525.300 2649.610 ;
        RECT 2825.420 2649.290 2825.680 2649.610 ;
        RECT 2525.100 2648.445 2525.240 2649.290 ;
        RECT 2525.030 2648.075 2525.310 2648.445 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2525.030 2648.120 2525.310 2648.400 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2506.000 2648.410 2510.000 2648.560 ;
        RECT 2525.005 2648.410 2525.335 2648.425 ;
        RECT 2506.000 2648.110 2525.335 2648.410 ;
        RECT 2506.000 2647.960 2510.000 2648.110 ;
        RECT 2525.005 2648.095 2525.335 2648.110 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2645.990 3250.300 2646.310 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2645.990 3250.160 2901.150 3250.300 ;
        RECT 2645.990 3250.100 2646.310 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2525.010 2815.100 2525.330 2815.160 ;
        RECT 2645.990 2815.100 2646.310 2815.160 ;
        RECT 2525.010 2814.960 2646.310 2815.100 ;
        RECT 2525.010 2814.900 2525.330 2814.960 ;
        RECT 2645.990 2814.900 2646.310 2814.960 ;
      LAYER via ;
        RECT 2646.020 3250.100 2646.280 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2525.040 2814.900 2525.300 2815.160 ;
        RECT 2646.020 2814.900 2646.280 2815.160 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2646.020 3250.070 2646.280 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2646.080 2815.190 2646.220 3250.070 ;
        RECT 2525.040 2815.045 2525.300 2815.190 ;
        RECT 2525.030 2814.675 2525.310 2815.045 ;
        RECT 2646.020 2814.870 2646.280 2815.190 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2525.030 2814.720 2525.310 2815.000 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2506.000 2815.010 2510.000 2815.160 ;
        RECT 2525.005 2815.010 2525.335 2815.025 ;
        RECT 2506.000 2814.710 2525.335 2815.010 ;
        RECT 2506.000 2814.560 2510.000 2814.710 ;
        RECT 2525.005 2814.695 2525.335 2814.710 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2694.290 3484.900 2694.610 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2694.290 3484.760 2901.150 3484.900 ;
        RECT 2694.290 3484.700 2694.610 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2525.010 2987.480 2525.330 2987.540 ;
        RECT 2694.290 2987.480 2694.610 2987.540 ;
        RECT 2525.010 2987.340 2694.610 2987.480 ;
        RECT 2525.010 2987.280 2525.330 2987.340 ;
        RECT 2694.290 2987.280 2694.610 2987.340 ;
      LAYER via ;
        RECT 2694.320 3484.700 2694.580 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2525.040 2987.280 2525.300 2987.540 ;
        RECT 2694.320 2987.280 2694.580 2987.540 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2694.320 3484.670 2694.580 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2694.380 2987.570 2694.520 3484.670 ;
        RECT 2525.040 2987.250 2525.300 2987.570 ;
        RECT 2694.320 2987.250 2694.580 2987.570 ;
        RECT 2525.100 2981.645 2525.240 2987.250 ;
        RECT 2525.030 2981.275 2525.310 2981.645 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2525.030 2981.320 2525.310 2981.600 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2506.000 2981.610 2510.000 2981.760 ;
        RECT 2525.005 2981.610 2525.335 2981.625 ;
        RECT 2506.000 2981.310 2525.335 2981.610 ;
        RECT 2506.000 2981.160 2510.000 2981.310 ;
        RECT 2525.005 2981.295 2525.335 2981.310 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2314.790 3018.760 2315.110 3018.820 ;
        RECT 2635.870 3018.760 2636.190 3018.820 ;
        RECT 2314.790 3018.620 2636.190 3018.760 ;
        RECT 2314.790 3018.560 2315.110 3018.620 ;
        RECT 2635.870 3018.560 2636.190 3018.620 ;
      LAYER via ;
        RECT 2314.820 3018.560 2315.080 3018.820 ;
        RECT 2635.900 3018.560 2636.160 3018.820 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3018.850 2636.100 3517.600 ;
        RECT 2314.820 3018.530 2315.080 3018.850 ;
        RECT 2635.900 3018.530 2636.160 3018.850 ;
        RECT 2314.880 3010.000 2315.020 3018.530 ;
        RECT 2314.880 3009.340 2315.230 3010.000 ;
        RECT 2314.950 3006.000 2315.230 3009.340 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2081.570 3018.760 2081.890 3018.820 ;
        RECT 2311.570 3018.760 2311.890 3018.820 ;
        RECT 2081.570 3018.620 2311.890 3018.760 ;
        RECT 2081.570 3018.560 2081.890 3018.620 ;
        RECT 2311.570 3018.560 2311.890 3018.620 ;
      LAYER via ;
        RECT 2081.600 3018.560 2081.860 3018.820 ;
        RECT 2311.600 3018.560 2311.860 3018.820 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3018.850 2311.800 3517.600 ;
        RECT 2081.600 3018.530 2081.860 3018.850 ;
        RECT 2311.600 3018.530 2311.860 3018.850 ;
        RECT 2081.660 3010.000 2081.800 3018.530 ;
        RECT 2081.660 3009.340 2082.010 3010.000 ;
        RECT 2081.730 3006.000 2082.010 3009.340 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.350 3018.760 1848.670 3018.820 ;
        RECT 1987.270 3018.760 1987.590 3018.820 ;
        RECT 1848.350 3018.620 1987.590 3018.760 ;
        RECT 1848.350 3018.560 1848.670 3018.620 ;
        RECT 1987.270 3018.560 1987.590 3018.620 ;
      LAYER via ;
        RECT 1848.380 3018.560 1848.640 3018.820 ;
        RECT 1987.300 3018.560 1987.560 3018.820 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3018.850 1987.500 3517.600 ;
        RECT 1848.380 3018.530 1848.640 3018.850 ;
        RECT 1987.300 3018.530 1987.560 3018.850 ;
        RECT 1848.440 3010.000 1848.580 3018.530 ;
        RECT 1848.440 3009.340 1848.790 3010.000 ;
        RECT 1848.510 3006.000 1848.790 3009.340 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.070 3487.960 1656.390 3488.020 ;
        RECT 1662.510 3487.960 1662.830 3488.020 ;
        RECT 1656.070 3487.820 1662.830 3487.960 ;
        RECT 1656.070 3487.760 1656.390 3487.820 ;
        RECT 1662.510 3487.760 1662.830 3487.820 ;
        RECT 1615.130 3018.760 1615.450 3018.820 ;
        RECT 1656.070 3018.760 1656.390 3018.820 ;
        RECT 1615.130 3018.620 1656.390 3018.760 ;
        RECT 1615.130 3018.560 1615.450 3018.620 ;
        RECT 1656.070 3018.560 1656.390 3018.620 ;
      LAYER via ;
        RECT 1656.100 3487.760 1656.360 3488.020 ;
        RECT 1662.540 3487.760 1662.800 3488.020 ;
        RECT 1615.160 3018.560 1615.420 3018.820 ;
        RECT 1656.100 3018.560 1656.360 3018.820 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3488.050 1662.740 3517.600 ;
        RECT 1656.100 3487.730 1656.360 3488.050 ;
        RECT 1662.540 3487.730 1662.800 3488.050 ;
        RECT 1656.160 3018.850 1656.300 3487.730 ;
        RECT 1615.160 3018.530 1615.420 3018.850 ;
        RECT 1656.100 3018.530 1656.360 3018.850 ;
        RECT 1615.220 3010.000 1615.360 3018.530 ;
        RECT 1615.220 3009.340 1615.570 3010.000 ;
        RECT 1615.290 3006.000 1615.570 3009.340 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3018.760 1338.530 3018.820 ;
        RECT 1381.450 3018.760 1381.770 3018.820 ;
        RECT 1338.210 3018.620 1381.770 3018.760 ;
        RECT 1338.210 3018.560 1338.530 3018.620 ;
        RECT 1381.450 3018.560 1381.770 3018.620 ;
      LAYER via ;
        RECT 1338.240 3018.560 1338.500 3018.820 ;
        RECT 1381.480 3018.560 1381.740 3018.820 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3018.850 1338.440 3517.600 ;
        RECT 1338.240 3018.530 1338.500 3018.850 ;
        RECT 1381.480 3018.530 1381.740 3018.850 ;
        RECT 1381.540 3010.000 1381.680 3018.530 ;
        RECT 1381.540 3009.340 1381.890 3010.000 ;
        RECT 1381.610 3006.000 1381.890 3009.340 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 441.560 2523.030 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2522.710 441.420 2901.150 441.560 ;
        RECT 2522.710 441.360 2523.030 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2522.740 441.360 2523.000 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2522.730 814.795 2523.010 815.165 ;
        RECT 2522.800 441.650 2522.940 814.795 ;
        RECT 2522.740 441.330 2523.000 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2522.730 814.840 2523.010 815.120 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2506.000 815.130 2510.000 815.280 ;
        RECT 2522.705 815.130 2523.035 815.145 ;
        RECT 2506.000 814.830 2523.035 815.130 ;
        RECT 2506.000 814.680 2510.000 814.830 ;
        RECT 2522.705 814.815 2523.035 814.830 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3019.100 1014.230 3019.160 ;
        RECT 1148.230 3019.100 1148.550 3019.160 ;
        RECT 1013.910 3018.960 1148.550 3019.100 ;
        RECT 1013.910 3018.900 1014.230 3018.960 ;
        RECT 1148.230 3018.900 1148.550 3018.960 ;
      LAYER via ;
        RECT 1013.940 3018.900 1014.200 3019.160 ;
        RECT 1148.260 3018.900 1148.520 3019.160 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3019.190 1014.140 3517.600 ;
        RECT 1013.940 3018.870 1014.200 3019.190 ;
        RECT 1148.260 3018.870 1148.520 3019.190 ;
        RECT 1148.320 3010.000 1148.460 3018.870 ;
        RECT 1148.320 3009.340 1148.670 3010.000 ;
        RECT 1148.390 3006.000 1148.670 3009.340 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3270.700 689.010 3270.760 ;
        RECT 689.610 3270.700 689.930 3270.760 ;
        RECT 688.690 3270.560 689.930 3270.700 ;
        RECT 688.690 3270.500 689.010 3270.560 ;
        RECT 689.610 3270.500 689.930 3270.560 ;
        RECT 688.690 3174.140 689.010 3174.200 ;
        RECT 689.610 3174.140 689.930 3174.200 ;
        RECT 688.690 3174.000 689.930 3174.140 ;
        RECT 688.690 3173.940 689.010 3174.000 ;
        RECT 689.610 3173.940 689.930 3174.000 ;
        RECT 688.690 3077.580 689.010 3077.640 ;
        RECT 689.610 3077.580 689.930 3077.640 ;
        RECT 688.690 3077.440 689.930 3077.580 ;
        RECT 688.690 3077.380 689.010 3077.440 ;
        RECT 689.610 3077.380 689.930 3077.440 ;
        RECT 688.690 3019.100 689.010 3019.160 ;
        RECT 915.010 3019.100 915.330 3019.160 ;
        RECT 688.690 3018.960 915.330 3019.100 ;
        RECT 688.690 3018.900 689.010 3018.960 ;
        RECT 915.010 3018.900 915.330 3018.960 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3270.500 688.980 3270.760 ;
        RECT 689.640 3270.500 689.900 3270.760 ;
        RECT 688.720 3173.940 688.980 3174.200 ;
        RECT 689.640 3173.940 689.900 3174.200 ;
        RECT 688.720 3077.380 688.980 3077.640 ;
        RECT 689.640 3077.380 689.900 3077.640 ;
        RECT 688.720 3018.900 688.980 3019.160 ;
        RECT 915.040 3018.900 915.300 3019.160 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3270.790 688.920 3318.670 ;
        RECT 688.720 3270.470 688.980 3270.790 ;
        RECT 689.640 3270.470 689.900 3270.790 ;
        RECT 689.700 3222.250 689.840 3270.470 ;
        RECT 688.780 3222.110 689.840 3222.250 ;
        RECT 688.780 3174.230 688.920 3222.110 ;
        RECT 688.720 3173.910 688.980 3174.230 ;
        RECT 689.640 3173.910 689.900 3174.230 ;
        RECT 689.700 3125.690 689.840 3173.910 ;
        RECT 688.780 3125.550 689.840 3125.690 ;
        RECT 688.780 3077.670 688.920 3125.550 ;
        RECT 688.720 3077.350 688.980 3077.670 ;
        RECT 689.640 3077.350 689.900 3077.670 ;
        RECT 689.700 3029.130 689.840 3077.350 ;
        RECT 688.780 3028.990 689.840 3029.130 ;
        RECT 688.780 3019.190 688.920 3028.990 ;
        RECT 688.720 3018.870 688.980 3019.190 ;
        RECT 915.040 3018.870 915.300 3019.190 ;
        RECT 915.100 3010.000 915.240 3018.870 ;
        RECT 915.100 3009.340 915.450 3010.000 ;
        RECT 915.170 3006.000 915.450 3009.340 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
        RECT 364.925 3236.205 365.095 3284.315 ;
        RECT 364.005 3139.645 364.175 3187.755 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
        RECT 364.925 3284.145 365.095 3284.315 ;
        RECT 364.005 3187.585 364.175 3187.755 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 364.390 3298.240 364.710 3298.300 ;
        RECT 365.310 3298.240 365.630 3298.300 ;
        RECT 364.390 3298.100 365.630 3298.240 ;
        RECT 364.390 3298.040 364.710 3298.100 ;
        RECT 365.310 3298.040 365.630 3298.100 ;
        RECT 364.865 3284.300 365.155 3284.345 ;
        RECT 365.310 3284.300 365.630 3284.360 ;
        RECT 364.865 3284.160 365.630 3284.300 ;
        RECT 364.865 3284.115 365.155 3284.160 ;
        RECT 365.310 3284.100 365.630 3284.160 ;
        RECT 364.850 3236.360 365.170 3236.420 ;
        RECT 364.655 3236.220 365.170 3236.360 ;
        RECT 364.850 3236.160 365.170 3236.220 ;
        RECT 364.850 3202.020 365.170 3202.080 ;
        RECT 364.020 3201.880 365.170 3202.020 ;
        RECT 364.020 3201.400 364.160 3201.880 ;
        RECT 364.850 3201.820 365.170 3201.880 ;
        RECT 363.930 3201.140 364.250 3201.400 ;
        RECT 363.930 3187.740 364.250 3187.800 ;
        RECT 363.735 3187.600 364.250 3187.740 ;
        RECT 363.930 3187.540 364.250 3187.600 ;
        RECT 363.945 3139.800 364.235 3139.845 ;
        RECT 365.310 3139.800 365.630 3139.860 ;
        RECT 363.945 3139.660 365.630 3139.800 ;
        RECT 363.945 3139.615 364.235 3139.660 ;
        RECT 365.310 3139.600 365.630 3139.660 ;
        RECT 365.310 3019.780 365.630 3019.840 ;
        RECT 681.790 3019.780 682.110 3019.840 ;
        RECT 365.310 3019.640 682.110 3019.780 ;
        RECT 365.310 3019.580 365.630 3019.640 ;
        RECT 681.790 3019.580 682.110 3019.640 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 364.420 3298.040 364.680 3298.300 ;
        RECT 365.340 3298.040 365.600 3298.300 ;
        RECT 365.340 3284.100 365.600 3284.360 ;
        RECT 364.880 3236.160 365.140 3236.420 ;
        RECT 364.880 3201.820 365.140 3202.080 ;
        RECT 363.960 3201.140 364.220 3201.400 ;
        RECT 363.960 3187.540 364.220 3187.800 ;
        RECT 365.340 3139.600 365.600 3139.860 ;
        RECT 365.340 3019.580 365.600 3019.840 ;
        RECT 681.820 3019.580 682.080 3019.840 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.330 364.620 3298.410 ;
        RECT 364.020 3298.270 364.680 3298.330 ;
        RECT 364.420 3298.010 364.680 3298.270 ;
        RECT 365.340 3298.010 365.600 3298.330 ;
        RECT 365.400 3284.390 365.540 3298.010 ;
        RECT 365.340 3284.070 365.600 3284.390 ;
        RECT 364.880 3236.130 365.140 3236.450 ;
        RECT 364.940 3202.110 365.080 3236.130 ;
        RECT 364.880 3201.790 365.140 3202.110 ;
        RECT 363.960 3201.110 364.220 3201.430 ;
        RECT 364.020 3187.830 364.160 3201.110 ;
        RECT 363.960 3187.510 364.220 3187.830 ;
        RECT 365.340 3139.570 365.600 3139.890 ;
        RECT 365.400 3019.870 365.540 3139.570 ;
        RECT 365.340 3019.550 365.600 3019.870 ;
        RECT 681.820 3019.550 682.080 3019.870 ;
        RECT 681.880 3010.000 682.020 3019.550 ;
        RECT 681.880 3009.340 682.230 3010.000 ;
        RECT 681.950 3006.000 682.230 3009.340 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 3018.760 40.410 3018.820 ;
        RECT 448.570 3018.760 448.890 3018.820 ;
        RECT 40.090 3018.620 448.890 3018.760 ;
        RECT 40.090 3018.560 40.410 3018.620 ;
        RECT 448.570 3018.560 448.890 3018.620 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 3018.560 40.380 3018.820 ;
        RECT 448.600 3018.560 448.860 3018.820 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 3018.850 40.320 3028.990 ;
        RECT 40.120 3018.530 40.380 3018.850 ;
        RECT 448.600 3018.530 448.860 3018.850 ;
        RECT 448.660 3010.000 448.800 3018.530 ;
        RECT 448.660 3009.340 449.010 3010.000 ;
        RECT 448.730 3006.000 449.010 3009.340 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 51.590 3263.900 51.910 3263.960 ;
        RECT 15.250 3263.760 51.910 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 51.590 3263.700 51.910 3263.760 ;
        RECT 51.590 2863.380 51.910 2863.440 ;
        RECT 393.370 2863.380 393.690 2863.440 ;
        RECT 51.590 2863.240 393.690 2863.380 ;
        RECT 51.590 2863.180 51.910 2863.240 ;
        RECT 393.370 2863.180 393.690 2863.240 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 51.620 3263.700 51.880 3263.960 ;
        RECT 51.620 2863.180 51.880 2863.440 ;
        RECT 393.400 2863.180 393.660 2863.440 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 51.620 3263.670 51.880 3263.990 ;
        RECT 51.680 2863.470 51.820 3263.670 ;
        RECT 51.620 2863.150 51.880 2863.470 ;
        RECT 393.400 2863.150 393.660 2863.470 ;
        RECT 393.460 2860.605 393.600 2863.150 ;
        RECT 393.390 2860.235 393.670 2860.605 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 393.390 2860.280 393.670 2860.560 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 393.365 2860.570 393.695 2860.585 ;
        RECT 410.000 2860.570 414.000 2860.720 ;
        RECT 393.365 2860.270 414.000 2860.570 ;
        RECT 393.365 2860.255 393.695 2860.270 ;
        RECT 410.000 2860.120 414.000 2860.270 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 65.390 2974.220 65.710 2974.280 ;
        RECT 16.630 2974.080 65.710 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 65.390 2974.020 65.710 2974.080 ;
        RECT 65.390 2683.860 65.710 2683.920 ;
        RECT 393.370 2683.860 393.690 2683.920 ;
        RECT 65.390 2683.720 393.690 2683.860 ;
        RECT 65.390 2683.660 65.710 2683.720 ;
        RECT 393.370 2683.660 393.690 2683.720 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 65.420 2974.020 65.680 2974.280 ;
        RECT 65.420 2683.660 65.680 2683.920 ;
        RECT 393.400 2683.660 393.660 2683.920 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 65.420 2973.990 65.680 2974.310 ;
        RECT 65.480 2683.950 65.620 2973.990 ;
        RECT 65.420 2683.630 65.680 2683.950 ;
        RECT 393.400 2683.630 393.660 2683.950 ;
        RECT 393.460 2681.765 393.600 2683.630 ;
        RECT 393.390 2681.395 393.670 2681.765 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
        RECT 393.390 2681.440 393.670 2681.720 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
        RECT 393.365 2681.730 393.695 2681.745 ;
        RECT 410.000 2681.730 414.000 2681.880 ;
        RECT 393.365 2681.430 414.000 2681.730 ;
        RECT 393.365 2681.415 393.695 2681.430 ;
        RECT 410.000 2681.280 414.000 2681.430 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2504.680 17.870 2504.740 ;
        RECT 393.370 2504.680 393.690 2504.740 ;
        RECT 17.550 2504.540 393.690 2504.680 ;
        RECT 17.550 2504.480 17.870 2504.540 ;
        RECT 393.370 2504.480 393.690 2504.540 ;
      LAYER via ;
        RECT 17.580 2504.480 17.840 2504.740 ;
        RECT 393.400 2504.480 393.660 2504.740 ;
      LAYER met2 ;
        RECT 17.570 2692.955 17.850 2693.325 ;
        RECT 17.640 2504.770 17.780 2692.955 ;
        RECT 17.580 2504.450 17.840 2504.770 ;
        RECT 393.400 2504.450 393.660 2504.770 ;
        RECT 393.460 2503.605 393.600 2504.450 ;
        RECT 393.390 2503.235 393.670 2503.605 ;
      LAYER via2 ;
        RECT 17.570 2693.000 17.850 2693.280 ;
        RECT 393.390 2503.280 393.670 2503.560 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.545 2693.290 17.875 2693.305 ;
        RECT -4.800 2692.990 17.875 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.545 2692.975 17.875 2692.990 ;
        RECT 393.365 2503.570 393.695 2503.585 ;
        RECT 410.000 2503.570 414.000 2503.720 ;
        RECT 393.365 2503.270 414.000 2503.570 ;
        RECT 393.365 2503.255 393.695 2503.270 ;
        RECT 410.000 2503.120 414.000 2503.270 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2325.160 17.410 2325.220 ;
        RECT 393.370 2325.160 393.690 2325.220 ;
        RECT 17.090 2325.020 393.690 2325.160 ;
        RECT 17.090 2324.960 17.410 2325.020 ;
        RECT 393.370 2324.960 393.690 2325.020 ;
      LAYER via ;
        RECT 17.120 2324.960 17.380 2325.220 ;
        RECT 393.400 2324.960 393.660 2325.220 ;
      LAYER met2 ;
        RECT 17.110 2405.315 17.390 2405.685 ;
        RECT 17.180 2325.250 17.320 2405.315 ;
        RECT 17.120 2324.930 17.380 2325.250 ;
        RECT 393.400 2324.930 393.660 2325.250 ;
        RECT 393.460 2324.765 393.600 2324.930 ;
        RECT 393.390 2324.395 393.670 2324.765 ;
      LAYER via2 ;
        RECT 17.110 2405.360 17.390 2405.640 ;
        RECT 393.390 2324.440 393.670 2324.720 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 17.085 2405.650 17.415 2405.665 ;
        RECT -4.800 2405.350 17.415 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 17.085 2405.335 17.415 2405.350 ;
        RECT 393.365 2324.730 393.695 2324.745 ;
        RECT 410.000 2324.730 414.000 2324.880 ;
        RECT 393.365 2324.430 414.000 2324.730 ;
        RECT 393.365 2324.415 393.695 2324.430 ;
        RECT 410.000 2324.280 414.000 2324.430 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 393.370 2125.240 393.690 2125.300 ;
        RECT 16.170 2125.100 393.690 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 393.370 2125.040 393.690 2125.100 ;
      LAYER via ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 393.400 2125.040 393.660 2125.300 ;
      LAYER met2 ;
        RECT 393.390 2146.235 393.670 2146.605 ;
        RECT 393.460 2125.330 393.600 2146.235 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 393.400 2125.010 393.660 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 393.390 2146.280 393.670 2146.560 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT 393.365 2146.570 393.695 2146.585 ;
        RECT 410.000 2146.570 414.000 2146.720 ;
        RECT 393.365 2146.270 414.000 2146.570 ;
        RECT 393.365 2146.255 393.695 2146.270 ;
        RECT 410.000 2146.120 414.000 2146.270 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 396.590 1835.220 396.910 1835.280 ;
        RECT 15.710 1835.080 396.910 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 396.590 1835.020 396.910 1835.080 ;
      LAYER via ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 396.620 1835.020 396.880 1835.280 ;
      LAYER met2 ;
        RECT 396.610 1967.395 396.890 1967.765 ;
        RECT 396.680 1835.310 396.820 1967.395 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 396.620 1834.990 396.880 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 396.610 1967.440 396.890 1967.720 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 396.585 1967.730 396.915 1967.745 ;
        RECT 410.000 1967.730 414.000 1967.880 ;
        RECT 396.585 1967.430 414.000 1967.730 ;
        RECT 396.585 1967.415 396.915 1967.430 ;
        RECT 410.000 1967.280 414.000 1967.430 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 676.160 2522.110 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2521.790 676.020 2901.150 676.160 ;
        RECT 2521.790 675.960 2522.110 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2521.820 675.960 2522.080 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2521.810 981.395 2522.090 981.765 ;
        RECT 2521.880 676.250 2522.020 981.395 ;
        RECT 2521.820 675.930 2522.080 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2521.810 981.440 2522.090 981.720 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2506.000 981.730 2510.000 981.880 ;
        RECT 2521.785 981.730 2522.115 981.745 ;
        RECT 2506.000 981.430 2522.115 981.730 ;
        RECT 2506.000 981.280 2510.000 981.430 ;
        RECT 2521.785 981.415 2522.115 981.430 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 397.050 1545.540 397.370 1545.600 ;
        RECT 16.630 1545.400 397.370 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 397.050 1545.340 397.370 1545.400 ;
      LAYER via ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 397.080 1545.340 397.340 1545.600 ;
      LAYER met2 ;
        RECT 397.070 1789.235 397.350 1789.605 ;
        RECT 397.140 1545.630 397.280 1789.235 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 397.080 1545.310 397.340 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 397.070 1789.280 397.350 1789.560 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 397.045 1789.570 397.375 1789.585 ;
        RECT 410.000 1789.570 414.000 1789.720 ;
        RECT 397.045 1789.270 414.000 1789.570 ;
        RECT 397.045 1789.255 397.375 1789.270 ;
        RECT 410.000 1789.120 414.000 1789.270 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 397.970 1331.680 398.290 1331.740 ;
        RECT 15.710 1331.540 398.290 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 397.970 1331.480 398.290 1331.540 ;
      LAYER via ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 398.000 1331.480 398.260 1331.740 ;
      LAYER met2 ;
        RECT 397.990 1610.395 398.270 1610.765 ;
        RECT 398.060 1331.770 398.200 1610.395 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 398.000 1331.450 398.260 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 397.990 1610.440 398.270 1610.720 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
        RECT 397.965 1610.730 398.295 1610.745 ;
        RECT 410.000 1610.730 414.000 1610.880 ;
        RECT 397.965 1610.430 414.000 1610.730 ;
        RECT 397.965 1610.415 398.295 1610.430 ;
        RECT 410.000 1610.280 414.000 1610.430 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 15.705 1328.215 16.035 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 396.590 1117.820 396.910 1117.880 ;
        RECT 15.710 1117.680 396.910 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 396.590 1117.620 396.910 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 396.620 1117.620 396.880 1117.880 ;
      LAYER met2 ;
        RECT 396.610 1431.555 396.890 1431.925 ;
        RECT 396.680 1117.910 396.820 1431.555 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 396.620 1117.590 396.880 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 396.610 1431.600 396.890 1431.880 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 396.585 1431.890 396.915 1431.905 ;
        RECT 410.000 1431.890 414.000 1432.040 ;
        RECT 396.585 1431.590 414.000 1431.890 ;
        RECT 396.585 1431.575 396.915 1431.590 ;
        RECT 410.000 1431.440 414.000 1431.590 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 397.510 903.960 397.830 904.020 ;
        RECT 16.170 903.820 397.830 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 397.510 903.760 397.830 903.820 ;
      LAYER via ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 397.540 903.760 397.800 904.020 ;
      LAYER met2 ;
        RECT 397.530 1253.395 397.810 1253.765 ;
        RECT 397.600 904.050 397.740 1253.395 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 397.540 903.730 397.800 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 397.530 1253.440 397.810 1253.720 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 397.505 1253.730 397.835 1253.745 ;
        RECT 410.000 1253.730 414.000 1253.880 ;
        RECT 397.505 1253.430 414.000 1253.730 ;
        RECT 397.505 1253.415 397.835 1253.430 ;
        RECT 410.000 1253.280 414.000 1253.430 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 396.590 682.960 396.910 683.020 ;
        RECT 16.170 682.820 396.910 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 396.590 682.760 396.910 682.820 ;
      LAYER via ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 396.620 682.760 396.880 683.020 ;
      LAYER met2 ;
        RECT 396.610 1074.555 396.890 1074.925 ;
        RECT 396.680 683.050 396.820 1074.555 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 396.620 682.730 396.880 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 396.610 1074.600 396.890 1074.880 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 396.585 1074.890 396.915 1074.905 ;
        RECT 410.000 1074.890 414.000 1075.040 ;
        RECT 396.585 1074.590 414.000 1074.890 ;
        RECT 396.585 1074.575 396.915 1074.590 ;
        RECT 410.000 1074.440 414.000 1074.590 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 398.430 469.100 398.750 469.160 ;
        RECT 17.090 468.960 398.750 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 398.430 468.900 398.750 468.960 ;
      LAYER via ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 398.460 468.900 398.720 469.160 ;
      LAYER met2 ;
        RECT 398.450 896.395 398.730 896.765 ;
        RECT 398.520 469.190 398.660 896.395 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 398.460 468.870 398.720 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 398.450 896.440 398.730 896.720 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 398.425 896.730 398.755 896.745 ;
        RECT 410.000 896.730 414.000 896.880 ;
        RECT 398.425 896.430 414.000 896.730 ;
        RECT 398.425 896.415 398.755 896.430 ;
        RECT 410.000 896.280 414.000 896.430 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 397.510 255.240 397.830 255.300 ;
        RECT 17.090 255.100 397.830 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 397.510 255.040 397.830 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 397.540 255.040 397.800 255.300 ;
      LAYER met2 ;
        RECT 397.530 717.555 397.810 717.925 ;
        RECT 397.600 255.330 397.740 717.555 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 397.540 255.010 397.800 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 397.530 717.600 397.810 717.880 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 397.505 717.890 397.835 717.905 ;
        RECT 410.000 717.890 414.000 718.040 ;
        RECT 397.505 717.590 414.000 717.890 ;
        RECT 397.505 717.575 397.835 717.590 ;
        RECT 410.000 717.440 414.000 717.590 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 396.590 41.380 396.910 41.440 ;
        RECT 17.090 41.240 396.910 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 396.590 41.180 396.910 41.240 ;
      LAYER via ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 396.620 41.180 396.880 41.440 ;
      LAYER met2 ;
        RECT 396.610 539.395 396.890 539.765 ;
        RECT 396.680 41.470 396.820 539.395 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 396.620 41.150 396.880 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 396.610 539.440 396.890 539.720 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 396.585 539.730 396.915 539.745 ;
        RECT 410.000 539.730 414.000 539.880 ;
        RECT 396.585 539.430 414.000 539.730 ;
        RECT 396.585 539.415 396.915 539.430 ;
        RECT 410.000 539.280 414.000 539.430 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 910.760 2523.030 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2522.710 910.620 2901.150 910.760 ;
        RECT 2522.710 910.560 2523.030 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2522.740 910.560 2523.000 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2522.730 1147.995 2523.010 1148.365 ;
        RECT 2522.800 910.850 2522.940 1147.995 ;
        RECT 2522.740 910.530 2523.000 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2522.730 1148.040 2523.010 1148.320 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2506.000 1148.330 2510.000 1148.480 ;
        RECT 2522.705 1148.330 2523.035 1148.345 ;
        RECT 2506.000 1148.030 2523.035 1148.330 ;
        RECT 2506.000 1147.880 2510.000 1148.030 ;
        RECT 2522.705 1148.015 2523.035 1148.030 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 1145.360 2522.570 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2522.250 1145.220 2901.150 1145.360 ;
        RECT 2522.250 1145.160 2522.570 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2522.280 1145.160 2522.540 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2522.270 1314.595 2522.550 1314.965 ;
        RECT 2522.340 1145.450 2522.480 1314.595 ;
        RECT 2522.280 1145.130 2522.540 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2522.270 1314.640 2522.550 1314.920 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2506.000 1314.930 2510.000 1315.080 ;
        RECT 2522.245 1314.930 2522.575 1314.945 ;
        RECT 2506.000 1314.630 2522.575 1314.930 ;
        RECT 2506.000 1314.480 2510.000 1314.630 ;
        RECT 2522.245 1314.615 2522.575 1314.630 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1379.960 2522.110 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2521.790 1379.820 2901.150 1379.960 ;
        RECT 2521.790 1379.760 2522.110 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2521.820 1379.760 2522.080 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2521.810 1481.195 2522.090 1481.565 ;
        RECT 2521.880 1380.050 2522.020 1481.195 ;
        RECT 2521.820 1379.730 2522.080 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2521.810 1481.240 2522.090 1481.520 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2506.000 1481.530 2510.000 1481.680 ;
        RECT 2521.785 1481.530 2522.115 1481.545 ;
        RECT 2506.000 1481.230 2522.115 1481.530 ;
        RECT 2506.000 1481.080 2510.000 1481.230 ;
        RECT 2521.785 1481.215 2522.115 1481.230 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1614.560 2522.110 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2521.790 1614.420 2901.150 1614.560 ;
        RECT 2521.790 1614.360 2522.110 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2521.820 1614.360 2522.080 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2521.810 1647.795 2522.090 1648.165 ;
        RECT 2521.880 1614.650 2522.020 1647.795 ;
        RECT 2521.820 1614.330 2522.080 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2521.810 1647.840 2522.090 1648.120 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2506.000 1648.130 2510.000 1648.280 ;
        RECT 2521.785 1648.130 2522.115 1648.145 ;
        RECT 2506.000 1647.830 2522.115 1648.130 ;
        RECT 2506.000 1647.680 2510.000 1647.830 ;
        RECT 2521.785 1647.815 2522.115 1647.830 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1814.480 2525.330 1814.540 ;
        RECT 2901.290 1814.480 2901.610 1814.540 ;
        RECT 2525.010 1814.340 2901.610 1814.480 ;
        RECT 2525.010 1814.280 2525.330 1814.340 ;
        RECT 2901.290 1814.280 2901.610 1814.340 ;
      LAYER via ;
        RECT 2525.040 1814.280 2525.300 1814.540 ;
        RECT 2901.320 1814.280 2901.580 1814.540 ;
      LAYER met2 ;
        RECT 2901.310 1847.715 2901.590 1848.085 ;
        RECT 2525.030 1814.395 2525.310 1814.765 ;
        RECT 2901.380 1814.570 2901.520 1847.715 ;
        RECT 2525.040 1814.250 2525.300 1814.395 ;
        RECT 2901.320 1814.250 2901.580 1814.570 ;
      LAYER via2 ;
        RECT 2901.310 1847.760 2901.590 1848.040 ;
        RECT 2525.030 1814.440 2525.310 1814.720 ;
      LAYER met3 ;
        RECT 2901.285 1848.050 2901.615 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.285 1847.750 2924.800 1848.050 ;
        RECT 2901.285 1847.735 2901.615 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2506.000 1814.730 2510.000 1814.880 ;
        RECT 2525.005 1814.730 2525.335 1814.745 ;
        RECT 2506.000 1814.430 2525.335 1814.730 ;
        RECT 2506.000 1814.280 2510.000 1814.430 ;
        RECT 2525.005 1814.415 2525.335 1814.430 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1987.200 2525.330 1987.260 ;
        RECT 2901.750 1987.200 2902.070 1987.260 ;
        RECT 2525.010 1987.060 2902.070 1987.200 ;
        RECT 2525.010 1987.000 2525.330 1987.060 ;
        RECT 2901.750 1987.000 2902.070 1987.060 ;
      LAYER via ;
        RECT 2525.040 1987.000 2525.300 1987.260 ;
        RECT 2901.780 1987.000 2902.040 1987.260 ;
      LAYER met2 ;
        RECT 2901.770 2082.315 2902.050 2082.685 ;
        RECT 2901.840 1987.290 2901.980 2082.315 ;
        RECT 2525.040 1986.970 2525.300 1987.290 ;
        RECT 2901.780 1986.970 2902.040 1987.290 ;
        RECT 2525.100 1981.365 2525.240 1986.970 ;
        RECT 2525.030 1980.995 2525.310 1981.365 ;
      LAYER via2 ;
        RECT 2901.770 2082.360 2902.050 2082.640 ;
        RECT 2525.030 1981.040 2525.310 1981.320 ;
      LAYER met3 ;
        RECT 2901.745 2082.650 2902.075 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2901.745 2082.350 2924.800 2082.650 ;
        RECT 2901.745 2082.335 2902.075 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2506.000 1981.330 2510.000 1981.480 ;
        RECT 2525.005 1981.330 2525.335 1981.345 ;
        RECT 2506.000 1981.030 2525.335 1981.330 ;
        RECT 2506.000 1980.880 2510.000 1981.030 ;
        RECT 2525.005 1981.015 2525.335 1981.030 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2152.780 2525.330 2152.840 ;
        RECT 2901.290 2152.780 2901.610 2152.840 ;
        RECT 2525.010 2152.640 2901.610 2152.780 ;
        RECT 2525.010 2152.580 2525.330 2152.640 ;
        RECT 2901.290 2152.580 2901.610 2152.640 ;
      LAYER via ;
        RECT 2525.040 2152.580 2525.300 2152.840 ;
        RECT 2901.320 2152.580 2901.580 2152.840 ;
      LAYER met2 ;
        RECT 2901.310 2316.915 2901.590 2317.285 ;
        RECT 2901.380 2152.870 2901.520 2316.915 ;
        RECT 2525.040 2152.550 2525.300 2152.870 ;
        RECT 2901.320 2152.550 2901.580 2152.870 ;
        RECT 2525.100 2147.965 2525.240 2152.550 ;
        RECT 2525.030 2147.595 2525.310 2147.965 ;
      LAYER via2 ;
        RECT 2901.310 2316.960 2901.590 2317.240 ;
        RECT 2525.030 2147.640 2525.310 2147.920 ;
      LAYER met3 ;
        RECT 2901.285 2317.250 2901.615 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2901.285 2316.950 2924.800 2317.250 ;
        RECT 2901.285 2316.935 2901.615 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2506.000 2147.930 2510.000 2148.080 ;
        RECT 2525.005 2147.930 2525.335 2147.945 ;
        RECT 2506.000 2147.630 2525.335 2147.930 ;
        RECT 2506.000 2147.480 2510.000 2147.630 ;
        RECT 2525.005 2147.615 2525.335 2147.630 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 151.540 2522.110 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2521.790 151.400 2901.150 151.540 ;
        RECT 2521.790 151.340 2522.110 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2521.820 151.340 2522.080 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2521.810 592.435 2522.090 592.805 ;
        RECT 2521.880 151.630 2522.020 592.435 ;
        RECT 2521.820 151.310 2522.080 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2521.810 592.480 2522.090 592.760 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2506.000 592.770 2510.000 592.920 ;
        RECT 2521.785 592.770 2522.115 592.785 ;
        RECT 2506.000 592.470 2522.115 592.770 ;
        RECT 2506.000 592.320 2510.000 592.470 ;
        RECT 2521.785 592.455 2522.115 592.470 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.870 2262.940 2521.190 2263.000 ;
        RECT 2901.750 2262.940 2902.070 2263.000 ;
        RECT 2520.870 2262.800 2902.070 2262.940 ;
        RECT 2520.870 2262.740 2521.190 2262.800 ;
        RECT 2901.750 2262.740 2902.070 2262.800 ;
      LAYER via ;
        RECT 2520.900 2262.740 2521.160 2263.000 ;
        RECT 2901.780 2262.740 2902.040 2263.000 ;
      LAYER met2 ;
        RECT 2901.770 2493.035 2902.050 2493.405 ;
        RECT 2901.840 2263.030 2901.980 2493.035 ;
        RECT 2520.900 2262.710 2521.160 2263.030 ;
        RECT 2901.780 2262.710 2902.040 2263.030 ;
        RECT 2520.960 2259.485 2521.100 2262.710 ;
        RECT 2520.890 2259.115 2521.170 2259.485 ;
      LAYER via2 ;
        RECT 2901.770 2493.080 2902.050 2493.360 ;
        RECT 2520.890 2259.160 2521.170 2259.440 ;
      LAYER met3 ;
        RECT 2901.745 2493.370 2902.075 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2901.745 2493.070 2924.800 2493.370 ;
        RECT 2901.745 2493.055 2902.075 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2506.000 2259.450 2510.000 2259.600 ;
        RECT 2520.865 2259.450 2521.195 2259.465 ;
        RECT 2506.000 2259.150 2521.195 2259.450 ;
        RECT 2506.000 2259.000 2510.000 2259.150 ;
        RECT 2520.865 2259.135 2521.195 2259.150 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2428.860 2525.330 2428.920 ;
        RECT 2901.290 2428.860 2901.610 2428.920 ;
        RECT 2525.010 2428.720 2901.610 2428.860 ;
        RECT 2525.010 2428.660 2525.330 2428.720 ;
        RECT 2901.290 2428.660 2901.610 2428.720 ;
      LAYER via ;
        RECT 2525.040 2428.660 2525.300 2428.920 ;
        RECT 2901.320 2428.660 2901.580 2428.920 ;
      LAYER met2 ;
        RECT 2901.310 2727.635 2901.590 2728.005 ;
        RECT 2901.380 2428.950 2901.520 2727.635 ;
        RECT 2525.040 2428.630 2525.300 2428.950 ;
        RECT 2901.320 2428.630 2901.580 2428.950 ;
        RECT 2525.100 2426.085 2525.240 2428.630 ;
        RECT 2525.030 2425.715 2525.310 2426.085 ;
      LAYER via2 ;
        RECT 2901.310 2727.680 2901.590 2727.960 ;
        RECT 2525.030 2425.760 2525.310 2426.040 ;
      LAYER met3 ;
        RECT 2901.285 2727.970 2901.615 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2901.285 2727.670 2924.800 2727.970 ;
        RECT 2901.285 2727.655 2901.615 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2506.000 2426.050 2510.000 2426.200 ;
        RECT 2525.005 2426.050 2525.335 2426.065 ;
        RECT 2506.000 2425.750 2525.335 2426.050 ;
        RECT 2506.000 2425.600 2510.000 2425.750 ;
        RECT 2525.005 2425.735 2525.335 2425.750 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2535.590 2960.280 2535.910 2960.340 ;
        RECT 2899.450 2960.280 2899.770 2960.340 ;
        RECT 2535.590 2960.140 2899.770 2960.280 ;
        RECT 2535.590 2960.080 2535.910 2960.140 ;
        RECT 2899.450 2960.080 2899.770 2960.140 ;
        RECT 2520.870 2592.740 2521.190 2592.800 ;
        RECT 2535.590 2592.740 2535.910 2592.800 ;
        RECT 2520.870 2592.600 2535.910 2592.740 ;
        RECT 2520.870 2592.540 2521.190 2592.600 ;
        RECT 2535.590 2592.540 2535.910 2592.600 ;
      LAYER via ;
        RECT 2535.620 2960.080 2535.880 2960.340 ;
        RECT 2899.480 2960.080 2899.740 2960.340 ;
        RECT 2520.900 2592.540 2521.160 2592.800 ;
        RECT 2535.620 2592.540 2535.880 2592.800 ;
      LAYER met2 ;
        RECT 2899.470 2962.235 2899.750 2962.605 ;
        RECT 2899.540 2960.370 2899.680 2962.235 ;
        RECT 2535.620 2960.050 2535.880 2960.370 ;
        RECT 2899.480 2960.050 2899.740 2960.370 ;
        RECT 2535.680 2592.830 2535.820 2960.050 ;
        RECT 2520.900 2592.685 2521.160 2592.830 ;
        RECT 2520.890 2592.315 2521.170 2592.685 ;
        RECT 2535.620 2592.510 2535.880 2592.830 ;
      LAYER via2 ;
        RECT 2899.470 2962.280 2899.750 2962.560 ;
        RECT 2520.890 2592.360 2521.170 2592.640 ;
      LAYER met3 ;
        RECT 2899.445 2962.570 2899.775 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2899.445 2962.270 2924.800 2962.570 ;
        RECT 2899.445 2962.255 2899.775 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2506.000 2592.650 2510.000 2592.800 ;
        RECT 2520.865 2592.650 2521.195 2592.665 ;
        RECT 2506.000 2592.350 2521.195 2592.650 ;
        RECT 2506.000 2592.200 2510.000 2592.350 ;
        RECT 2520.865 2592.335 2521.195 2592.350 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2760.020 2525.330 2760.080 ;
        RECT 2901.750 2760.020 2902.070 2760.080 ;
        RECT 2525.010 2759.880 2902.070 2760.020 ;
        RECT 2525.010 2759.820 2525.330 2759.880 ;
        RECT 2901.750 2759.820 2902.070 2759.880 ;
      LAYER via ;
        RECT 2525.040 2759.820 2525.300 2760.080 ;
        RECT 2901.780 2759.820 2902.040 2760.080 ;
      LAYER met2 ;
        RECT 2901.770 3196.835 2902.050 3197.205 ;
        RECT 2901.840 2760.110 2901.980 3196.835 ;
        RECT 2525.040 2759.790 2525.300 2760.110 ;
        RECT 2901.780 2759.790 2902.040 2760.110 ;
        RECT 2525.100 2759.285 2525.240 2759.790 ;
        RECT 2525.030 2758.915 2525.310 2759.285 ;
      LAYER via2 ;
        RECT 2901.770 3196.880 2902.050 3197.160 ;
        RECT 2525.030 2758.960 2525.310 2759.240 ;
      LAYER met3 ;
        RECT 2901.745 3197.170 2902.075 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.745 3196.870 2924.800 3197.170 ;
        RECT 2901.745 3196.855 2902.075 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2506.000 2759.250 2510.000 2759.400 ;
        RECT 2525.005 2759.250 2525.335 2759.265 ;
        RECT 2506.000 2758.950 2525.335 2759.250 ;
        RECT 2506.000 2758.800 2510.000 2758.950 ;
        RECT 2525.005 2758.935 2525.335 2758.950 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 2932.400 2523.490 2932.460 ;
        RECT 2901.290 2932.400 2901.610 2932.460 ;
        RECT 2523.170 2932.260 2901.610 2932.400 ;
        RECT 2523.170 2932.200 2523.490 2932.260 ;
        RECT 2901.290 2932.200 2901.610 2932.260 ;
      LAYER via ;
        RECT 2523.200 2932.200 2523.460 2932.460 ;
        RECT 2901.320 2932.200 2901.580 2932.460 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 2901.380 2932.490 2901.520 3431.435 ;
        RECT 2523.200 2932.170 2523.460 2932.490 ;
        RECT 2901.320 2932.170 2901.580 2932.490 ;
        RECT 2523.260 2925.885 2523.400 2932.170 ;
        RECT 2523.190 2925.515 2523.470 2925.885 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
        RECT 2523.190 2925.560 2523.470 2925.840 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2506.000 2925.850 2510.000 2926.000 ;
        RECT 2523.165 2925.850 2523.495 2925.865 ;
        RECT 2506.000 2925.550 2523.495 2925.850 ;
        RECT 2506.000 2925.400 2510.000 2925.550 ;
        RECT 2523.165 2925.535 2523.495 2925.550 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3415.555 ;
      LAYER mcon ;
        RECT 2713.685 3415.385 2713.855 3415.555 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2712.690 3470.620 2713.010 3470.680 ;
        RECT 2713.610 3470.620 2713.930 3470.680 ;
        RECT 2712.690 3470.480 2713.930 3470.620 ;
        RECT 2712.690 3470.420 2713.010 3470.480 ;
        RECT 2713.610 3470.420 2713.930 3470.480 ;
        RECT 2712.690 3463.820 2713.010 3463.880 ;
        RECT 2713.610 3463.820 2713.930 3463.880 ;
        RECT 2712.690 3463.680 2713.930 3463.820 ;
        RECT 2712.690 3463.620 2713.010 3463.680 ;
        RECT 2713.610 3463.620 2713.930 3463.680 ;
        RECT 2711.770 3415.540 2712.090 3415.600 ;
        RECT 2713.625 3415.540 2713.915 3415.585 ;
        RECT 2711.770 3415.400 2713.915 3415.540 ;
        RECT 2711.770 3415.340 2712.090 3415.400 ;
        RECT 2713.625 3415.355 2713.915 3415.400 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2392.530 3019.100 2392.850 3019.160 ;
        RECT 2712.230 3019.100 2712.550 3019.160 ;
        RECT 2392.530 3018.960 2712.550 3019.100 ;
        RECT 2392.530 3018.900 2392.850 3018.960 ;
        RECT 2712.230 3018.900 2712.550 3018.960 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2712.720 3470.420 2712.980 3470.680 ;
        RECT 2713.640 3470.420 2713.900 3470.680 ;
        RECT 2712.720 3463.620 2712.980 3463.880 ;
        RECT 2713.640 3463.620 2713.900 3463.880 ;
        RECT 2711.800 3415.340 2712.060 3415.600 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2392.560 3018.900 2392.820 3019.160 ;
        RECT 2712.260 3018.900 2712.520 3019.160 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3470.710 2713.840 3491.130 ;
        RECT 2712.720 3470.390 2712.980 3470.710 ;
        RECT 2713.640 3470.390 2713.900 3470.710 ;
        RECT 2712.780 3463.910 2712.920 3470.390 ;
        RECT 2712.720 3463.590 2712.980 3463.910 ;
        RECT 2713.640 3463.590 2713.900 3463.910 ;
        RECT 2713.700 3416.165 2713.840 3463.590 ;
        RECT 2711.790 3415.795 2712.070 3416.165 ;
        RECT 2713.630 3415.795 2713.910 3416.165 ;
        RECT 2711.860 3415.630 2712.000 3415.795 ;
        RECT 2711.800 3415.310 2712.060 3415.630 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3019.190 2712.460 3056.610 ;
        RECT 2392.560 3018.870 2392.820 3019.190 ;
        RECT 2712.260 3018.870 2712.520 3019.190 ;
        RECT 2392.620 3010.000 2392.760 3018.870 ;
        RECT 2392.620 3009.340 2392.970 3010.000 ;
        RECT 2392.690 3006.000 2392.970 3009.340 ;
      LAYER via2 ;
        RECT 2711.790 3415.840 2712.070 3416.120 ;
        RECT 2713.630 3415.840 2713.910 3416.120 ;
      LAYER met3 ;
        RECT 2711.765 3416.130 2712.095 3416.145 ;
        RECT 2713.605 3416.130 2713.935 3416.145 ;
        RECT 2711.765 3415.830 2713.935 3416.130 ;
        RECT 2711.765 3415.815 2712.095 3415.830 ;
        RECT 2713.605 3415.815 2713.935 3415.830 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.470 3464.160 2387.790 3464.220 ;
        RECT 2392.990 3464.160 2393.310 3464.220 ;
        RECT 2387.470 3464.020 2393.310 3464.160 ;
        RECT 2387.470 3463.960 2387.790 3464.020 ;
        RECT 2392.990 3463.960 2393.310 3464.020 ;
        RECT 2387.470 3367.600 2387.790 3367.660 ;
        RECT 2388.390 3367.600 2388.710 3367.660 ;
        RECT 2387.470 3367.460 2388.710 3367.600 ;
        RECT 2387.470 3367.400 2387.790 3367.460 ;
        RECT 2388.390 3367.400 2388.710 3367.460 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 2387.470 3077.580 2387.790 3077.640 ;
        RECT 2388.390 3077.580 2388.710 3077.640 ;
        RECT 2387.470 3077.440 2388.710 3077.580 ;
        RECT 2387.470 3077.380 2387.790 3077.440 ;
        RECT 2388.390 3077.380 2388.710 3077.440 ;
        RECT 2159.310 3019.100 2159.630 3019.160 ;
        RECT 2388.390 3019.100 2388.710 3019.160 ;
        RECT 2159.310 3018.960 2388.710 3019.100 ;
        RECT 2159.310 3018.900 2159.630 3018.960 ;
        RECT 2388.390 3018.900 2388.710 3018.960 ;
      LAYER via ;
        RECT 2387.500 3463.960 2387.760 3464.220 ;
        RECT 2393.020 3463.960 2393.280 3464.220 ;
        RECT 2387.500 3367.400 2387.760 3367.660 ;
        RECT 2388.420 3367.400 2388.680 3367.660 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 2387.500 3077.380 2387.760 3077.640 ;
        RECT 2388.420 3077.380 2388.680 3077.640 ;
        RECT 2159.340 3018.900 2159.600 3019.160 ;
        RECT 2388.420 3018.900 2388.680 3019.160 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3464.250 2393.220 3517.230 ;
        RECT 2387.500 3463.930 2387.760 3464.250 ;
        RECT 2393.020 3463.930 2393.280 3464.250 ;
        RECT 2387.560 3415.370 2387.700 3463.930 ;
        RECT 2387.560 3415.230 2388.620 3415.370 ;
        RECT 2388.480 3367.690 2388.620 3415.230 ;
        RECT 2387.500 3367.370 2387.760 3367.690 ;
        RECT 2388.420 3367.370 2388.680 3367.690 ;
        RECT 2387.560 3318.810 2387.700 3367.370 ;
        RECT 2387.560 3318.670 2388.620 3318.810 ;
        RECT 2388.480 3270.790 2388.620 3318.670 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 3019.190 2388.620 3028.990 ;
        RECT 2159.340 3018.870 2159.600 3019.190 ;
        RECT 2388.420 3018.870 2388.680 3019.190 ;
        RECT 2159.400 3010.000 2159.540 3018.870 ;
        RECT 2159.400 3009.340 2159.750 3010.000 ;
        RECT 2159.470 3006.000 2159.750 3009.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2063.245 3416.065 2063.415 3463.835 ;
        RECT 2065.085 3332.765 2065.255 3415.555 ;
      LAYER mcon ;
        RECT 2063.245 3463.665 2063.415 3463.835 ;
        RECT 2065.085 3415.385 2065.255 3415.555 ;
      LAYER met1 ;
        RECT 2065.010 3491.360 2065.330 3491.420 ;
        RECT 2068.690 3491.360 2069.010 3491.420 ;
        RECT 2065.010 3491.220 2069.010 3491.360 ;
        RECT 2065.010 3491.160 2065.330 3491.220 ;
        RECT 2068.690 3491.160 2069.010 3491.220 ;
        RECT 2064.090 3470.620 2064.410 3470.680 ;
        RECT 2065.010 3470.620 2065.330 3470.680 ;
        RECT 2064.090 3470.480 2065.330 3470.620 ;
        RECT 2064.090 3470.420 2064.410 3470.480 ;
        RECT 2065.010 3470.420 2065.330 3470.480 ;
        RECT 2063.185 3463.820 2063.475 3463.865 ;
        RECT 2064.090 3463.820 2064.410 3463.880 ;
        RECT 2063.185 3463.680 2064.410 3463.820 ;
        RECT 2063.185 3463.635 2063.475 3463.680 ;
        RECT 2064.090 3463.620 2064.410 3463.680 ;
        RECT 2063.170 3416.220 2063.490 3416.280 ;
        RECT 2063.170 3416.080 2063.685 3416.220 ;
        RECT 2063.170 3416.020 2063.490 3416.080 ;
        RECT 2063.170 3415.540 2063.490 3415.600 ;
        RECT 2065.025 3415.540 2065.315 3415.585 ;
        RECT 2063.170 3415.400 2065.315 3415.540 ;
        RECT 2063.170 3415.340 2063.490 3415.400 ;
        RECT 2065.025 3415.355 2065.315 3415.400 ;
        RECT 2065.025 3332.920 2065.315 3332.965 ;
        RECT 2065.470 3332.920 2065.790 3332.980 ;
        RECT 2065.025 3332.780 2065.790 3332.920 ;
        RECT 2065.025 3332.735 2065.315 3332.780 ;
        RECT 2065.470 3332.720 2065.790 3332.780 ;
        RECT 2064.090 3236.360 2064.410 3236.420 ;
        RECT 2064.550 3236.360 2064.870 3236.420 ;
        RECT 2064.090 3236.220 2064.870 3236.360 ;
        RECT 2064.090 3236.160 2064.410 3236.220 ;
        RECT 2064.550 3236.160 2064.870 3236.220 ;
        RECT 2064.090 3202.020 2064.410 3202.080 ;
        RECT 2064.550 3202.020 2064.870 3202.080 ;
        RECT 2064.090 3201.880 2064.870 3202.020 ;
        RECT 2064.090 3201.820 2064.410 3201.880 ;
        RECT 2064.550 3201.820 2064.870 3201.880 ;
        RECT 2063.630 3153.400 2063.950 3153.460 ;
        RECT 2064.550 3153.400 2064.870 3153.460 ;
        RECT 2063.630 3153.260 2064.870 3153.400 ;
        RECT 2063.630 3153.200 2063.950 3153.260 ;
        RECT 2064.550 3153.200 2064.870 3153.260 ;
        RECT 2063.630 3056.840 2063.950 3056.900 ;
        RECT 2064.550 3056.840 2064.870 3056.900 ;
        RECT 2063.630 3056.700 2064.870 3056.840 ;
        RECT 2063.630 3056.640 2063.950 3056.700 ;
        RECT 2064.550 3056.640 2064.870 3056.700 ;
        RECT 1926.090 3019.440 1926.410 3019.500 ;
        RECT 2063.630 3019.440 2063.950 3019.500 ;
        RECT 1926.090 3019.300 2063.950 3019.440 ;
        RECT 1926.090 3019.240 1926.410 3019.300 ;
        RECT 2063.630 3019.240 2063.950 3019.300 ;
      LAYER via ;
        RECT 2065.040 3491.160 2065.300 3491.420 ;
        RECT 2068.720 3491.160 2068.980 3491.420 ;
        RECT 2064.120 3470.420 2064.380 3470.680 ;
        RECT 2065.040 3470.420 2065.300 3470.680 ;
        RECT 2064.120 3463.620 2064.380 3463.880 ;
        RECT 2063.200 3416.020 2063.460 3416.280 ;
        RECT 2063.200 3415.340 2063.460 3415.600 ;
        RECT 2065.500 3332.720 2065.760 3332.980 ;
        RECT 2064.120 3236.160 2064.380 3236.420 ;
        RECT 2064.580 3236.160 2064.840 3236.420 ;
        RECT 2064.120 3201.820 2064.380 3202.080 ;
        RECT 2064.580 3201.820 2064.840 3202.080 ;
        RECT 2063.660 3153.200 2063.920 3153.460 ;
        RECT 2064.580 3153.200 2064.840 3153.460 ;
        RECT 2063.660 3056.640 2063.920 3056.900 ;
        RECT 2064.580 3056.640 2064.840 3056.900 ;
        RECT 1926.120 3019.240 1926.380 3019.500 ;
        RECT 2063.660 3019.240 2063.920 3019.500 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3470.710 2065.240 3491.130 ;
        RECT 2064.120 3470.390 2064.380 3470.710 ;
        RECT 2065.040 3470.390 2065.300 3470.710 ;
        RECT 2064.180 3463.910 2064.320 3470.390 ;
        RECT 2064.120 3463.590 2064.380 3463.910 ;
        RECT 2063.200 3415.990 2063.460 3416.310 ;
        RECT 2063.260 3415.630 2063.400 3415.990 ;
        RECT 2063.200 3415.310 2063.460 3415.630 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3019.530 2063.860 3056.610 ;
        RECT 1926.120 3019.210 1926.380 3019.530 ;
        RECT 2063.660 3019.210 2063.920 3019.530 ;
        RECT 1926.180 3010.000 1926.320 3019.210 ;
        RECT 1926.180 3009.340 1926.530 3010.000 ;
        RECT 1926.250 3006.000 1926.530 3009.340 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.870 3464.160 1739.190 3464.220 ;
        RECT 1744.390 3464.160 1744.710 3464.220 ;
        RECT 1738.870 3464.020 1744.710 3464.160 ;
        RECT 1738.870 3463.960 1739.190 3464.020 ;
        RECT 1744.390 3463.960 1744.710 3464.020 ;
        RECT 1738.870 3367.600 1739.190 3367.660 ;
        RECT 1739.790 3367.600 1740.110 3367.660 ;
        RECT 1738.870 3367.460 1740.110 3367.600 ;
        RECT 1738.870 3367.400 1739.190 3367.460 ;
        RECT 1739.790 3367.400 1740.110 3367.460 ;
        RECT 1738.870 3270.700 1739.190 3270.760 ;
        RECT 1739.790 3270.700 1740.110 3270.760 ;
        RECT 1738.870 3270.560 1740.110 3270.700 ;
        RECT 1738.870 3270.500 1739.190 3270.560 ;
        RECT 1739.790 3270.500 1740.110 3270.560 ;
        RECT 1738.870 3174.140 1739.190 3174.200 ;
        RECT 1739.790 3174.140 1740.110 3174.200 ;
        RECT 1738.870 3174.000 1740.110 3174.140 ;
        RECT 1738.870 3173.940 1739.190 3174.000 ;
        RECT 1739.790 3173.940 1740.110 3174.000 ;
        RECT 1738.870 3077.580 1739.190 3077.640 ;
        RECT 1739.790 3077.580 1740.110 3077.640 ;
        RECT 1738.870 3077.440 1740.110 3077.580 ;
        RECT 1738.870 3077.380 1739.190 3077.440 ;
        RECT 1739.790 3077.380 1740.110 3077.440 ;
        RECT 1692.870 3018.760 1693.190 3018.820 ;
        RECT 1739.790 3018.760 1740.110 3018.820 ;
        RECT 1692.870 3018.620 1740.110 3018.760 ;
        RECT 1692.870 3018.560 1693.190 3018.620 ;
        RECT 1739.790 3018.560 1740.110 3018.620 ;
      LAYER via ;
        RECT 1738.900 3463.960 1739.160 3464.220 ;
        RECT 1744.420 3463.960 1744.680 3464.220 ;
        RECT 1738.900 3367.400 1739.160 3367.660 ;
        RECT 1739.820 3367.400 1740.080 3367.660 ;
        RECT 1738.900 3270.500 1739.160 3270.760 ;
        RECT 1739.820 3270.500 1740.080 3270.760 ;
        RECT 1738.900 3173.940 1739.160 3174.200 ;
        RECT 1739.820 3173.940 1740.080 3174.200 ;
        RECT 1738.900 3077.380 1739.160 3077.640 ;
        RECT 1739.820 3077.380 1740.080 3077.640 ;
        RECT 1692.900 3018.560 1693.160 3018.820 ;
        RECT 1739.820 3018.560 1740.080 3018.820 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3517.370 1744.160 3517.600 ;
        RECT 1744.020 3517.230 1744.620 3517.370 ;
        RECT 1744.480 3464.250 1744.620 3517.230 ;
        RECT 1738.900 3463.930 1739.160 3464.250 ;
        RECT 1744.420 3463.930 1744.680 3464.250 ;
        RECT 1738.960 3415.370 1739.100 3463.930 ;
        RECT 1738.960 3415.230 1740.020 3415.370 ;
        RECT 1739.880 3367.690 1740.020 3415.230 ;
        RECT 1738.900 3367.370 1739.160 3367.690 ;
        RECT 1739.820 3367.370 1740.080 3367.690 ;
        RECT 1738.960 3318.810 1739.100 3367.370 ;
        RECT 1738.960 3318.670 1740.020 3318.810 ;
        RECT 1739.880 3270.790 1740.020 3318.670 ;
        RECT 1738.900 3270.470 1739.160 3270.790 ;
        RECT 1739.820 3270.470 1740.080 3270.790 ;
        RECT 1738.960 3222.250 1739.100 3270.470 ;
        RECT 1738.960 3222.110 1740.020 3222.250 ;
        RECT 1739.880 3174.230 1740.020 3222.110 ;
        RECT 1738.900 3173.910 1739.160 3174.230 ;
        RECT 1739.820 3173.910 1740.080 3174.230 ;
        RECT 1738.960 3125.690 1739.100 3173.910 ;
        RECT 1738.960 3125.550 1740.020 3125.690 ;
        RECT 1739.880 3077.670 1740.020 3125.550 ;
        RECT 1738.900 3077.350 1739.160 3077.670 ;
        RECT 1739.820 3077.350 1740.080 3077.670 ;
        RECT 1738.960 3029.130 1739.100 3077.350 ;
        RECT 1738.960 3028.990 1740.020 3029.130 ;
        RECT 1739.880 3018.850 1740.020 3028.990 ;
        RECT 1692.900 3018.530 1693.160 3018.850 ;
        RECT 1739.820 3018.530 1740.080 3018.850 ;
        RECT 1692.960 3010.000 1693.100 3018.530 ;
        RECT 1692.960 3009.340 1693.310 3010.000 ;
        RECT 1693.030 3006.000 1693.310 3009.340 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3270.700 1420.410 3270.760 ;
        RECT 1421.010 3270.700 1421.330 3270.760 ;
        RECT 1420.090 3270.560 1421.330 3270.700 ;
        RECT 1420.090 3270.500 1420.410 3270.560 ;
        RECT 1421.010 3270.500 1421.330 3270.560 ;
        RECT 1420.090 3174.140 1420.410 3174.200 ;
        RECT 1421.010 3174.140 1421.330 3174.200 ;
        RECT 1420.090 3174.000 1421.330 3174.140 ;
        RECT 1420.090 3173.940 1420.410 3174.000 ;
        RECT 1421.010 3173.940 1421.330 3174.000 ;
        RECT 1420.090 3077.580 1420.410 3077.640 ;
        RECT 1421.010 3077.580 1421.330 3077.640 ;
        RECT 1420.090 3077.440 1421.330 3077.580 ;
        RECT 1420.090 3077.380 1420.410 3077.440 ;
        RECT 1421.010 3077.380 1421.330 3077.440 ;
        RECT 1420.090 3018.760 1420.410 3018.820 ;
        RECT 1459.190 3018.760 1459.510 3018.820 ;
        RECT 1420.090 3018.620 1459.510 3018.760 ;
        RECT 1420.090 3018.560 1420.410 3018.620 ;
        RECT 1459.190 3018.560 1459.510 3018.620 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3270.500 1420.380 3270.760 ;
        RECT 1421.040 3270.500 1421.300 3270.760 ;
        RECT 1420.120 3173.940 1420.380 3174.200 ;
        RECT 1421.040 3173.940 1421.300 3174.200 ;
        RECT 1420.120 3077.380 1420.380 3077.640 ;
        RECT 1421.040 3077.380 1421.300 3077.640 ;
        RECT 1420.120 3018.560 1420.380 3018.820 ;
        RECT 1459.220 3018.560 1459.480 3018.820 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3222.250 1421.240 3270.470 ;
        RECT 1420.180 3222.110 1421.240 3222.250 ;
        RECT 1420.180 3174.230 1420.320 3222.110 ;
        RECT 1420.120 3173.910 1420.380 3174.230 ;
        RECT 1421.040 3173.910 1421.300 3174.230 ;
        RECT 1421.100 3125.690 1421.240 3173.910 ;
        RECT 1420.180 3125.550 1421.240 3125.690 ;
        RECT 1420.180 3077.670 1420.320 3125.550 ;
        RECT 1420.120 3077.350 1420.380 3077.670 ;
        RECT 1421.040 3077.350 1421.300 3077.670 ;
        RECT 1421.100 3029.130 1421.240 3077.350 ;
        RECT 1420.180 3028.990 1421.240 3029.130 ;
        RECT 1420.180 3018.850 1420.320 3028.990 ;
        RECT 1420.120 3018.530 1420.380 3018.850 ;
        RECT 1459.220 3018.530 1459.480 3018.850 ;
        RECT 1459.280 3010.000 1459.420 3018.530 ;
        RECT 1459.280 3009.340 1459.630 3010.000 ;
        RECT 1459.350 3006.000 1459.630 3009.340 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 386.140 2523.490 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2523.170 386.000 2901.150 386.140 ;
        RECT 2523.170 385.940 2523.490 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2523.200 385.940 2523.460 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2523.190 759.035 2523.470 759.405 ;
        RECT 2523.260 386.230 2523.400 759.035 ;
        RECT 2523.200 385.910 2523.460 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2523.190 759.080 2523.470 759.360 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2506.000 759.370 2510.000 759.520 ;
        RECT 2523.165 759.370 2523.495 759.385 ;
        RECT 2506.000 759.070 2523.495 759.370 ;
        RECT 2506.000 758.920 2510.000 759.070 ;
        RECT 2523.165 759.055 2523.495 759.070 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1095.405 3139.645 1095.575 3187.755 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1095.405 3187.585 1095.575 3187.755 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.135 3187.600 1095.650 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.345 3139.800 1095.635 3139.845 ;
        RECT 1096.710 3139.800 1097.030 3139.860 ;
        RECT 1095.345 3139.660 1097.030 3139.800 ;
        RECT 1095.345 3139.615 1095.635 3139.660 ;
        RECT 1096.710 3139.600 1097.030 3139.660 ;
        RECT 1096.710 3018.760 1097.030 3018.820 ;
        RECT 1225.970 3018.760 1226.290 3018.820 ;
        RECT 1096.710 3018.620 1226.290 3018.760 ;
        RECT 1096.710 3018.560 1097.030 3018.620 ;
        RECT 1225.970 3018.560 1226.290 3018.620 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1096.740 3139.600 1097.000 3139.860 ;
        RECT 1096.740 3018.560 1097.000 3018.820 ;
        RECT 1226.000 3018.560 1226.260 3018.820 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1096.740 3139.570 1097.000 3139.890 ;
        RECT 1096.800 3018.850 1096.940 3139.570 ;
        RECT 1096.740 3018.530 1097.000 3018.850 ;
        RECT 1226.000 3018.530 1226.260 3018.850 ;
        RECT 1226.060 3010.000 1226.200 3018.530 ;
        RECT 1226.060 3009.340 1226.410 3010.000 ;
        RECT 1226.130 3006.000 1226.410 3009.340 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 3019.440 771.810 3019.500 ;
        RECT 992.750 3019.440 993.070 3019.500 ;
        RECT 771.490 3019.300 993.070 3019.440 ;
        RECT 771.490 3019.240 771.810 3019.300 ;
        RECT 992.750 3019.240 993.070 3019.300 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 3019.240 771.780 3019.500 ;
        RECT 992.780 3019.240 993.040 3019.500 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 3019.530 771.720 3028.990 ;
        RECT 771.520 3019.210 771.780 3019.530 ;
        RECT 992.780 3019.210 993.040 3019.530 ;
        RECT 992.840 3010.000 992.980 3019.210 ;
        RECT 992.840 3009.340 993.190 3010.000 ;
        RECT 992.910 3006.000 993.190 3009.340 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 3020.120 448.430 3020.180 ;
        RECT 759.530 3020.120 759.850 3020.180 ;
        RECT 448.110 3019.980 759.850 3020.120 ;
        RECT 448.110 3019.920 448.430 3019.980 ;
        RECT 759.530 3019.920 759.850 3019.980 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 3019.920 448.400 3020.180 ;
        RECT 759.560 3019.920 759.820 3020.180 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 3020.210 448.340 3498.270 ;
        RECT 448.140 3019.890 448.400 3020.210 ;
        RECT 759.560 3019.890 759.820 3020.210 ;
        RECT 759.620 3010.000 759.760 3019.890 ;
        RECT 759.620 3009.340 759.970 3010.000 ;
        RECT 759.690 3006.000 759.970 3009.340 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 3019.100 124.130 3019.160 ;
        RECT 526.310 3019.100 526.630 3019.160 ;
        RECT 123.810 3018.960 526.630 3019.100 ;
        RECT 123.810 3018.900 124.130 3018.960 ;
        RECT 526.310 3018.900 526.630 3018.960 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 3018.900 124.100 3019.160 ;
        RECT 526.340 3018.900 526.600 3019.160 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 3019.190 124.040 3498.270 ;
        RECT 123.840 3018.870 124.100 3019.190 ;
        RECT 526.340 3018.870 526.600 3019.190 ;
        RECT 526.400 3010.000 526.540 3018.870 ;
        RECT 526.400 3009.340 526.750 3010.000 ;
        RECT 526.470 3006.000 526.750 3009.340 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2925.600 17.410 2925.660 ;
        RECT 393.370 2925.600 393.690 2925.660 ;
        RECT 17.090 2925.460 393.690 2925.600 ;
        RECT 17.090 2925.400 17.410 2925.460 ;
        RECT 393.370 2925.400 393.690 2925.460 ;
      LAYER via ;
        RECT 17.120 2925.400 17.380 2925.660 ;
        RECT 393.400 2925.400 393.660 2925.660 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 2925.690 17.320 3339.635 ;
        RECT 17.120 2925.370 17.380 2925.690 ;
        RECT 393.400 2925.370 393.660 2925.690 ;
        RECT 393.460 2919.765 393.600 2925.370 ;
        RECT 393.390 2919.395 393.670 2919.765 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 393.390 2919.440 393.670 2919.720 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 393.365 2919.730 393.695 2919.745 ;
        RECT 410.000 2919.730 414.000 2919.880 ;
        RECT 393.365 2919.430 414.000 2919.730 ;
        RECT 393.365 2919.415 393.695 2919.430 ;
        RECT 410.000 2919.280 414.000 2919.430 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2746.080 17.870 2746.140 ;
        RECT 393.370 2746.080 393.690 2746.140 ;
        RECT 17.550 2745.940 393.690 2746.080 ;
        RECT 17.550 2745.880 17.870 2745.940 ;
        RECT 393.370 2745.880 393.690 2745.940 ;
      LAYER via ;
        RECT 17.580 2745.880 17.840 2746.140 ;
        RECT 393.400 2745.880 393.660 2746.140 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 2746.170 17.780 3051.995 ;
        RECT 17.580 2745.850 17.840 2746.170 ;
        RECT 393.400 2745.850 393.660 2746.170 ;
        RECT 393.460 2741.605 393.600 2745.850 ;
        RECT 393.390 2741.235 393.670 2741.605 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 393.390 2741.280 393.670 2741.560 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 393.365 2741.570 393.695 2741.585 ;
        RECT 410.000 2741.570 414.000 2741.720 ;
        RECT 393.365 2741.270 414.000 2741.570 ;
        RECT 393.365 2741.255 393.695 2741.270 ;
        RECT 410.000 2741.120 414.000 2741.270 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2566.560 17.410 2566.620 ;
        RECT 393.370 2566.560 393.690 2566.620 ;
        RECT 17.090 2566.420 393.690 2566.560 ;
        RECT 17.090 2566.360 17.410 2566.420 ;
        RECT 393.370 2566.360 393.690 2566.420 ;
      LAYER via ;
        RECT 17.120 2566.360 17.380 2566.620 ;
        RECT 393.400 2566.360 393.660 2566.620 ;
      LAYER met2 ;
        RECT 17.110 2765.035 17.390 2765.405 ;
        RECT 17.180 2566.650 17.320 2765.035 ;
        RECT 17.120 2566.330 17.380 2566.650 ;
        RECT 393.400 2566.330 393.660 2566.650 ;
        RECT 393.460 2562.765 393.600 2566.330 ;
        RECT 393.390 2562.395 393.670 2562.765 ;
      LAYER via2 ;
        RECT 17.110 2765.080 17.390 2765.360 ;
        RECT 393.390 2562.440 393.670 2562.720 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.085 2765.370 17.415 2765.385 ;
        RECT -4.800 2765.070 17.415 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.085 2765.055 17.415 2765.070 ;
        RECT 393.365 2562.730 393.695 2562.745 ;
        RECT 410.000 2562.730 414.000 2562.880 ;
        RECT 393.365 2562.430 414.000 2562.730 ;
        RECT 393.365 2562.415 393.695 2562.430 ;
        RECT 410.000 2562.280 414.000 2562.430 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2387.380 17.870 2387.440 ;
        RECT 393.370 2387.380 393.690 2387.440 ;
        RECT 17.550 2387.240 393.690 2387.380 ;
        RECT 17.550 2387.180 17.870 2387.240 ;
        RECT 393.370 2387.180 393.690 2387.240 ;
      LAYER via ;
        RECT 17.580 2387.180 17.840 2387.440 ;
        RECT 393.400 2387.180 393.660 2387.440 ;
      LAYER met2 ;
        RECT 17.570 2477.395 17.850 2477.765 ;
        RECT 17.640 2387.470 17.780 2477.395 ;
        RECT 17.580 2387.150 17.840 2387.470 ;
        RECT 393.400 2387.150 393.660 2387.470 ;
        RECT 393.460 2384.605 393.600 2387.150 ;
        RECT 393.390 2384.235 393.670 2384.605 ;
      LAYER via2 ;
        RECT 17.570 2477.440 17.850 2477.720 ;
        RECT 393.390 2384.280 393.670 2384.560 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.545 2477.730 17.875 2477.745 ;
        RECT -4.800 2477.430 17.875 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.545 2477.415 17.875 2477.430 ;
        RECT 393.365 2384.570 393.695 2384.585 ;
        RECT 410.000 2384.570 414.000 2384.720 ;
        RECT 393.365 2384.270 414.000 2384.570 ;
        RECT 393.365 2384.255 393.695 2384.270 ;
        RECT 410.000 2384.120 414.000 2384.270 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2194.260 16.030 2194.320 ;
        RECT 393.370 2194.260 393.690 2194.320 ;
        RECT 15.710 2194.120 393.690 2194.260 ;
        RECT 15.710 2194.060 16.030 2194.120 ;
        RECT 393.370 2194.060 393.690 2194.120 ;
      LAYER via ;
        RECT 15.740 2194.060 16.000 2194.320 ;
        RECT 393.400 2194.060 393.660 2194.320 ;
      LAYER met2 ;
        RECT 393.390 2205.395 393.670 2205.765 ;
        RECT 393.460 2194.350 393.600 2205.395 ;
        RECT 15.740 2194.030 16.000 2194.350 ;
        RECT 393.400 2194.030 393.660 2194.350 ;
        RECT 15.800 2190.125 15.940 2194.030 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 393.390 2205.440 393.670 2205.720 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT 393.365 2205.730 393.695 2205.745 ;
        RECT 410.000 2205.730 414.000 2205.880 ;
        RECT 393.365 2205.430 414.000 2205.730 ;
        RECT 393.365 2205.415 393.695 2205.430 ;
        RECT 410.000 2205.280 414.000 2205.430 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 397.050 1904.240 397.370 1904.300 ;
        RECT 16.170 1904.100 397.370 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 397.050 1904.040 397.370 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 397.080 1904.040 397.340 1904.300 ;
      LAYER met2 ;
        RECT 397.070 2027.235 397.350 2027.605 ;
        RECT 397.140 1904.330 397.280 2027.235 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 397.080 1904.010 397.340 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 397.070 2027.280 397.350 2027.560 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 397.045 2027.570 397.375 2027.585 ;
        RECT 410.000 2027.570 414.000 2027.720 ;
        RECT 397.045 2027.270 414.000 2027.570 ;
        RECT 397.045 2027.255 397.375 2027.270 ;
        RECT 410.000 2027.120 414.000 2027.270 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2524.090 620.740 2524.410 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2524.090 620.600 2901.150 620.740 ;
        RECT 2524.090 620.540 2524.410 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2524.120 620.540 2524.380 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2524.110 925.635 2524.390 926.005 ;
        RECT 2524.180 620.830 2524.320 925.635 ;
        RECT 2524.120 620.510 2524.380 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2524.110 925.680 2524.390 925.960 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2506.000 925.970 2510.000 926.120 ;
        RECT 2524.085 925.970 2524.415 925.985 ;
        RECT 2506.000 925.670 2524.415 925.970 ;
        RECT 2506.000 925.520 2510.000 925.670 ;
        RECT 2524.085 925.655 2524.415 925.670 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 397.510 1621.360 397.830 1621.420 ;
        RECT 16.170 1621.220 397.830 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 397.510 1621.160 397.830 1621.220 ;
      LAYER via ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 397.540 1621.160 397.800 1621.420 ;
      LAYER met2 ;
        RECT 397.530 1848.395 397.810 1848.765 ;
        RECT 397.600 1621.450 397.740 1848.395 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 397.540 1621.130 397.800 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 397.530 1848.440 397.810 1848.720 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 397.505 1848.730 397.835 1848.745 ;
        RECT 410.000 1848.730 414.000 1848.880 ;
        RECT 397.505 1848.430 414.000 1848.730 ;
        RECT 397.505 1848.415 397.835 1848.430 ;
        RECT 410.000 1848.280 414.000 1848.430 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 398.430 1400.700 398.750 1400.760 ;
        RECT 17.090 1400.560 398.750 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 398.430 1400.500 398.750 1400.560 ;
      LAYER via ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 398.460 1400.500 398.720 1400.760 ;
      LAYER met2 ;
        RECT 398.450 1669.555 398.730 1669.925 ;
        RECT 398.520 1400.790 398.660 1669.555 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 398.460 1400.470 398.720 1400.790 ;
      LAYER via2 ;
        RECT 398.450 1669.600 398.730 1669.880 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 398.425 1669.890 398.755 1669.905 ;
        RECT 410.000 1669.890 414.000 1670.040 ;
        RECT 398.425 1669.590 414.000 1669.890 ;
        RECT 398.425 1669.575 398.755 1669.590 ;
        RECT 410.000 1669.440 414.000 1669.590 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 397.050 1186.840 397.370 1186.900 ;
        RECT 17.090 1186.700 397.370 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 397.050 1186.640 397.370 1186.700 ;
      LAYER via ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 397.080 1186.640 397.340 1186.900 ;
      LAYER met2 ;
        RECT 397.070 1491.395 397.350 1491.765 ;
        RECT 397.140 1186.930 397.280 1491.395 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 397.080 1186.610 397.340 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 397.070 1491.440 397.350 1491.720 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 397.045 1491.730 397.375 1491.745 ;
        RECT 410.000 1491.730 414.000 1491.880 ;
        RECT 397.045 1491.430 414.000 1491.730 ;
        RECT 397.045 1491.415 397.375 1491.430 ;
        RECT 410.000 1491.280 414.000 1491.430 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 397.970 972.640 398.290 972.700 ;
        RECT 15.710 972.500 398.290 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 397.970 972.440 398.290 972.500 ;
      LAYER via ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 398.000 972.440 398.260 972.700 ;
      LAYER met2 ;
        RECT 397.990 1312.555 398.270 1312.925 ;
        RECT 398.060 972.730 398.200 1312.555 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 398.000 972.410 398.260 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 397.990 1312.600 398.270 1312.880 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 397.965 1312.890 398.295 1312.905 ;
        RECT 410.000 1312.890 414.000 1313.040 ;
        RECT 397.965 1312.590 414.000 1312.890 ;
        RECT 397.965 1312.575 398.295 1312.590 ;
        RECT 410.000 1312.440 414.000 1312.590 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 397.050 758.780 397.370 758.840 ;
        RECT 15.710 758.640 397.370 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 397.050 758.580 397.370 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 397.080 758.580 397.340 758.840 ;
      LAYER met2 ;
        RECT 397.070 1134.395 397.350 1134.765 ;
        RECT 397.140 758.870 397.280 1134.395 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 397.080 758.550 397.340 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 397.070 1134.440 397.350 1134.720 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 397.045 1134.730 397.375 1134.745 ;
        RECT 410.000 1134.730 414.000 1134.880 ;
        RECT 397.045 1134.430 414.000 1134.730 ;
        RECT 397.045 1134.415 397.375 1134.430 ;
        RECT 410.000 1134.280 414.000 1134.430 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 398.890 544.920 399.210 544.980 ;
        RECT 16.170 544.780 399.210 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 398.890 544.720 399.210 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 398.920 544.720 399.180 544.980 ;
      LAYER met2 ;
        RECT 398.910 955.555 399.190 955.925 ;
        RECT 398.980 545.010 399.120 955.555 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 398.920 544.690 399.180 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 398.910 955.600 399.190 955.880 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 398.885 955.890 399.215 955.905 ;
        RECT 410.000 955.890 414.000 956.040 ;
        RECT 398.885 955.590 414.000 955.890 ;
        RECT 398.885 955.575 399.215 955.590 ;
        RECT 410.000 955.440 414.000 955.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 397.970 324.260 398.290 324.320 ;
        RECT 16.630 324.120 398.290 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 397.970 324.060 398.290 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 398.000 324.060 398.260 324.320 ;
      LAYER met2 ;
        RECT 397.990 777.395 398.270 777.765 ;
        RECT 398.060 324.350 398.200 777.395 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 398.000 324.030 398.260 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 397.990 777.440 398.270 777.720 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 397.965 777.730 398.295 777.745 ;
        RECT 410.000 777.730 414.000 777.880 ;
        RECT 397.965 777.430 414.000 777.730 ;
        RECT 397.965 777.415 398.295 777.430 ;
        RECT 410.000 777.280 414.000 777.430 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 397.050 110.400 397.370 110.460 ;
        RECT 15.710 110.260 397.370 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 397.050 110.200 397.370 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 397.080 110.200 397.340 110.460 ;
      LAYER met2 ;
        RECT 397.070 598.555 397.350 598.925 ;
        RECT 397.140 110.490 397.280 598.555 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 397.080 110.170 397.340 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 397.070 598.600 397.350 598.880 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 397.045 598.890 397.375 598.905 ;
        RECT 410.000 598.890 414.000 599.040 ;
        RECT 397.045 598.590 414.000 598.890 ;
        RECT 397.045 598.575 397.375 598.590 ;
        RECT 410.000 598.440 414.000 598.590 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 855.340 2523.490 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2523.170 855.200 2901.150 855.340 ;
        RECT 2523.170 855.140 2523.490 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2523.200 855.140 2523.460 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2523.190 1092.235 2523.470 1092.605 ;
        RECT 2523.260 855.430 2523.400 1092.235 ;
        RECT 2523.200 855.110 2523.460 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2523.190 1092.280 2523.470 1092.560 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2506.000 1092.570 2510.000 1092.720 ;
        RECT 2523.165 1092.570 2523.495 1092.585 ;
        RECT 2506.000 1092.270 2523.495 1092.570 ;
        RECT 2506.000 1092.120 2510.000 1092.270 ;
        RECT 2523.165 1092.255 2523.495 1092.270 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.630 1089.940 2523.950 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2523.630 1089.800 2901.150 1089.940 ;
        RECT 2523.630 1089.740 2523.950 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2523.660 1089.740 2523.920 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2523.650 1258.835 2523.930 1259.205 ;
        RECT 2523.720 1090.030 2523.860 1258.835 ;
        RECT 2523.660 1089.710 2523.920 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2523.650 1258.880 2523.930 1259.160 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2506.000 1259.170 2510.000 1259.320 ;
        RECT 2523.625 1259.170 2523.955 1259.185 ;
        RECT 2506.000 1258.870 2523.955 1259.170 ;
        RECT 2506.000 1258.720 2510.000 1258.870 ;
        RECT 2523.625 1258.855 2523.955 1258.870 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 1324.540 2522.570 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2522.250 1324.400 2901.150 1324.540 ;
        RECT 2522.250 1324.340 2522.570 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2522.280 1324.340 2522.540 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2522.270 1426.115 2522.550 1426.485 ;
        RECT 2522.340 1324.630 2522.480 1426.115 ;
        RECT 2522.280 1324.310 2522.540 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2522.270 1426.160 2522.550 1426.440 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2506.000 1426.450 2510.000 1426.600 ;
        RECT 2522.245 1426.450 2522.575 1426.465 ;
        RECT 2506.000 1426.150 2522.575 1426.450 ;
        RECT 2506.000 1426.000 2510.000 1426.150 ;
        RECT 2522.245 1426.135 2522.575 1426.150 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.030 1559.140 2519.350 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2519.030 1559.000 2901.150 1559.140 ;
        RECT 2519.030 1558.940 2519.350 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2519.060 1558.940 2519.320 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2519.050 1592.715 2519.330 1593.085 ;
        RECT 2519.120 1559.230 2519.260 1592.715 ;
        RECT 2519.060 1558.910 2519.320 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2519.050 1592.760 2519.330 1593.040 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2506.000 1593.050 2510.000 1593.200 ;
        RECT 2519.025 1593.050 2519.355 1593.065 ;
        RECT 2506.000 1592.750 2519.355 1593.050 ;
        RECT 2506.000 1592.600 2510.000 1592.750 ;
        RECT 2519.025 1592.735 2519.355 1592.750 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 1766.200 2523.490 1766.260 ;
        RECT 2901.290 1766.200 2901.610 1766.260 ;
        RECT 2523.170 1766.060 2901.610 1766.200 ;
        RECT 2523.170 1766.000 2523.490 1766.060 ;
        RECT 2901.290 1766.000 2901.610 1766.060 ;
      LAYER via ;
        RECT 2523.200 1766.000 2523.460 1766.260 ;
        RECT 2901.320 1766.000 2901.580 1766.260 ;
      LAYER met2 ;
        RECT 2901.310 1789.235 2901.590 1789.605 ;
        RECT 2901.380 1766.290 2901.520 1789.235 ;
        RECT 2523.200 1765.970 2523.460 1766.290 ;
        RECT 2901.320 1765.970 2901.580 1766.290 ;
        RECT 2523.260 1759.685 2523.400 1765.970 ;
        RECT 2523.190 1759.315 2523.470 1759.685 ;
      LAYER via2 ;
        RECT 2901.310 1789.280 2901.590 1789.560 ;
        RECT 2523.190 1759.360 2523.470 1759.640 ;
      LAYER met3 ;
        RECT 2901.285 1789.570 2901.615 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.285 1789.270 2924.800 1789.570 ;
        RECT 2901.285 1789.255 2901.615 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2506.000 1759.650 2510.000 1759.800 ;
        RECT 2523.165 1759.650 2523.495 1759.665 ;
        RECT 2506.000 1759.350 2523.495 1759.650 ;
        RECT 2506.000 1759.200 2510.000 1759.350 ;
        RECT 2523.165 1759.335 2523.495 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 1931.780 2523.030 1931.840 ;
        RECT 2901.290 1931.780 2901.610 1931.840 ;
        RECT 2522.710 1931.640 2901.610 1931.780 ;
        RECT 2522.710 1931.580 2523.030 1931.640 ;
        RECT 2901.290 1931.580 2901.610 1931.640 ;
      LAYER via ;
        RECT 2522.740 1931.580 2523.000 1931.840 ;
        RECT 2901.320 1931.580 2901.580 1931.840 ;
      LAYER met2 ;
        RECT 2901.310 2023.835 2901.590 2024.205 ;
        RECT 2901.380 1931.870 2901.520 2023.835 ;
        RECT 2522.740 1931.550 2523.000 1931.870 ;
        RECT 2901.320 1931.550 2901.580 1931.870 ;
        RECT 2522.800 1926.285 2522.940 1931.550 ;
        RECT 2522.730 1925.915 2523.010 1926.285 ;
      LAYER via2 ;
        RECT 2901.310 2023.880 2901.590 2024.160 ;
        RECT 2522.730 1925.960 2523.010 1926.240 ;
      LAYER met3 ;
        RECT 2901.285 2024.170 2901.615 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.285 2023.870 2924.800 2024.170 ;
        RECT 2901.285 2023.855 2901.615 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2506.000 1926.250 2510.000 1926.400 ;
        RECT 2522.705 1926.250 2523.035 1926.265 ;
        RECT 2506.000 1925.950 2523.035 1926.250 ;
        RECT 2506.000 1925.800 2510.000 1925.950 ;
        RECT 2522.705 1925.935 2523.035 1925.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2097.360 2525.330 2097.420 ;
        RECT 2902.210 2097.360 2902.530 2097.420 ;
        RECT 2525.010 2097.220 2902.530 2097.360 ;
        RECT 2525.010 2097.160 2525.330 2097.220 ;
        RECT 2902.210 2097.160 2902.530 2097.220 ;
      LAYER via ;
        RECT 2525.040 2097.160 2525.300 2097.420 ;
        RECT 2902.240 2097.160 2902.500 2097.420 ;
      LAYER met2 ;
        RECT 2902.230 2258.435 2902.510 2258.805 ;
        RECT 2902.300 2097.450 2902.440 2258.435 ;
        RECT 2525.040 2097.130 2525.300 2097.450 ;
        RECT 2902.240 2097.130 2902.500 2097.450 ;
        RECT 2525.100 2092.885 2525.240 2097.130 ;
        RECT 2525.030 2092.515 2525.310 2092.885 ;
      LAYER via2 ;
        RECT 2902.230 2258.480 2902.510 2258.760 ;
        RECT 2525.030 2092.560 2525.310 2092.840 ;
      LAYER met3 ;
        RECT 2902.205 2258.770 2902.535 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2902.205 2258.470 2924.800 2258.770 ;
        RECT 2902.205 2258.455 2902.535 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2506.000 2092.850 2510.000 2093.000 ;
        RECT 2525.005 2092.850 2525.335 2092.865 ;
        RECT 2506.000 2092.550 2525.335 2092.850 ;
        RECT 2506.000 2092.400 2510.000 2092.550 ;
        RECT 2525.005 2092.535 2525.335 2092.550 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 422.810 503.440 423.130 503.500 ;
        RECT 427.410 503.440 427.730 503.500 ;
        RECT 422.810 503.300 427.730 503.440 ;
        RECT 422.810 503.240 423.130 503.300 ;
        RECT 427.410 503.240 427.730 503.300 ;
        RECT 427.410 24.040 427.730 24.100 ;
        RECT 633.030 24.040 633.350 24.100 ;
        RECT 427.410 23.900 633.350 24.040 ;
        RECT 427.410 23.840 427.730 23.900 ;
        RECT 633.030 23.840 633.350 23.900 ;
      LAYER via ;
        RECT 422.840 503.240 423.100 503.500 ;
        RECT 427.440 503.240 427.700 503.500 ;
        RECT 427.440 23.840 427.700 24.100 ;
        RECT 633.060 23.840 633.320 24.100 ;
      LAYER met2 ;
        RECT 422.970 510.340 423.250 514.000 ;
        RECT 422.900 510.000 423.250 510.340 ;
        RECT 422.900 503.530 423.040 510.000 ;
        RECT 422.840 503.210 423.100 503.530 ;
        RECT 427.440 503.210 427.700 503.530 ;
        RECT 427.500 24.130 427.640 503.210 ;
        RECT 427.440 23.810 427.700 24.130 ;
        RECT 633.060 23.810 633.320 24.130 ;
        RECT 633.120 2.400 633.260 23.810 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2054.965 386.665 2055.135 410.635 ;
        RECT 2053.585 254.745 2053.755 282.795 ;
        RECT 2054.505 131.325 2054.675 179.435 ;
        RECT 2054.505 41.905 2054.675 110.755 ;
        RECT 2054.505 30.685 2054.675 41.395 ;
      LAYER mcon ;
        RECT 2054.965 410.465 2055.135 410.635 ;
        RECT 2053.585 282.625 2053.755 282.795 ;
        RECT 2054.505 179.265 2054.675 179.435 ;
        RECT 2054.505 110.585 2054.675 110.755 ;
        RECT 2054.505 41.225 2054.675 41.395 ;
      LAYER met1 ;
        RECT 2054.890 435.100 2055.210 435.160 ;
        RECT 2055.350 435.100 2055.670 435.160 ;
        RECT 2054.890 434.960 2055.670 435.100 ;
        RECT 2054.890 434.900 2055.210 434.960 ;
        RECT 2055.350 434.900 2055.670 434.960 ;
        RECT 2054.890 410.620 2055.210 410.680 ;
        RECT 2054.695 410.480 2055.210 410.620 ;
        RECT 2054.890 410.420 2055.210 410.480 ;
        RECT 2054.890 386.820 2055.210 386.880 ;
        RECT 2054.695 386.680 2055.210 386.820 ;
        RECT 2054.890 386.620 2055.210 386.680 ;
        RECT 2054.430 351.940 2054.750 352.200 ;
        RECT 2054.520 351.460 2054.660 351.940 ;
        RECT 2054.890 351.460 2055.210 351.520 ;
        RECT 2054.520 351.320 2055.210 351.460 ;
        RECT 2054.890 351.260 2055.210 351.320 ;
        RECT 2053.510 307.260 2053.830 307.320 ;
        RECT 2054.890 307.260 2055.210 307.320 ;
        RECT 2053.510 307.120 2055.210 307.260 ;
        RECT 2053.510 307.060 2053.830 307.120 ;
        RECT 2054.890 307.060 2055.210 307.120 ;
        RECT 2053.510 282.780 2053.830 282.840 ;
        RECT 2053.315 282.640 2053.830 282.780 ;
        RECT 2053.510 282.580 2053.830 282.640 ;
        RECT 2053.525 254.900 2053.815 254.945 ;
        RECT 2054.890 254.900 2055.210 254.960 ;
        RECT 2053.525 254.760 2055.210 254.900 ;
        RECT 2053.525 254.715 2053.815 254.760 ;
        RECT 2054.890 254.700 2055.210 254.760 ;
        RECT 2054.430 179.420 2054.750 179.480 ;
        RECT 2054.235 179.280 2054.750 179.420 ;
        RECT 2054.430 179.220 2054.750 179.280 ;
        RECT 2054.445 131.480 2054.735 131.525 ;
        RECT 2054.890 131.480 2055.210 131.540 ;
        RECT 2054.445 131.340 2055.210 131.480 ;
        RECT 2054.445 131.295 2054.735 131.340 ;
        RECT 2054.890 131.280 2055.210 131.340 ;
        RECT 2054.445 110.740 2054.735 110.785 ;
        RECT 2054.890 110.740 2055.210 110.800 ;
        RECT 2054.445 110.600 2055.210 110.740 ;
        RECT 2054.445 110.555 2054.735 110.600 ;
        RECT 2054.890 110.540 2055.210 110.600 ;
        RECT 2054.430 42.060 2054.750 42.120 ;
        RECT 2054.235 41.920 2054.750 42.060 ;
        RECT 2054.430 41.860 2054.750 41.920 ;
        RECT 2054.430 41.380 2054.750 41.440 ;
        RECT 2054.235 41.240 2054.750 41.380 ;
        RECT 2054.430 41.180 2054.750 41.240 ;
        RECT 2054.445 30.840 2054.735 30.885 ;
        RECT 2417.370 30.840 2417.690 30.900 ;
        RECT 2054.445 30.700 2417.690 30.840 ;
        RECT 2054.445 30.655 2054.735 30.700 ;
        RECT 2417.370 30.640 2417.690 30.700 ;
      LAYER via ;
        RECT 2054.920 434.900 2055.180 435.160 ;
        RECT 2055.380 434.900 2055.640 435.160 ;
        RECT 2054.920 410.420 2055.180 410.680 ;
        RECT 2054.920 386.620 2055.180 386.880 ;
        RECT 2054.460 351.940 2054.720 352.200 ;
        RECT 2054.920 351.260 2055.180 351.520 ;
        RECT 2053.540 307.060 2053.800 307.320 ;
        RECT 2054.920 307.060 2055.180 307.320 ;
        RECT 2053.540 282.580 2053.800 282.840 ;
        RECT 2054.920 254.700 2055.180 254.960 ;
        RECT 2054.460 179.220 2054.720 179.480 ;
        RECT 2054.920 131.280 2055.180 131.540 ;
        RECT 2054.920 110.540 2055.180 110.800 ;
        RECT 2054.460 41.860 2054.720 42.120 ;
        RECT 2054.460 41.180 2054.720 41.440 ;
        RECT 2417.400 30.640 2417.660 30.900 ;
      LAYER met2 ;
        RECT 2055.050 511.090 2055.330 514.000 ;
        RECT 2055.050 510.950 2056.040 511.090 ;
        RECT 2055.050 510.000 2055.330 510.950 ;
        RECT 2055.900 499.530 2056.040 510.950 ;
        RECT 2055.440 499.390 2056.040 499.530 ;
        RECT 2055.440 435.190 2055.580 499.390 ;
        RECT 2054.920 434.870 2055.180 435.190 ;
        RECT 2055.380 434.870 2055.640 435.190 ;
        RECT 2054.980 410.710 2055.120 434.870 ;
        RECT 2054.920 410.390 2055.180 410.710 ;
        RECT 2054.920 386.650 2055.180 386.910 ;
        RECT 2054.520 386.590 2055.180 386.650 ;
        RECT 2054.520 386.510 2055.120 386.590 ;
        RECT 2054.520 352.230 2054.660 386.510 ;
        RECT 2054.460 351.910 2054.720 352.230 ;
        RECT 2054.920 351.230 2055.180 351.550 ;
        RECT 2054.980 307.350 2055.120 351.230 ;
        RECT 2053.540 307.030 2053.800 307.350 ;
        RECT 2054.920 307.030 2055.180 307.350 ;
        RECT 2053.600 282.870 2053.740 307.030 ;
        RECT 2053.540 282.550 2053.800 282.870 ;
        RECT 2054.920 254.670 2055.180 254.990 ;
        RECT 2054.980 207.925 2055.120 254.670 ;
        RECT 2054.910 207.555 2055.190 207.925 ;
        RECT 2054.450 179.675 2054.730 180.045 ;
        RECT 2054.520 179.510 2054.660 179.675 ;
        RECT 2054.460 179.190 2054.720 179.510 ;
        RECT 2054.920 131.250 2055.180 131.570 ;
        RECT 2054.980 110.830 2055.120 131.250 ;
        RECT 2054.920 110.510 2055.180 110.830 ;
        RECT 2054.460 41.830 2054.720 42.150 ;
        RECT 2054.520 41.470 2054.660 41.830 ;
        RECT 2054.460 41.150 2054.720 41.470 ;
        RECT 2417.400 30.610 2417.660 30.930 ;
        RECT 2417.460 2.400 2417.600 30.610 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 2054.910 207.600 2055.190 207.880 ;
        RECT 2054.450 179.720 2054.730 180.000 ;
      LAYER met3 ;
        RECT 2054.885 207.900 2055.215 207.905 ;
        RECT 2054.630 207.890 2055.215 207.900 ;
        RECT 2054.430 207.590 2055.215 207.890 ;
        RECT 2054.630 207.580 2055.215 207.590 ;
        RECT 2054.885 207.575 2055.215 207.580 ;
        RECT 2054.425 180.020 2054.755 180.025 ;
        RECT 2054.425 180.010 2055.010 180.020 ;
        RECT 2054.425 179.710 2055.210 180.010 ;
        RECT 2054.425 179.700 2055.010 179.710 ;
        RECT 2054.425 179.695 2054.755 179.700 ;
      LAYER via3 ;
        RECT 2054.660 207.580 2054.980 207.900 ;
        RECT 2054.660 179.700 2054.980 180.020 ;
      LAYER met4 ;
        RECT 2054.655 207.575 2054.985 207.905 ;
        RECT 2054.670 180.025 2054.970 207.575 ;
        RECT 2054.655 179.695 2054.985 180.025 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2071.450 500.380 2071.770 500.440 ;
        RECT 2190.590 500.380 2190.910 500.440 ;
        RECT 2071.450 500.240 2190.910 500.380 ;
        RECT 2071.450 500.180 2071.770 500.240 ;
        RECT 2190.590 500.180 2190.910 500.240 ;
        RECT 2190.590 44.780 2190.910 44.840 ;
        RECT 2434.850 44.780 2435.170 44.840 ;
        RECT 2190.590 44.640 2435.170 44.780 ;
        RECT 2190.590 44.580 2190.910 44.640 ;
        RECT 2434.850 44.580 2435.170 44.640 ;
      LAYER via ;
        RECT 2071.480 500.180 2071.740 500.440 ;
        RECT 2190.620 500.180 2190.880 500.440 ;
        RECT 2190.620 44.580 2190.880 44.840 ;
        RECT 2434.880 44.580 2435.140 44.840 ;
      LAYER met2 ;
        RECT 2071.610 510.340 2071.890 514.000 ;
        RECT 2071.540 510.000 2071.890 510.340 ;
        RECT 2071.540 500.470 2071.680 510.000 ;
        RECT 2071.480 500.150 2071.740 500.470 ;
        RECT 2190.620 500.150 2190.880 500.470 ;
        RECT 2190.680 44.870 2190.820 500.150 ;
        RECT 2190.620 44.550 2190.880 44.870 ;
        RECT 2434.880 44.550 2435.140 44.870 ;
        RECT 2434.940 2.400 2435.080 44.550 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 24.040 2090.630 24.100 ;
        RECT 2452.790 24.040 2453.110 24.100 ;
        RECT 2090.310 23.900 2453.110 24.040 ;
        RECT 2090.310 23.840 2090.630 23.900 ;
        RECT 2452.790 23.840 2453.110 23.900 ;
      LAYER via ;
        RECT 2090.340 23.840 2090.600 24.100 ;
        RECT 2452.820 23.840 2453.080 24.100 ;
      LAYER met2 ;
        RECT 2087.710 510.410 2087.990 514.000 ;
        RECT 2087.710 510.270 2090.540 510.410 ;
        RECT 2087.710 510.000 2087.990 510.270 ;
        RECT 2090.400 24.130 2090.540 510.270 ;
        RECT 2090.340 23.810 2090.600 24.130 ;
        RECT 2452.820 23.810 2453.080 24.130 ;
        RECT 2452.880 2.400 2453.020 23.810 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 37.980 2104.430 38.040 ;
        RECT 2470.730 37.980 2471.050 38.040 ;
        RECT 2104.110 37.840 2471.050 37.980 ;
        RECT 2104.110 37.780 2104.430 37.840 ;
        RECT 2470.730 37.780 2471.050 37.840 ;
      LAYER via ;
        RECT 2104.140 37.780 2104.400 38.040 ;
        RECT 2470.760 37.780 2471.020 38.040 ;
      LAYER met2 ;
        RECT 2104.270 510.340 2104.550 514.000 ;
        RECT 2104.200 510.000 2104.550 510.340 ;
        RECT 2104.200 38.070 2104.340 510.000 ;
        RECT 2104.140 37.750 2104.400 38.070 ;
        RECT 2470.760 37.750 2471.020 38.070 ;
        RECT 2470.820 2.400 2470.960 37.750 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2120.210 503.440 2120.530 503.500 ;
        RECT 2124.810 503.440 2125.130 503.500 ;
        RECT 2120.210 503.300 2125.130 503.440 ;
        RECT 2120.210 503.240 2120.530 503.300 ;
        RECT 2124.810 503.240 2125.130 503.300 ;
        RECT 2124.810 51.580 2125.130 51.640 ;
        RECT 2488.670 51.580 2488.990 51.640 ;
        RECT 2124.810 51.440 2488.990 51.580 ;
        RECT 2124.810 51.380 2125.130 51.440 ;
        RECT 2488.670 51.380 2488.990 51.440 ;
      LAYER via ;
        RECT 2120.240 503.240 2120.500 503.500 ;
        RECT 2124.840 503.240 2125.100 503.500 ;
        RECT 2124.840 51.380 2125.100 51.640 ;
        RECT 2488.700 51.380 2488.960 51.640 ;
      LAYER met2 ;
        RECT 2120.370 510.340 2120.650 514.000 ;
        RECT 2120.300 510.000 2120.650 510.340 ;
        RECT 2120.300 503.530 2120.440 510.000 ;
        RECT 2120.240 503.210 2120.500 503.530 ;
        RECT 2124.840 503.210 2125.100 503.530 ;
        RECT 2124.900 51.670 2125.040 503.210 ;
        RECT 2124.840 51.350 2125.100 51.670 ;
        RECT 2488.700 51.350 2488.960 51.670 ;
        RECT 2488.760 2.400 2488.900 51.350 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2138.610 59.060 2138.930 59.120 ;
        RECT 2506.150 59.060 2506.470 59.120 ;
        RECT 2138.610 58.920 2506.470 59.060 ;
        RECT 2138.610 58.860 2138.930 58.920 ;
        RECT 2506.150 58.860 2506.470 58.920 ;
      LAYER via ;
        RECT 2138.640 58.860 2138.900 59.120 ;
        RECT 2506.180 58.860 2506.440 59.120 ;
      LAYER met2 ;
        RECT 2136.470 510.410 2136.750 514.000 ;
        RECT 2136.470 510.270 2138.840 510.410 ;
        RECT 2136.470 510.000 2136.750 510.270 ;
        RECT 2138.700 59.150 2138.840 510.270 ;
        RECT 2138.640 58.830 2138.900 59.150 ;
        RECT 2506.180 58.830 2506.440 59.150 ;
        RECT 2506.240 2.400 2506.380 58.830 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.870 500.040 2153.190 500.100 ;
        RECT 2514.890 500.040 2515.210 500.100 ;
        RECT 2152.870 499.900 2515.210 500.040 ;
        RECT 2152.870 499.840 2153.190 499.900 ;
        RECT 2514.890 499.840 2515.210 499.900 ;
        RECT 2514.890 27.440 2515.210 27.500 ;
        RECT 2524.090 27.440 2524.410 27.500 ;
        RECT 2514.890 27.300 2524.410 27.440 ;
        RECT 2514.890 27.240 2515.210 27.300 ;
        RECT 2524.090 27.240 2524.410 27.300 ;
      LAYER via ;
        RECT 2152.900 499.840 2153.160 500.100 ;
        RECT 2514.920 499.840 2515.180 500.100 ;
        RECT 2514.920 27.240 2515.180 27.500 ;
        RECT 2524.120 27.240 2524.380 27.500 ;
      LAYER met2 ;
        RECT 2153.030 510.340 2153.310 514.000 ;
        RECT 2152.960 510.000 2153.310 510.340 ;
        RECT 2152.960 500.130 2153.100 510.000 ;
        RECT 2152.900 499.810 2153.160 500.130 ;
        RECT 2514.920 499.810 2515.180 500.130 ;
        RECT 2514.980 27.530 2515.120 499.810 ;
        RECT 2514.920 27.210 2515.180 27.530 ;
        RECT 2524.120 27.210 2524.380 27.530 ;
        RECT 2524.180 2.400 2524.320 27.210 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2168.970 496.980 2169.290 497.040 ;
        RECT 2173.110 496.980 2173.430 497.040 ;
        RECT 2168.970 496.840 2173.430 496.980 ;
        RECT 2168.970 496.780 2169.290 496.840 ;
        RECT 2173.110 496.780 2173.430 496.840 ;
        RECT 2173.110 65.520 2173.430 65.580 ;
        RECT 2539.270 65.520 2539.590 65.580 ;
        RECT 2173.110 65.380 2539.590 65.520 ;
        RECT 2173.110 65.320 2173.430 65.380 ;
        RECT 2539.270 65.320 2539.590 65.380 ;
      LAYER via ;
        RECT 2169.000 496.780 2169.260 497.040 ;
        RECT 2173.140 496.780 2173.400 497.040 ;
        RECT 2173.140 65.320 2173.400 65.580 ;
        RECT 2539.300 65.320 2539.560 65.580 ;
      LAYER met2 ;
        RECT 2169.130 510.340 2169.410 514.000 ;
        RECT 2169.060 510.000 2169.410 510.340 ;
        RECT 2169.060 497.070 2169.200 510.000 ;
        RECT 2169.000 496.750 2169.260 497.070 ;
        RECT 2173.140 496.750 2173.400 497.070 ;
        RECT 2173.200 65.610 2173.340 496.750 ;
        RECT 2173.140 65.290 2173.400 65.610 ;
        RECT 2539.300 65.290 2539.560 65.610 ;
        RECT 2539.360 17.410 2539.500 65.290 ;
        RECT 2539.360 17.270 2542.260 17.410 ;
        RECT 2542.120 2.400 2542.260 17.270 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 79.460 2187.230 79.520 ;
        RECT 2560.430 79.460 2560.750 79.520 ;
        RECT 2186.910 79.320 2560.750 79.460 ;
        RECT 2186.910 79.260 2187.230 79.320 ;
        RECT 2560.430 79.260 2560.750 79.320 ;
      LAYER via ;
        RECT 2186.940 79.260 2187.200 79.520 ;
        RECT 2560.460 79.260 2560.720 79.520 ;
      LAYER met2 ;
        RECT 2185.690 510.410 2185.970 514.000 ;
        RECT 2185.690 510.270 2187.140 510.410 ;
        RECT 2185.690 510.000 2185.970 510.270 ;
        RECT 2187.000 79.550 2187.140 510.270 ;
        RECT 2186.940 79.230 2187.200 79.550 ;
        RECT 2560.460 79.230 2560.720 79.550 ;
        RECT 2560.520 7.210 2560.660 79.230 ;
        RECT 2560.060 7.070 2560.660 7.210 ;
        RECT 2560.060 2.400 2560.200 7.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2201.630 493.240 2201.950 493.300 ;
        RECT 2573.770 493.240 2574.090 493.300 ;
        RECT 2201.630 493.100 2574.090 493.240 ;
        RECT 2201.630 493.040 2201.950 493.100 ;
        RECT 2573.770 493.040 2574.090 493.100 ;
      LAYER via ;
        RECT 2201.660 493.040 2201.920 493.300 ;
        RECT 2573.800 493.040 2574.060 493.300 ;
      LAYER met2 ;
        RECT 2201.790 510.340 2202.070 514.000 ;
        RECT 2201.720 510.000 2202.070 510.340 ;
        RECT 2201.720 493.330 2201.860 510.000 ;
        RECT 2201.660 493.010 2201.920 493.330 ;
        RECT 2573.800 493.010 2574.060 493.330 ;
        RECT 2573.860 17.410 2574.000 493.010 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 500.040 586.430 500.100 ;
        RECT 807.830 500.040 808.150 500.100 ;
        RECT 586.110 499.900 808.150 500.040 ;
        RECT 586.110 499.840 586.430 499.900 ;
        RECT 807.830 499.840 808.150 499.900 ;
      LAYER via ;
        RECT 586.140 499.840 586.400 500.100 ;
        RECT 807.860 499.840 808.120 500.100 ;
      LAYER met2 ;
        RECT 586.270 510.340 586.550 514.000 ;
        RECT 586.200 510.000 586.550 510.340 ;
        RECT 586.200 500.130 586.340 510.000 ;
        RECT 586.140 499.810 586.400 500.130 ;
        RECT 807.860 499.810 808.120 500.130 ;
        RECT 807.920 17.410 808.060 499.810 ;
        RECT 807.920 17.270 811.740 17.410 ;
        RECT 811.600 2.400 811.740 17.270 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2218.190 486.440 2218.510 486.500 ;
        RECT 2594.470 486.440 2594.790 486.500 ;
        RECT 2218.190 486.300 2594.790 486.440 ;
        RECT 2218.190 486.240 2218.510 486.300 ;
        RECT 2594.470 486.240 2594.790 486.300 ;
      LAYER via ;
        RECT 2218.220 486.240 2218.480 486.500 ;
        RECT 2594.500 486.240 2594.760 486.500 ;
      LAYER met2 ;
        RECT 2218.350 510.340 2218.630 514.000 ;
        RECT 2218.280 510.000 2218.630 510.340 ;
        RECT 2218.280 486.530 2218.420 510.000 ;
        RECT 2218.220 486.210 2218.480 486.530 ;
        RECT 2594.500 486.210 2594.760 486.530 ;
        RECT 2594.560 17.410 2594.700 486.210 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2234.290 479.640 2234.610 479.700 ;
        RECT 2608.270 479.640 2608.590 479.700 ;
        RECT 2234.290 479.500 2608.590 479.640 ;
        RECT 2234.290 479.440 2234.610 479.500 ;
        RECT 2608.270 479.440 2608.590 479.500 ;
      LAYER via ;
        RECT 2234.320 479.440 2234.580 479.700 ;
        RECT 2608.300 479.440 2608.560 479.700 ;
      LAYER met2 ;
        RECT 2234.450 510.340 2234.730 514.000 ;
        RECT 2234.380 510.000 2234.730 510.340 ;
        RECT 2234.380 479.730 2234.520 510.000 ;
        RECT 2234.320 479.410 2234.580 479.730 ;
        RECT 2608.300 479.410 2608.560 479.730 ;
        RECT 2608.360 17.410 2608.500 479.410 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2250.850 496.980 2251.170 497.040 ;
        RECT 2255.910 496.980 2256.230 497.040 ;
        RECT 2250.850 496.840 2256.230 496.980 ;
        RECT 2250.850 496.780 2251.170 496.840 ;
        RECT 2255.910 496.780 2256.230 496.840 ;
        RECT 2255.910 86.260 2256.230 86.320 ;
        RECT 2628.970 86.260 2629.290 86.320 ;
        RECT 2255.910 86.120 2629.290 86.260 ;
        RECT 2255.910 86.060 2256.230 86.120 ;
        RECT 2628.970 86.060 2629.290 86.120 ;
      LAYER via ;
        RECT 2250.880 496.780 2251.140 497.040 ;
        RECT 2255.940 496.780 2256.200 497.040 ;
        RECT 2255.940 86.060 2256.200 86.320 ;
        RECT 2629.000 86.060 2629.260 86.320 ;
      LAYER met2 ;
        RECT 2251.010 510.340 2251.290 514.000 ;
        RECT 2250.940 510.000 2251.290 510.340 ;
        RECT 2250.940 497.070 2251.080 510.000 ;
        RECT 2250.880 496.750 2251.140 497.070 ;
        RECT 2255.940 496.750 2256.200 497.070 ;
        RECT 2256.000 86.350 2256.140 496.750 ;
        RECT 2255.940 86.030 2256.200 86.350 ;
        RECT 2629.000 86.030 2629.260 86.350 ;
        RECT 2629.060 17.410 2629.200 86.030 ;
        RECT 2629.060 17.270 2631.500 17.410 ;
        RECT 2631.360 2.400 2631.500 17.270 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 113.800 2270.030 113.860 ;
        RECT 2643.230 113.800 2643.550 113.860 ;
        RECT 2269.710 113.660 2643.550 113.800 ;
        RECT 2269.710 113.600 2270.030 113.660 ;
        RECT 2643.230 113.600 2643.550 113.660 ;
        RECT 2643.230 20.980 2643.550 21.040 ;
        RECT 2649.210 20.980 2649.530 21.040 ;
        RECT 2643.230 20.840 2649.530 20.980 ;
        RECT 2643.230 20.780 2643.550 20.840 ;
        RECT 2649.210 20.780 2649.530 20.840 ;
      LAYER via ;
        RECT 2269.740 113.600 2270.000 113.860 ;
        RECT 2643.260 113.600 2643.520 113.860 ;
        RECT 2643.260 20.780 2643.520 21.040 ;
        RECT 2649.240 20.780 2649.500 21.040 ;
      LAYER met2 ;
        RECT 2267.110 510.410 2267.390 514.000 ;
        RECT 2267.110 510.270 2269.940 510.410 ;
        RECT 2267.110 510.000 2267.390 510.270 ;
        RECT 2269.800 113.890 2269.940 510.270 ;
        RECT 2269.740 113.570 2270.000 113.890 ;
        RECT 2643.260 113.570 2643.520 113.890 ;
        RECT 2643.320 21.070 2643.460 113.570 ;
        RECT 2643.260 20.750 2643.520 21.070 ;
        RECT 2649.240 20.750 2649.500 21.070 ;
        RECT 2649.300 2.400 2649.440 20.750 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2283.510 93.060 2283.830 93.120 ;
        RECT 2663.470 93.060 2663.790 93.120 ;
        RECT 2283.510 92.920 2663.790 93.060 ;
        RECT 2283.510 92.860 2283.830 92.920 ;
        RECT 2663.470 92.860 2663.790 92.920 ;
      LAYER via ;
        RECT 2283.540 92.860 2283.800 93.120 ;
        RECT 2663.500 92.860 2663.760 93.120 ;
      LAYER met2 ;
        RECT 2283.670 510.340 2283.950 514.000 ;
        RECT 2283.600 510.000 2283.950 510.340 ;
        RECT 2283.600 93.150 2283.740 510.000 ;
        RECT 2283.540 92.830 2283.800 93.150 ;
        RECT 2663.500 92.830 2663.760 93.150 ;
        RECT 2663.560 17.410 2663.700 92.830 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2299.610 503.440 2299.930 503.500 ;
        RECT 2304.210 503.440 2304.530 503.500 ;
        RECT 2299.610 503.300 2304.530 503.440 ;
        RECT 2299.610 503.240 2299.930 503.300 ;
        RECT 2304.210 503.240 2304.530 503.300 ;
        RECT 2304.210 72.320 2304.530 72.380 ;
        RECT 2684.630 72.320 2684.950 72.380 ;
        RECT 2304.210 72.180 2684.950 72.320 ;
        RECT 2304.210 72.120 2304.530 72.180 ;
        RECT 2684.630 72.120 2684.950 72.180 ;
      LAYER via ;
        RECT 2299.640 503.240 2299.900 503.500 ;
        RECT 2304.240 503.240 2304.500 503.500 ;
        RECT 2304.240 72.120 2304.500 72.380 ;
        RECT 2684.660 72.120 2684.920 72.380 ;
      LAYER met2 ;
        RECT 2299.770 510.340 2300.050 514.000 ;
        RECT 2299.700 510.000 2300.050 510.340 ;
        RECT 2299.700 503.530 2299.840 510.000 ;
        RECT 2299.640 503.210 2299.900 503.530 ;
        RECT 2304.240 503.210 2304.500 503.530 ;
        RECT 2304.300 72.410 2304.440 503.210 ;
        RECT 2304.240 72.090 2304.500 72.410 ;
        RECT 2684.660 72.090 2684.920 72.410 ;
        RECT 2684.720 2.400 2684.860 72.090 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2318.010 99.860 2318.330 99.920 ;
        RECT 2697.970 99.860 2698.290 99.920 ;
        RECT 2318.010 99.720 2698.290 99.860 ;
        RECT 2318.010 99.660 2318.330 99.720 ;
        RECT 2697.970 99.660 2698.290 99.720 ;
      LAYER via ;
        RECT 2318.040 99.660 2318.300 99.920 ;
        RECT 2698.000 99.660 2698.260 99.920 ;
      LAYER met2 ;
        RECT 2316.330 510.410 2316.610 514.000 ;
        RECT 2316.330 510.270 2318.240 510.410 ;
        RECT 2316.330 510.000 2316.610 510.270 ;
        RECT 2318.100 99.950 2318.240 510.270 ;
        RECT 2318.040 99.630 2318.300 99.950 ;
        RECT 2698.000 99.630 2698.260 99.950 ;
        RECT 2698.060 17.410 2698.200 99.630 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2332.270 496.980 2332.590 497.040 ;
        RECT 2338.710 496.980 2339.030 497.040 ;
        RECT 2332.270 496.840 2339.030 496.980 ;
        RECT 2332.270 496.780 2332.590 496.840 ;
        RECT 2338.710 496.780 2339.030 496.840 ;
        RECT 2338.710 107.000 2339.030 107.060 ;
        RECT 2718.670 107.000 2718.990 107.060 ;
        RECT 2338.710 106.860 2718.990 107.000 ;
        RECT 2338.710 106.800 2339.030 106.860 ;
        RECT 2718.670 106.800 2718.990 106.860 ;
      LAYER via ;
        RECT 2332.300 496.780 2332.560 497.040 ;
        RECT 2338.740 496.780 2339.000 497.040 ;
        RECT 2338.740 106.800 2339.000 107.060 ;
        RECT 2718.700 106.800 2718.960 107.060 ;
      LAYER met2 ;
        RECT 2332.430 510.340 2332.710 514.000 ;
        RECT 2332.360 510.000 2332.710 510.340 ;
        RECT 2332.360 497.070 2332.500 510.000 ;
        RECT 2332.300 496.750 2332.560 497.070 ;
        RECT 2338.740 496.750 2339.000 497.070 ;
        RECT 2338.800 107.090 2338.940 496.750 ;
        RECT 2338.740 106.770 2339.000 107.090 ;
        RECT 2718.700 106.770 2718.960 107.090 ;
        RECT 2718.760 17.410 2718.900 106.770 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2348.830 496.980 2349.150 497.040 ;
        RECT 2352.510 496.980 2352.830 497.040 ;
        RECT 2348.830 496.840 2352.830 496.980 ;
        RECT 2348.830 496.780 2349.150 496.840 ;
        RECT 2352.510 496.780 2352.830 496.840 ;
        RECT 2352.510 120.600 2352.830 120.660 ;
        RECT 2732.930 120.600 2733.250 120.660 ;
        RECT 2352.510 120.460 2733.250 120.600 ;
        RECT 2352.510 120.400 2352.830 120.460 ;
        RECT 2732.930 120.400 2733.250 120.460 ;
      LAYER via ;
        RECT 2348.860 496.780 2349.120 497.040 ;
        RECT 2352.540 496.780 2352.800 497.040 ;
        RECT 2352.540 120.400 2352.800 120.660 ;
        RECT 2732.960 120.400 2733.220 120.660 ;
      LAYER met2 ;
        RECT 2348.990 510.340 2349.270 514.000 ;
        RECT 2348.920 510.000 2349.270 510.340 ;
        RECT 2348.920 497.070 2349.060 510.000 ;
        RECT 2348.860 496.750 2349.120 497.070 ;
        RECT 2352.540 496.750 2352.800 497.070 ;
        RECT 2352.600 120.690 2352.740 496.750 ;
        RECT 2352.540 120.370 2352.800 120.690 ;
        RECT 2732.960 120.370 2733.220 120.690 ;
        RECT 2733.020 17.410 2733.160 120.370 ;
        RECT 2733.020 17.270 2738.680 17.410 ;
        RECT 2738.540 2.400 2738.680 17.270 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2366.310 237.900 2366.630 237.960 ;
        RECT 2753.170 237.900 2753.490 237.960 ;
        RECT 2366.310 237.760 2753.490 237.900 ;
        RECT 2366.310 237.700 2366.630 237.760 ;
        RECT 2753.170 237.700 2753.490 237.760 ;
      LAYER via ;
        RECT 2366.340 237.700 2366.600 237.960 ;
        RECT 2753.200 237.700 2753.460 237.960 ;
      LAYER met2 ;
        RECT 2365.090 510.410 2365.370 514.000 ;
        RECT 2365.090 510.270 2366.540 510.410 ;
        RECT 2365.090 510.000 2365.370 510.270 ;
        RECT 2366.400 237.990 2366.540 510.270 ;
        RECT 2366.340 237.670 2366.600 237.990 ;
        RECT 2753.200 237.670 2753.460 237.990 ;
        RECT 2753.260 17.410 2753.400 237.670 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 602.210 496.980 602.530 497.040 ;
        RECT 606.810 496.980 607.130 497.040 ;
        RECT 602.210 496.840 607.130 496.980 ;
        RECT 602.210 496.780 602.530 496.840 ;
        RECT 606.810 496.780 607.130 496.840 ;
        RECT 606.810 31.180 607.130 31.240 ;
        RECT 829.450 31.180 829.770 31.240 ;
        RECT 606.810 31.040 829.770 31.180 ;
        RECT 606.810 30.980 607.130 31.040 ;
        RECT 829.450 30.980 829.770 31.040 ;
      LAYER via ;
        RECT 602.240 496.780 602.500 497.040 ;
        RECT 606.840 496.780 607.100 497.040 ;
        RECT 606.840 30.980 607.100 31.240 ;
        RECT 829.480 30.980 829.740 31.240 ;
      LAYER met2 ;
        RECT 602.370 510.340 602.650 514.000 ;
        RECT 602.300 510.000 602.650 510.340 ;
        RECT 602.300 497.070 602.440 510.000 ;
        RECT 602.240 496.750 602.500 497.070 ;
        RECT 606.840 496.750 607.100 497.070 ;
        RECT 606.900 31.270 607.040 496.750 ;
        RECT 606.840 30.950 607.100 31.270 ;
        RECT 829.480 30.950 829.740 31.270 ;
        RECT 829.540 2.400 829.680 30.950 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2381.490 503.440 2381.810 503.500 ;
        RECT 2391.150 503.440 2391.470 503.500 ;
        RECT 2381.490 503.300 2391.470 503.440 ;
        RECT 2381.490 503.240 2381.810 503.300 ;
        RECT 2391.150 503.240 2391.470 503.300 ;
        RECT 2391.150 472.500 2391.470 472.560 ;
        RECT 2773.870 472.500 2774.190 472.560 ;
        RECT 2391.150 472.360 2774.190 472.500 ;
        RECT 2391.150 472.300 2391.470 472.360 ;
        RECT 2773.870 472.300 2774.190 472.360 ;
      LAYER via ;
        RECT 2381.520 503.240 2381.780 503.500 ;
        RECT 2391.180 503.240 2391.440 503.500 ;
        RECT 2391.180 472.300 2391.440 472.560 ;
        RECT 2773.900 472.300 2774.160 472.560 ;
      LAYER met2 ;
        RECT 2381.650 510.340 2381.930 514.000 ;
        RECT 2381.580 510.000 2381.930 510.340 ;
        RECT 2381.580 503.530 2381.720 510.000 ;
        RECT 2381.520 503.210 2381.780 503.530 ;
        RECT 2391.180 503.210 2391.440 503.530 ;
        RECT 2391.240 472.590 2391.380 503.210 ;
        RECT 2391.180 472.270 2391.440 472.590 ;
        RECT 2773.900 472.270 2774.160 472.590 ;
        RECT 2773.960 2.400 2774.100 472.270 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.810 465.700 2401.130 465.760 ;
        RECT 2787.670 465.700 2787.990 465.760 ;
        RECT 2400.810 465.560 2787.990 465.700 ;
        RECT 2400.810 465.500 2401.130 465.560 ;
        RECT 2787.670 465.500 2787.990 465.560 ;
        RECT 2787.670 62.120 2787.990 62.180 ;
        RECT 2791.810 62.120 2792.130 62.180 ;
        RECT 2787.670 61.980 2792.130 62.120 ;
        RECT 2787.670 61.920 2787.990 61.980 ;
        RECT 2791.810 61.920 2792.130 61.980 ;
      LAYER via ;
        RECT 2400.840 465.500 2401.100 465.760 ;
        RECT 2787.700 465.500 2787.960 465.760 ;
        RECT 2787.700 61.920 2787.960 62.180 ;
        RECT 2791.840 61.920 2792.100 62.180 ;
      LAYER met2 ;
        RECT 2397.750 510.410 2398.030 514.000 ;
        RECT 2397.750 510.270 2401.040 510.410 ;
        RECT 2397.750 510.000 2398.030 510.270 ;
        RECT 2400.900 465.790 2401.040 510.270 ;
        RECT 2400.840 465.470 2401.100 465.790 ;
        RECT 2787.700 465.470 2787.960 465.790 ;
        RECT 2787.760 62.210 2787.900 465.470 ;
        RECT 2787.700 61.890 2787.960 62.210 ;
        RECT 2791.840 61.890 2792.100 62.210 ;
        RECT 2791.900 2.400 2792.040 61.890 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2808.445 48.365 2808.615 96.475 ;
      LAYER mcon ;
        RECT 2808.445 96.305 2808.615 96.475 ;
      LAYER met1 ;
        RECT 2414.150 127.740 2414.470 127.800 ;
        RECT 2808.370 127.740 2808.690 127.800 ;
        RECT 2414.150 127.600 2808.690 127.740 ;
        RECT 2414.150 127.540 2414.470 127.600 ;
        RECT 2808.370 127.540 2808.690 127.600 ;
        RECT 2808.370 96.460 2808.690 96.520 ;
        RECT 2808.175 96.320 2808.690 96.460 ;
        RECT 2808.370 96.260 2808.690 96.320 ;
        RECT 2808.385 48.520 2808.675 48.565 ;
        RECT 2809.750 48.520 2810.070 48.580 ;
        RECT 2808.385 48.380 2810.070 48.520 ;
        RECT 2808.385 48.335 2808.675 48.380 ;
        RECT 2809.750 48.320 2810.070 48.380 ;
      LAYER via ;
        RECT 2414.180 127.540 2414.440 127.800 ;
        RECT 2808.400 127.540 2808.660 127.800 ;
        RECT 2808.400 96.260 2808.660 96.520 ;
        RECT 2809.780 48.320 2810.040 48.580 ;
      LAYER met2 ;
        RECT 2414.310 510.340 2414.590 514.000 ;
        RECT 2414.240 510.000 2414.590 510.340 ;
        RECT 2414.240 127.830 2414.380 510.000 ;
        RECT 2414.180 127.510 2414.440 127.830 ;
        RECT 2808.400 127.510 2808.660 127.830 ;
        RECT 2808.460 96.550 2808.600 127.510 ;
        RECT 2808.400 96.230 2808.660 96.550 ;
        RECT 2809.780 48.290 2810.040 48.610 ;
        RECT 2809.840 2.400 2809.980 48.290 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2430.250 496.980 2430.570 497.040 ;
        RECT 2435.310 496.980 2435.630 497.040 ;
        RECT 2430.250 496.840 2435.630 496.980 ;
        RECT 2430.250 496.780 2430.570 496.840 ;
        RECT 2435.310 496.780 2435.630 496.840 ;
        RECT 2435.310 44.780 2435.630 44.840 ;
        RECT 2827.690 44.780 2828.010 44.840 ;
        RECT 2435.310 44.640 2828.010 44.780 ;
        RECT 2435.310 44.580 2435.630 44.640 ;
        RECT 2827.690 44.580 2828.010 44.640 ;
      LAYER via ;
        RECT 2430.280 496.780 2430.540 497.040 ;
        RECT 2435.340 496.780 2435.600 497.040 ;
        RECT 2435.340 44.580 2435.600 44.840 ;
        RECT 2827.720 44.580 2827.980 44.840 ;
      LAYER met2 ;
        RECT 2430.410 510.340 2430.690 514.000 ;
        RECT 2430.340 510.000 2430.690 510.340 ;
        RECT 2430.340 497.070 2430.480 510.000 ;
        RECT 2430.280 496.750 2430.540 497.070 ;
        RECT 2435.340 496.750 2435.600 497.070 ;
        RECT 2435.400 44.870 2435.540 496.750 ;
        RECT 2435.340 44.550 2435.600 44.870 ;
        RECT 2827.720 44.550 2827.980 44.870 ;
        RECT 2827.780 2.400 2827.920 44.550 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2449.110 30.840 2449.430 30.900 ;
        RECT 2845.170 30.840 2845.490 30.900 ;
        RECT 2449.110 30.700 2845.490 30.840 ;
        RECT 2449.110 30.640 2449.430 30.700 ;
        RECT 2845.170 30.640 2845.490 30.700 ;
      LAYER via ;
        RECT 2449.140 30.640 2449.400 30.900 ;
        RECT 2845.200 30.640 2845.460 30.900 ;
      LAYER met2 ;
        RECT 2446.970 510.410 2447.250 514.000 ;
        RECT 2446.970 510.270 2449.340 510.410 ;
        RECT 2446.970 510.000 2447.250 510.270 ;
        RECT 2449.200 30.930 2449.340 510.270 ;
        RECT 2449.140 30.610 2449.400 30.930 ;
        RECT 2845.200 30.610 2845.460 30.930 ;
        RECT 2845.260 2.400 2845.400 30.610 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2462.910 500.380 2463.230 500.440 ;
        RECT 2804.690 500.380 2805.010 500.440 ;
        RECT 2462.910 500.240 2805.010 500.380 ;
        RECT 2462.910 500.180 2463.230 500.240 ;
        RECT 2804.690 500.180 2805.010 500.240 ;
        RECT 2804.690 24.040 2805.010 24.100 ;
        RECT 2863.110 24.040 2863.430 24.100 ;
        RECT 2804.690 23.900 2863.430 24.040 ;
        RECT 2804.690 23.840 2805.010 23.900 ;
        RECT 2863.110 23.840 2863.430 23.900 ;
      LAYER via ;
        RECT 2462.940 500.180 2463.200 500.440 ;
        RECT 2804.720 500.180 2804.980 500.440 ;
        RECT 2804.720 23.840 2804.980 24.100 ;
        RECT 2863.140 23.840 2863.400 24.100 ;
      LAYER met2 ;
        RECT 2463.070 510.340 2463.350 514.000 ;
        RECT 2463.000 510.000 2463.350 510.340 ;
        RECT 2463.000 500.470 2463.140 510.000 ;
        RECT 2462.940 500.150 2463.200 500.470 ;
        RECT 2804.720 500.150 2804.980 500.470 ;
        RECT 2804.780 24.130 2804.920 500.150 ;
        RECT 2804.720 23.810 2804.980 24.130 ;
        RECT 2863.140 23.810 2863.400 24.130 ;
        RECT 2863.200 2.400 2863.340 23.810 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2479.470 496.980 2479.790 497.040 ;
        RECT 2483.610 496.980 2483.930 497.040 ;
        RECT 2479.470 496.840 2483.930 496.980 ;
        RECT 2479.470 496.780 2479.790 496.840 ;
        RECT 2483.610 496.780 2483.930 496.840 ;
        RECT 2483.610 37.980 2483.930 38.040 ;
        RECT 2881.050 37.980 2881.370 38.040 ;
        RECT 2483.610 37.840 2881.370 37.980 ;
        RECT 2483.610 37.780 2483.930 37.840 ;
        RECT 2881.050 37.780 2881.370 37.840 ;
      LAYER via ;
        RECT 2479.500 496.780 2479.760 497.040 ;
        RECT 2483.640 496.780 2483.900 497.040 ;
        RECT 2483.640 37.780 2483.900 38.040 ;
        RECT 2881.080 37.780 2881.340 38.040 ;
      LAYER met2 ;
        RECT 2479.630 510.340 2479.910 514.000 ;
        RECT 2479.560 510.000 2479.910 510.340 ;
        RECT 2479.560 497.070 2479.700 510.000 ;
        RECT 2479.500 496.750 2479.760 497.070 ;
        RECT 2483.640 496.750 2483.900 497.070 ;
        RECT 2483.700 38.070 2483.840 496.750 ;
        RECT 2483.640 37.750 2483.900 38.070 ;
        RECT 2881.080 37.750 2881.340 38.070 ;
        RECT 2881.140 2.400 2881.280 37.750 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2497.410 51.580 2497.730 51.640 ;
        RECT 2898.070 51.580 2898.390 51.640 ;
        RECT 2497.410 51.440 2898.390 51.580 ;
        RECT 2497.410 51.380 2497.730 51.440 ;
        RECT 2898.070 51.380 2898.390 51.440 ;
        RECT 2898.070 2.960 2898.390 3.020 ;
        RECT 2898.990 2.960 2899.310 3.020 ;
        RECT 2898.070 2.820 2899.310 2.960 ;
        RECT 2898.070 2.760 2898.390 2.820 ;
        RECT 2898.990 2.760 2899.310 2.820 ;
      LAYER via ;
        RECT 2497.440 51.380 2497.700 51.640 ;
        RECT 2898.100 51.380 2898.360 51.640 ;
        RECT 2898.100 2.760 2898.360 3.020 ;
        RECT 2899.020 2.760 2899.280 3.020 ;
      LAYER met2 ;
        RECT 2495.730 510.410 2496.010 514.000 ;
        RECT 2495.730 510.270 2497.640 510.410 ;
        RECT 2495.730 510.000 2496.010 510.270 ;
        RECT 2497.500 51.670 2497.640 510.270 ;
        RECT 2497.440 51.350 2497.700 51.670 ;
        RECT 2898.100 51.350 2898.360 51.670 ;
        RECT 2898.160 3.050 2898.300 51.350 ;
        RECT 2898.100 2.730 2898.360 3.050 ;
        RECT 2899.020 2.730 2899.280 3.050 ;
        RECT 2899.080 2.400 2899.220 2.730 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 37.980 620.930 38.040 ;
        RECT 846.930 37.980 847.250 38.040 ;
        RECT 620.610 37.840 847.250 37.980 ;
        RECT 620.610 37.780 620.930 37.840 ;
        RECT 846.930 37.780 847.250 37.840 ;
      LAYER via ;
        RECT 620.640 37.780 620.900 38.040 ;
        RECT 846.960 37.780 847.220 38.040 ;
      LAYER met2 ;
        RECT 618.930 510.410 619.210 514.000 ;
        RECT 618.930 510.270 620.840 510.410 ;
        RECT 618.930 510.000 619.210 510.270 ;
        RECT 620.700 38.070 620.840 510.270 ;
        RECT 620.640 37.750 620.900 38.070 ;
        RECT 846.960 37.750 847.220 38.070 ;
        RECT 847.020 2.400 847.160 37.750 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.870 496.980 635.190 497.040 ;
        RECT 644.990 496.980 645.310 497.040 ;
        RECT 634.870 496.840 645.310 496.980 ;
        RECT 634.870 496.780 635.190 496.840 ;
        RECT 644.990 496.780 645.310 496.840 ;
        RECT 644.990 24.040 645.310 24.100 ;
        RECT 864.870 24.040 865.190 24.100 ;
        RECT 644.990 23.900 865.190 24.040 ;
        RECT 644.990 23.840 645.310 23.900 ;
        RECT 864.870 23.840 865.190 23.900 ;
      LAYER via ;
        RECT 634.900 496.780 635.160 497.040 ;
        RECT 645.020 496.780 645.280 497.040 ;
        RECT 645.020 23.840 645.280 24.100 ;
        RECT 864.900 23.840 865.160 24.100 ;
      LAYER met2 ;
        RECT 635.030 510.340 635.310 514.000 ;
        RECT 634.960 510.000 635.310 510.340 ;
        RECT 634.960 497.070 635.100 510.000 ;
        RECT 634.900 496.750 635.160 497.070 ;
        RECT 645.020 496.750 645.280 497.070 ;
        RECT 645.080 24.130 645.220 496.750 ;
        RECT 645.020 23.810 645.280 24.130 ;
        RECT 864.900 23.810 865.160 24.130 ;
        RECT 864.960 2.400 865.100 23.810 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 651.430 496.980 651.750 497.040 ;
        RECT 655.110 496.980 655.430 497.040 ;
        RECT 651.430 496.840 655.430 496.980 ;
        RECT 651.430 496.780 651.750 496.840 ;
        RECT 655.110 496.780 655.430 496.840 ;
        RECT 655.110 44.780 655.430 44.840 ;
        RECT 882.810 44.780 883.130 44.840 ;
        RECT 655.110 44.640 883.130 44.780 ;
        RECT 655.110 44.580 655.430 44.640 ;
        RECT 882.810 44.580 883.130 44.640 ;
      LAYER via ;
        RECT 651.460 496.780 651.720 497.040 ;
        RECT 655.140 496.780 655.400 497.040 ;
        RECT 655.140 44.580 655.400 44.840 ;
        RECT 882.840 44.580 883.100 44.840 ;
      LAYER met2 ;
        RECT 651.590 510.340 651.870 514.000 ;
        RECT 651.520 510.000 651.870 510.340 ;
        RECT 651.520 497.070 651.660 510.000 ;
        RECT 651.460 496.750 651.720 497.070 ;
        RECT 655.140 496.750 655.400 497.070 ;
        RECT 655.200 44.870 655.340 496.750 ;
        RECT 655.140 44.550 655.400 44.870 ;
        RECT 882.840 44.550 883.100 44.870 ;
        RECT 882.900 2.400 883.040 44.550 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 58.720 669.230 58.780 ;
        RECT 897.070 58.720 897.390 58.780 ;
        RECT 668.910 58.580 897.390 58.720 ;
        RECT 668.910 58.520 669.230 58.580 ;
        RECT 897.070 58.520 897.390 58.580 ;
      LAYER via ;
        RECT 668.940 58.520 669.200 58.780 ;
        RECT 897.100 58.520 897.360 58.780 ;
      LAYER met2 ;
        RECT 667.690 510.410 667.970 514.000 ;
        RECT 667.690 510.270 669.140 510.410 ;
        RECT 667.690 510.000 667.970 510.270 ;
        RECT 669.000 58.810 669.140 510.270 ;
        RECT 668.940 58.490 669.200 58.810 ;
        RECT 897.100 58.490 897.360 58.810 ;
        RECT 897.160 17.410 897.300 58.490 ;
        RECT 897.160 17.270 900.980 17.410 ;
        RECT 900.840 2.400 900.980 17.270 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 684.090 496.980 684.410 497.040 ;
        RECT 693.290 496.980 693.610 497.040 ;
        RECT 684.090 496.840 693.610 496.980 ;
        RECT 684.090 496.780 684.410 496.840 ;
        RECT 693.290 496.780 693.610 496.840 ;
        RECT 693.290 51.580 693.610 51.640 ;
        RECT 918.230 51.580 918.550 51.640 ;
        RECT 693.290 51.440 918.550 51.580 ;
        RECT 693.290 51.380 693.610 51.440 ;
        RECT 918.230 51.380 918.550 51.440 ;
      LAYER via ;
        RECT 684.120 496.780 684.380 497.040 ;
        RECT 693.320 496.780 693.580 497.040 ;
        RECT 693.320 51.380 693.580 51.640 ;
        RECT 918.260 51.380 918.520 51.640 ;
      LAYER met2 ;
        RECT 684.250 510.340 684.530 514.000 ;
        RECT 684.180 510.000 684.530 510.340 ;
        RECT 684.180 497.070 684.320 510.000 ;
        RECT 684.120 496.750 684.380 497.070 ;
        RECT 693.320 496.750 693.580 497.070 ;
        RECT 693.380 51.670 693.520 496.750 ;
        RECT 693.320 51.350 693.580 51.670 ;
        RECT 918.260 51.350 918.520 51.670 ;
        RECT 918.320 17.410 918.460 51.350 ;
        RECT 918.320 17.270 918.920 17.410 ;
        RECT 918.780 2.400 918.920 17.270 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 65.520 703.730 65.580 ;
        RECT 931.570 65.520 931.890 65.580 ;
        RECT 703.410 65.380 931.890 65.520 ;
        RECT 703.410 65.320 703.730 65.380 ;
        RECT 931.570 65.320 931.890 65.380 ;
      LAYER via ;
        RECT 703.440 65.320 703.700 65.580 ;
        RECT 931.600 65.320 931.860 65.580 ;
      LAYER met2 ;
        RECT 700.350 510.410 700.630 514.000 ;
        RECT 700.350 510.270 703.640 510.410 ;
        RECT 700.350 510.000 700.630 510.270 ;
        RECT 703.500 65.610 703.640 510.270 ;
        RECT 703.440 65.290 703.700 65.610 ;
        RECT 931.600 65.290 931.860 65.610 ;
        RECT 931.660 17.410 931.800 65.290 ;
        RECT 931.660 17.270 936.400 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 72.320 717.530 72.380 ;
        RECT 952.270 72.320 952.590 72.380 ;
        RECT 717.210 72.180 952.590 72.320 ;
        RECT 717.210 72.120 717.530 72.180 ;
        RECT 952.270 72.120 952.590 72.180 ;
      LAYER via ;
        RECT 717.240 72.120 717.500 72.380 ;
        RECT 952.300 72.120 952.560 72.380 ;
      LAYER met2 ;
        RECT 716.910 510.340 717.190 514.000 ;
        RECT 716.840 510.000 717.190 510.340 ;
        RECT 716.840 497.490 716.980 510.000 ;
        RECT 716.840 497.350 717.440 497.490 ;
        RECT 717.300 72.410 717.440 497.350 ;
        RECT 717.240 72.090 717.500 72.410 ;
        RECT 952.300 72.090 952.560 72.410 ;
        RECT 952.360 17.410 952.500 72.090 ;
        RECT 952.360 17.270 954.340 17.410 ;
        RECT 954.200 2.400 954.340 17.270 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 732.850 496.980 733.170 497.040 ;
        RECT 737.910 496.980 738.230 497.040 ;
        RECT 732.850 496.840 738.230 496.980 ;
        RECT 732.850 496.780 733.170 496.840 ;
        RECT 737.910 496.780 738.230 496.840 ;
        RECT 737.910 79.460 738.230 79.520 ;
        RECT 966.530 79.460 966.850 79.520 ;
        RECT 737.910 79.320 966.850 79.460 ;
        RECT 737.910 79.260 738.230 79.320 ;
        RECT 966.530 79.260 966.850 79.320 ;
      LAYER via ;
        RECT 732.880 496.780 733.140 497.040 ;
        RECT 737.940 496.780 738.200 497.040 ;
        RECT 737.940 79.260 738.200 79.520 ;
        RECT 966.560 79.260 966.820 79.520 ;
      LAYER met2 ;
        RECT 733.010 510.340 733.290 514.000 ;
        RECT 732.940 510.000 733.290 510.340 ;
        RECT 732.940 497.070 733.080 510.000 ;
        RECT 732.880 496.750 733.140 497.070 ;
        RECT 737.940 496.750 738.200 497.070 ;
        RECT 738.000 79.550 738.140 496.750 ;
        RECT 737.940 79.230 738.200 79.550 ;
        RECT 966.560 79.230 966.820 79.550 ;
        RECT 966.620 17.410 966.760 79.230 ;
        RECT 966.620 17.270 972.280 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 44.780 441.530 44.840 ;
        RECT 650.970 44.780 651.290 44.840 ;
        RECT 441.210 44.640 651.290 44.780 ;
        RECT 441.210 44.580 441.530 44.640 ;
        RECT 650.970 44.580 651.290 44.640 ;
      LAYER via ;
        RECT 441.240 44.580 441.500 44.840 ;
        RECT 651.000 44.580 651.260 44.840 ;
      LAYER met2 ;
        RECT 439.530 510.410 439.810 514.000 ;
        RECT 439.530 510.270 441.440 510.410 ;
        RECT 439.530 510.000 439.810 510.270 ;
        RECT 441.300 44.870 441.440 510.270 ;
        RECT 441.240 44.550 441.500 44.870 ;
        RECT 651.000 44.550 651.260 44.870 ;
        RECT 651.060 2.400 651.200 44.550 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 751.710 86.260 752.030 86.320 ;
        RECT 986.770 86.260 987.090 86.320 ;
        RECT 751.710 86.120 987.090 86.260 ;
        RECT 751.710 86.060 752.030 86.120 ;
        RECT 986.770 86.060 987.090 86.120 ;
      LAYER via ;
        RECT 751.740 86.060 752.000 86.320 ;
        RECT 986.800 86.060 987.060 86.320 ;
      LAYER met2 ;
        RECT 749.570 510.410 749.850 514.000 ;
        RECT 749.570 510.270 751.940 510.410 ;
        RECT 749.570 510.000 749.850 510.270 ;
        RECT 751.800 86.350 751.940 510.270 ;
        RECT 751.740 86.030 752.000 86.350 ;
        RECT 986.800 86.030 987.060 86.350 ;
        RECT 986.860 17.410 987.000 86.030 ;
        RECT 986.860 17.270 990.220 17.410 ;
        RECT 990.080 2.400 990.220 17.270 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.510 502.420 765.830 502.480 ;
        RECT 769.190 502.420 769.510 502.480 ;
        RECT 765.510 502.280 769.510 502.420 ;
        RECT 765.510 502.220 765.830 502.280 ;
        RECT 769.190 502.220 769.510 502.280 ;
        RECT 769.190 93.060 769.510 93.120 ;
        RECT 1007.930 93.060 1008.250 93.120 ;
        RECT 769.190 92.920 1008.250 93.060 ;
        RECT 769.190 92.860 769.510 92.920 ;
        RECT 1007.930 92.860 1008.250 92.920 ;
      LAYER via ;
        RECT 765.540 502.220 765.800 502.480 ;
        RECT 769.220 502.220 769.480 502.480 ;
        RECT 769.220 92.860 769.480 93.120 ;
        RECT 1007.960 92.860 1008.220 93.120 ;
      LAYER met2 ;
        RECT 765.670 510.340 765.950 514.000 ;
        RECT 765.600 510.000 765.950 510.340 ;
        RECT 765.600 502.510 765.740 510.000 ;
        RECT 765.540 502.190 765.800 502.510 ;
        RECT 769.220 502.190 769.480 502.510 ;
        RECT 769.280 93.150 769.420 502.190 ;
        RECT 769.220 92.830 769.480 93.150 ;
        RECT 1007.960 92.830 1008.220 93.150 ;
        RECT 1008.020 17.410 1008.160 92.830 ;
        RECT 1007.560 17.270 1008.160 17.410 ;
        RECT 1007.560 2.400 1007.700 17.270 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 782.070 503.440 782.390 503.500 ;
        RECT 786.210 503.440 786.530 503.500 ;
        RECT 782.070 503.300 786.530 503.440 ;
        RECT 782.070 503.240 782.390 503.300 ;
        RECT 786.210 503.240 786.530 503.300 ;
        RECT 786.210 99.860 786.530 99.920 ;
        RECT 1021.270 99.860 1021.590 99.920 ;
        RECT 786.210 99.720 1021.590 99.860 ;
        RECT 786.210 99.660 786.530 99.720 ;
        RECT 1021.270 99.660 1021.590 99.720 ;
      LAYER via ;
        RECT 782.100 503.240 782.360 503.500 ;
        RECT 786.240 503.240 786.500 503.500 ;
        RECT 786.240 99.660 786.500 99.920 ;
        RECT 1021.300 99.660 1021.560 99.920 ;
      LAYER met2 ;
        RECT 782.230 510.340 782.510 514.000 ;
        RECT 782.160 510.000 782.510 510.340 ;
        RECT 782.160 503.530 782.300 510.000 ;
        RECT 782.100 503.210 782.360 503.530 ;
        RECT 786.240 503.210 786.500 503.530 ;
        RECT 786.300 99.950 786.440 503.210 ;
        RECT 786.240 99.630 786.500 99.950 ;
        RECT 1021.300 99.630 1021.560 99.950 ;
        RECT 1021.360 17.410 1021.500 99.630 ;
        RECT 1021.360 17.270 1025.640 17.410 ;
        RECT 1025.500 2.400 1025.640 17.270 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 800.010 30.840 800.330 30.900 ;
        RECT 1043.350 30.840 1043.670 30.900 ;
        RECT 800.010 30.700 1043.670 30.840 ;
        RECT 800.010 30.640 800.330 30.700 ;
        RECT 1043.350 30.640 1043.670 30.700 ;
      LAYER via ;
        RECT 800.040 30.640 800.300 30.900 ;
        RECT 1043.380 30.640 1043.640 30.900 ;
      LAYER met2 ;
        RECT 798.330 510.410 798.610 514.000 ;
        RECT 798.330 510.270 800.240 510.410 ;
        RECT 798.330 510.000 798.610 510.270 ;
        RECT 800.100 30.930 800.240 510.270 ;
        RECT 800.040 30.610 800.300 30.930 ;
        RECT 1043.380 30.610 1043.640 30.930 ;
        RECT 1043.440 2.400 1043.580 30.610 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 814.730 500.040 815.050 500.100 ;
        RECT 1055.770 500.040 1056.090 500.100 ;
        RECT 814.730 499.900 1056.090 500.040 ;
        RECT 814.730 499.840 815.050 499.900 ;
        RECT 1055.770 499.840 1056.090 499.900 ;
      LAYER via ;
        RECT 814.760 499.840 815.020 500.100 ;
        RECT 1055.800 499.840 1056.060 500.100 ;
      LAYER met2 ;
        RECT 814.890 510.340 815.170 514.000 ;
        RECT 814.820 510.000 815.170 510.340 ;
        RECT 814.820 500.130 814.960 510.000 ;
        RECT 814.760 499.810 815.020 500.130 ;
        RECT 1055.800 499.810 1056.060 500.130 ;
        RECT 1055.860 17.410 1056.000 499.810 ;
        RECT 1055.860 17.270 1061.520 17.410 ;
        RECT 1061.380 2.400 1061.520 17.270 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 830.830 496.980 831.150 497.040 ;
        RECT 834.510 496.980 834.830 497.040 ;
        RECT 830.830 496.840 834.830 496.980 ;
        RECT 830.830 496.780 831.150 496.840 ;
        RECT 834.510 496.780 834.830 496.840 ;
        RECT 834.510 107.000 834.830 107.060 ;
        RECT 1076.470 107.000 1076.790 107.060 ;
        RECT 834.510 106.860 1076.790 107.000 ;
        RECT 834.510 106.800 834.830 106.860 ;
        RECT 1076.470 106.800 1076.790 106.860 ;
      LAYER via ;
        RECT 830.860 496.780 831.120 497.040 ;
        RECT 834.540 496.780 834.800 497.040 ;
        RECT 834.540 106.800 834.800 107.060 ;
        RECT 1076.500 106.800 1076.760 107.060 ;
      LAYER met2 ;
        RECT 830.990 510.340 831.270 514.000 ;
        RECT 830.920 510.000 831.270 510.340 ;
        RECT 830.920 497.070 831.060 510.000 ;
        RECT 830.860 496.750 831.120 497.070 ;
        RECT 834.540 496.750 834.800 497.070 ;
        RECT 834.600 107.090 834.740 496.750 ;
        RECT 834.540 106.770 834.800 107.090 ;
        RECT 1076.500 106.770 1076.760 107.090 ;
        RECT 1076.560 17.410 1076.700 106.770 ;
        RECT 1076.560 17.270 1079.460 17.410 ;
        RECT 1079.320 2.400 1079.460 17.270 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.310 224.300 848.630 224.360 ;
        RECT 1090.730 224.300 1091.050 224.360 ;
        RECT 848.310 224.160 1091.050 224.300 ;
        RECT 848.310 224.100 848.630 224.160 ;
        RECT 1090.730 224.100 1091.050 224.160 ;
        RECT 1090.730 17.920 1091.050 17.980 ;
        RECT 1096.710 17.920 1097.030 17.980 ;
        RECT 1090.730 17.780 1097.030 17.920 ;
        RECT 1090.730 17.720 1091.050 17.780 ;
        RECT 1096.710 17.720 1097.030 17.780 ;
      LAYER via ;
        RECT 848.340 224.100 848.600 224.360 ;
        RECT 1090.760 224.100 1091.020 224.360 ;
        RECT 1090.760 17.720 1091.020 17.980 ;
        RECT 1096.740 17.720 1097.000 17.980 ;
      LAYER met2 ;
        RECT 847.550 510.410 847.830 514.000 ;
        RECT 847.550 510.270 848.540 510.410 ;
        RECT 847.550 510.000 847.830 510.270 ;
        RECT 848.400 224.390 848.540 510.270 ;
        RECT 848.340 224.070 848.600 224.390 ;
        RECT 1090.760 224.070 1091.020 224.390 ;
        RECT 1090.820 18.010 1090.960 224.070 ;
        RECT 1090.760 17.690 1091.020 18.010 ;
        RECT 1096.740 17.690 1097.000 18.010 ;
        RECT 1096.800 2.400 1096.940 17.690 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 863.490 496.980 863.810 497.040 ;
        RECT 869.010 496.980 869.330 497.040 ;
        RECT 863.490 496.840 869.330 496.980 ;
        RECT 863.490 496.780 863.810 496.840 ;
        RECT 869.010 496.780 869.330 496.840 ;
        RECT 869.010 24.040 869.330 24.100 ;
        RECT 1114.650 24.040 1114.970 24.100 ;
        RECT 869.010 23.900 1114.970 24.040 ;
        RECT 869.010 23.840 869.330 23.900 ;
        RECT 1114.650 23.840 1114.970 23.900 ;
      LAYER via ;
        RECT 863.520 496.780 863.780 497.040 ;
        RECT 869.040 496.780 869.300 497.040 ;
        RECT 869.040 23.840 869.300 24.100 ;
        RECT 1114.680 23.840 1114.940 24.100 ;
      LAYER met2 ;
        RECT 863.650 510.340 863.930 514.000 ;
        RECT 863.580 510.000 863.930 510.340 ;
        RECT 863.580 497.070 863.720 510.000 ;
        RECT 863.520 496.750 863.780 497.070 ;
        RECT 869.040 496.750 869.300 497.070 ;
        RECT 869.100 24.130 869.240 496.750 ;
        RECT 869.040 23.810 869.300 24.130 ;
        RECT 1114.680 23.810 1114.940 24.130 ;
        RECT 1114.740 2.400 1114.880 23.810 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 881.890 37.980 882.210 38.040 ;
        RECT 1132.590 37.980 1132.910 38.040 ;
        RECT 881.890 37.840 1132.910 37.980 ;
        RECT 881.890 37.780 882.210 37.840 ;
        RECT 1132.590 37.780 1132.910 37.840 ;
      LAYER via ;
        RECT 881.920 37.780 882.180 38.040 ;
        RECT 1132.620 37.780 1132.880 38.040 ;
      LAYER met2 ;
        RECT 880.210 510.410 880.490 514.000 ;
        RECT 880.210 510.270 883.040 510.410 ;
        RECT 880.210 510.000 880.490 510.270 ;
        RECT 882.900 60.250 883.040 510.270 ;
        RECT 881.980 60.110 883.040 60.250 ;
        RECT 881.980 38.070 882.120 60.110 ;
        RECT 881.920 37.750 882.180 38.070 ;
        RECT 1132.620 37.750 1132.880 38.070 ;
        RECT 1132.680 2.400 1132.820 37.750 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 44.780 896.930 44.840 ;
        RECT 1150.530 44.780 1150.850 44.840 ;
        RECT 896.610 44.640 1150.850 44.780 ;
        RECT 896.610 44.580 896.930 44.640 ;
        RECT 1150.530 44.580 1150.850 44.640 ;
      LAYER via ;
        RECT 896.640 44.580 896.900 44.840 ;
        RECT 1150.560 44.580 1150.820 44.840 ;
      LAYER met2 ;
        RECT 896.310 510.340 896.590 514.000 ;
        RECT 896.240 510.000 896.590 510.340 ;
        RECT 896.240 497.490 896.380 510.000 ;
        RECT 896.240 497.350 896.840 497.490 ;
        RECT 896.700 44.870 896.840 497.350 ;
        RECT 896.640 44.550 896.900 44.870 ;
        RECT 1150.560 44.550 1150.820 44.870 ;
        RECT 1150.620 2.400 1150.760 44.550 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.470 503.100 455.790 503.160 ;
        RECT 461.910 503.100 462.230 503.160 ;
        RECT 455.470 502.960 462.230 503.100 ;
        RECT 455.470 502.900 455.790 502.960 ;
        RECT 461.910 502.900 462.230 502.960 ;
        RECT 461.910 58.720 462.230 58.780 ;
        RECT 662.930 58.720 663.250 58.780 ;
        RECT 461.910 58.580 663.250 58.720 ;
        RECT 461.910 58.520 462.230 58.580 ;
        RECT 662.930 58.520 663.250 58.580 ;
        RECT 662.930 16.900 663.250 16.960 ;
        RECT 668.910 16.900 669.230 16.960 ;
        RECT 662.930 16.760 669.230 16.900 ;
        RECT 662.930 16.700 663.250 16.760 ;
        RECT 668.910 16.700 669.230 16.760 ;
      LAYER via ;
        RECT 455.500 502.900 455.760 503.160 ;
        RECT 461.940 502.900 462.200 503.160 ;
        RECT 461.940 58.520 462.200 58.780 ;
        RECT 662.960 58.520 663.220 58.780 ;
        RECT 662.960 16.700 663.220 16.960 ;
        RECT 668.940 16.700 669.200 16.960 ;
      LAYER met2 ;
        RECT 455.630 510.340 455.910 514.000 ;
        RECT 455.560 510.000 455.910 510.340 ;
        RECT 455.560 503.190 455.700 510.000 ;
        RECT 455.500 502.870 455.760 503.190 ;
        RECT 461.940 502.870 462.200 503.190 ;
        RECT 462.000 58.810 462.140 502.870 ;
        RECT 461.940 58.490 462.200 58.810 ;
        RECT 662.960 58.490 663.220 58.810 ;
        RECT 663.020 16.990 663.160 58.490 ;
        RECT 662.960 16.670 663.220 16.990 ;
        RECT 668.940 16.670 669.200 16.990 ;
        RECT 669.000 2.400 669.140 16.670 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 496.980 913.030 497.040 ;
        RECT 917.310 496.980 917.630 497.040 ;
        RECT 912.710 496.840 917.630 496.980 ;
        RECT 912.710 496.780 913.030 496.840 ;
        RECT 917.310 496.780 917.630 496.840 ;
        RECT 917.310 58.720 917.630 58.780 ;
        RECT 1166.170 58.720 1166.490 58.780 ;
        RECT 917.310 58.580 1166.490 58.720 ;
        RECT 917.310 58.520 917.630 58.580 ;
        RECT 1166.170 58.520 1166.490 58.580 ;
      LAYER via ;
        RECT 912.740 496.780 913.000 497.040 ;
        RECT 917.340 496.780 917.600 497.040 ;
        RECT 917.340 58.520 917.600 58.780 ;
        RECT 1166.200 58.520 1166.460 58.780 ;
      LAYER met2 ;
        RECT 912.870 510.340 913.150 514.000 ;
        RECT 912.800 510.000 913.150 510.340 ;
        RECT 912.800 497.070 912.940 510.000 ;
        RECT 912.740 496.750 913.000 497.070 ;
        RECT 917.340 496.750 917.600 497.070 ;
        RECT 917.400 58.810 917.540 496.750 ;
        RECT 917.340 58.490 917.600 58.810 ;
        RECT 1166.200 58.490 1166.460 58.810 ;
        RECT 1166.260 17.410 1166.400 58.490 ;
        RECT 1166.260 17.270 1168.700 17.410 ;
        RECT 1168.560 2.400 1168.700 17.270 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 51.580 931.430 51.640 ;
        RECT 1180.430 51.580 1180.750 51.640 ;
        RECT 931.110 51.440 1180.750 51.580 ;
        RECT 931.110 51.380 931.430 51.440 ;
        RECT 1180.430 51.380 1180.750 51.440 ;
      LAYER via ;
        RECT 931.140 51.380 931.400 51.640 ;
        RECT 1180.460 51.380 1180.720 51.640 ;
      LAYER met2 ;
        RECT 928.970 510.410 929.250 514.000 ;
        RECT 928.970 510.270 931.340 510.410 ;
        RECT 928.970 510.000 929.250 510.270 ;
        RECT 931.200 51.670 931.340 510.270 ;
        RECT 931.140 51.350 931.400 51.670 ;
        RECT 1180.460 51.350 1180.720 51.670 ;
        RECT 1180.520 17.410 1180.660 51.350 ;
        RECT 1180.520 17.270 1186.180 17.410 ;
        RECT 1186.040 2.400 1186.180 17.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 944.910 496.980 945.230 497.040 ;
        RECT 948.590 496.980 948.910 497.040 ;
        RECT 944.910 496.840 948.910 496.980 ;
        RECT 944.910 496.780 945.230 496.840 ;
        RECT 948.590 496.780 948.910 496.840 ;
        RECT 948.590 65.520 948.910 65.580 ;
        RECT 1200.670 65.520 1200.990 65.580 ;
        RECT 948.590 65.380 1200.990 65.520 ;
        RECT 948.590 65.320 948.910 65.380 ;
        RECT 1200.670 65.320 1200.990 65.380 ;
      LAYER via ;
        RECT 944.940 496.780 945.200 497.040 ;
        RECT 948.620 496.780 948.880 497.040 ;
        RECT 948.620 65.320 948.880 65.580 ;
        RECT 1200.700 65.320 1200.960 65.580 ;
      LAYER met2 ;
        RECT 945.070 510.340 945.350 514.000 ;
        RECT 945.000 510.000 945.350 510.340 ;
        RECT 945.000 497.070 945.140 510.000 ;
        RECT 944.940 496.750 945.200 497.070 ;
        RECT 948.620 496.750 948.880 497.070 ;
        RECT 948.680 65.610 948.820 496.750 ;
        RECT 948.620 65.290 948.880 65.610 ;
        RECT 1200.700 65.290 1200.960 65.610 ;
        RECT 1200.760 17.410 1200.900 65.290 ;
        RECT 1200.760 17.270 1204.120 17.410 ;
        RECT 1203.980 2.400 1204.120 17.270 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 961.470 496.980 961.790 497.040 ;
        RECT 965.610 496.980 965.930 497.040 ;
        RECT 961.470 496.840 965.930 496.980 ;
        RECT 961.470 496.780 961.790 496.840 ;
        RECT 965.610 496.780 965.930 496.840 ;
        RECT 965.610 72.320 965.930 72.380 ;
        RECT 1221.830 72.320 1222.150 72.380 ;
        RECT 965.610 72.180 1222.150 72.320 ;
        RECT 965.610 72.120 965.930 72.180 ;
        RECT 1221.830 72.120 1222.150 72.180 ;
      LAYER via ;
        RECT 961.500 496.780 961.760 497.040 ;
        RECT 965.640 496.780 965.900 497.040 ;
        RECT 965.640 72.120 965.900 72.380 ;
        RECT 1221.860 72.120 1222.120 72.380 ;
      LAYER met2 ;
        RECT 961.630 510.340 961.910 514.000 ;
        RECT 961.560 510.000 961.910 510.340 ;
        RECT 961.560 497.070 961.700 510.000 ;
        RECT 961.500 496.750 961.760 497.070 ;
        RECT 965.640 496.750 965.900 497.070 ;
        RECT 965.700 72.410 965.840 496.750 ;
        RECT 965.640 72.090 965.900 72.410 ;
        RECT 1221.860 72.090 1222.120 72.410 ;
        RECT 1221.920 2.400 1222.060 72.090 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.410 79.460 979.730 79.520 ;
        RECT 1235.170 79.460 1235.490 79.520 ;
        RECT 979.410 79.320 1235.490 79.460 ;
        RECT 979.410 79.260 979.730 79.320 ;
        RECT 1235.170 79.260 1235.490 79.320 ;
      LAYER via ;
        RECT 979.440 79.260 979.700 79.520 ;
        RECT 1235.200 79.260 1235.460 79.520 ;
      LAYER met2 ;
        RECT 977.730 510.410 978.010 514.000 ;
        RECT 977.730 510.270 979.640 510.410 ;
        RECT 977.730 510.000 978.010 510.270 ;
        RECT 979.500 79.550 979.640 510.270 ;
        RECT 979.440 79.230 979.700 79.550 ;
        RECT 1235.200 79.230 1235.460 79.550 ;
        RECT 1235.260 17.410 1235.400 79.230 ;
        RECT 1235.260 17.270 1240.000 17.410 ;
        RECT 1239.860 2.400 1240.000 17.270 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 994.130 493.240 994.450 493.300 ;
        RECT 1255.870 493.240 1256.190 493.300 ;
        RECT 994.130 493.100 1256.190 493.240 ;
        RECT 994.130 493.040 994.450 493.100 ;
        RECT 1255.870 493.040 1256.190 493.100 ;
      LAYER via ;
        RECT 994.160 493.040 994.420 493.300 ;
        RECT 1255.900 493.040 1256.160 493.300 ;
      LAYER met2 ;
        RECT 994.290 510.340 994.570 514.000 ;
        RECT 994.220 510.000 994.570 510.340 ;
        RECT 994.220 493.330 994.360 510.000 ;
        RECT 994.160 493.010 994.420 493.330 ;
        RECT 1255.900 493.010 1256.160 493.330 ;
        RECT 1255.960 17.410 1256.100 493.010 ;
        RECT 1255.960 17.270 1257.480 17.410 ;
        RECT 1257.340 2.400 1257.480 17.270 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1010.230 496.980 1010.550 497.040 ;
        RECT 1013.910 496.980 1014.230 497.040 ;
        RECT 1010.230 496.840 1014.230 496.980 ;
        RECT 1010.230 496.780 1010.550 496.840 ;
        RECT 1013.910 496.780 1014.230 496.840 ;
        RECT 1013.910 120.940 1014.230 121.000 ;
        RECT 1269.670 120.940 1269.990 121.000 ;
        RECT 1013.910 120.800 1269.990 120.940 ;
        RECT 1013.910 120.740 1014.230 120.800 ;
        RECT 1269.670 120.740 1269.990 120.800 ;
      LAYER via ;
        RECT 1010.260 496.780 1010.520 497.040 ;
        RECT 1013.940 496.780 1014.200 497.040 ;
        RECT 1013.940 120.740 1014.200 121.000 ;
        RECT 1269.700 120.740 1269.960 121.000 ;
      LAYER met2 ;
        RECT 1010.390 510.340 1010.670 514.000 ;
        RECT 1010.320 510.000 1010.670 510.340 ;
        RECT 1010.320 497.070 1010.460 510.000 ;
        RECT 1010.260 496.750 1010.520 497.070 ;
        RECT 1013.940 496.750 1014.200 497.070 ;
        RECT 1014.000 121.030 1014.140 496.750 ;
        RECT 1013.940 120.710 1014.200 121.030 ;
        RECT 1269.700 120.710 1269.960 121.030 ;
        RECT 1269.760 17.410 1269.900 120.710 ;
        RECT 1269.760 17.270 1275.420 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 99.860 1028.030 99.920 ;
        RECT 1290.370 99.860 1290.690 99.920 ;
        RECT 1027.710 99.720 1290.690 99.860 ;
        RECT 1027.710 99.660 1028.030 99.720 ;
        RECT 1290.370 99.660 1290.690 99.720 ;
      LAYER via ;
        RECT 1027.740 99.660 1028.000 99.920 ;
        RECT 1290.400 99.660 1290.660 99.920 ;
      LAYER met2 ;
        RECT 1026.950 510.410 1027.230 514.000 ;
        RECT 1026.950 510.270 1027.940 510.410 ;
        RECT 1026.950 510.000 1027.230 510.270 ;
        RECT 1027.800 99.950 1027.940 510.270 ;
        RECT 1027.740 99.630 1028.000 99.950 ;
        RECT 1290.400 99.630 1290.660 99.950 ;
        RECT 1290.460 17.410 1290.600 99.630 ;
        RECT 1290.460 17.270 1293.360 17.410 ;
        RECT 1293.220 2.400 1293.360 17.270 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1042.890 496.980 1043.210 497.040 ;
        RECT 1048.410 496.980 1048.730 497.040 ;
        RECT 1042.890 496.840 1048.730 496.980 ;
        RECT 1042.890 496.780 1043.210 496.840 ;
        RECT 1048.410 496.780 1048.730 496.840 ;
        RECT 1048.410 86.260 1048.730 86.320 ;
        RECT 1311.530 86.260 1311.850 86.320 ;
        RECT 1048.410 86.120 1311.850 86.260 ;
        RECT 1048.410 86.060 1048.730 86.120 ;
        RECT 1311.530 86.060 1311.850 86.120 ;
      LAYER via ;
        RECT 1042.920 496.780 1043.180 497.040 ;
        RECT 1048.440 496.780 1048.700 497.040 ;
        RECT 1048.440 86.060 1048.700 86.320 ;
        RECT 1311.560 86.060 1311.820 86.320 ;
      LAYER met2 ;
        RECT 1043.050 510.340 1043.330 514.000 ;
        RECT 1042.980 510.000 1043.330 510.340 ;
        RECT 1042.980 497.070 1043.120 510.000 ;
        RECT 1042.920 496.750 1043.180 497.070 ;
        RECT 1048.440 496.750 1048.700 497.070 ;
        RECT 1048.500 86.350 1048.640 496.750 ;
        RECT 1048.440 86.030 1048.700 86.350 ;
        RECT 1311.560 86.030 1311.820 86.350 ;
        RECT 1311.620 17.410 1311.760 86.030 ;
        RECT 1311.160 17.270 1311.760 17.410 ;
        RECT 1311.160 2.400 1311.300 17.270 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1059.450 500.380 1059.770 500.440 ;
        RECT 1155.590 500.380 1155.910 500.440 ;
        RECT 1059.450 500.240 1155.910 500.380 ;
        RECT 1059.450 500.180 1059.770 500.240 ;
        RECT 1155.590 500.180 1155.910 500.240 ;
        RECT 1155.590 24.380 1155.910 24.440 ;
        RECT 1329.010 24.380 1329.330 24.440 ;
        RECT 1155.590 24.240 1329.330 24.380 ;
        RECT 1155.590 24.180 1155.910 24.240 ;
        RECT 1329.010 24.180 1329.330 24.240 ;
      LAYER via ;
        RECT 1059.480 500.180 1059.740 500.440 ;
        RECT 1155.620 500.180 1155.880 500.440 ;
        RECT 1155.620 24.180 1155.880 24.440 ;
        RECT 1329.040 24.180 1329.300 24.440 ;
      LAYER met2 ;
        RECT 1059.610 510.340 1059.890 514.000 ;
        RECT 1059.540 510.000 1059.890 510.340 ;
        RECT 1059.540 500.470 1059.680 510.000 ;
        RECT 1059.480 500.150 1059.740 500.470 ;
        RECT 1155.620 500.150 1155.880 500.470 ;
        RECT 1155.680 24.470 1155.820 500.150 ;
        RECT 1155.620 24.150 1155.880 24.470 ;
        RECT 1329.040 24.150 1329.300 24.470 ;
        RECT 1329.100 2.400 1329.240 24.150 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.030 503.440 472.350 503.500 ;
        RECT 475.710 503.440 476.030 503.500 ;
        RECT 472.030 503.300 476.030 503.440 ;
        RECT 472.030 503.240 472.350 503.300 ;
        RECT 475.710 503.240 476.030 503.300 ;
        RECT 475.710 51.580 476.030 51.640 ;
        RECT 683.170 51.580 683.490 51.640 ;
        RECT 475.710 51.440 683.490 51.580 ;
        RECT 475.710 51.380 476.030 51.440 ;
        RECT 683.170 51.380 683.490 51.440 ;
      LAYER via ;
        RECT 472.060 503.240 472.320 503.500 ;
        RECT 475.740 503.240 476.000 503.500 ;
        RECT 475.740 51.380 476.000 51.640 ;
        RECT 683.200 51.380 683.460 51.640 ;
      LAYER met2 ;
        RECT 472.190 510.340 472.470 514.000 ;
        RECT 472.120 510.000 472.470 510.340 ;
        RECT 472.120 503.530 472.260 510.000 ;
        RECT 472.060 503.210 472.320 503.530 ;
        RECT 475.740 503.210 476.000 503.530 ;
        RECT 475.800 51.670 475.940 503.210 ;
        RECT 475.740 51.350 476.000 51.670 ;
        RECT 683.200 51.350 683.460 51.670 ;
        RECT 683.260 17.410 683.400 51.350 ;
        RECT 683.260 17.270 686.620 17.410 ;
        RECT 686.480 2.400 686.620 17.270 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 196.760 1076.330 196.820 ;
        RECT 1345.570 196.760 1345.890 196.820 ;
        RECT 1076.010 196.620 1345.890 196.760 ;
        RECT 1076.010 196.560 1076.330 196.620 ;
        RECT 1345.570 196.560 1345.890 196.620 ;
      LAYER via ;
        RECT 1076.040 196.560 1076.300 196.820 ;
        RECT 1345.600 196.560 1345.860 196.820 ;
      LAYER met2 ;
        RECT 1075.710 510.340 1075.990 514.000 ;
        RECT 1075.640 510.000 1075.990 510.340 ;
        RECT 1075.640 497.490 1075.780 510.000 ;
        RECT 1075.640 497.350 1076.240 497.490 ;
        RECT 1076.100 196.850 1076.240 497.350 ;
        RECT 1076.040 196.530 1076.300 196.850 ;
        RECT 1345.600 196.530 1345.860 196.850 ;
        RECT 1345.660 17.410 1345.800 196.530 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1092.110 496.980 1092.430 497.040 ;
        RECT 1096.710 496.980 1097.030 497.040 ;
        RECT 1092.110 496.840 1097.030 496.980 ;
        RECT 1092.110 496.780 1092.430 496.840 ;
        RECT 1096.710 496.780 1097.030 496.840 ;
        RECT 1096.710 30.840 1097.030 30.900 ;
        RECT 1364.430 30.840 1364.750 30.900 ;
        RECT 1096.710 30.700 1364.750 30.840 ;
        RECT 1096.710 30.640 1097.030 30.700 ;
        RECT 1364.430 30.640 1364.750 30.700 ;
      LAYER via ;
        RECT 1092.140 496.780 1092.400 497.040 ;
        RECT 1096.740 496.780 1097.000 497.040 ;
        RECT 1096.740 30.640 1097.000 30.900 ;
        RECT 1364.460 30.640 1364.720 30.900 ;
      LAYER met2 ;
        RECT 1092.270 510.340 1092.550 514.000 ;
        RECT 1092.200 510.000 1092.550 510.340 ;
        RECT 1092.200 497.070 1092.340 510.000 ;
        RECT 1092.140 496.750 1092.400 497.070 ;
        RECT 1096.740 496.750 1097.000 497.070 ;
        RECT 1096.800 30.930 1096.940 496.750 ;
        RECT 1096.740 30.610 1097.000 30.930 ;
        RECT 1364.460 30.610 1364.720 30.930 ;
        RECT 1364.520 2.400 1364.660 30.610 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 93.060 1110.830 93.120 ;
        RECT 1380.070 93.060 1380.390 93.120 ;
        RECT 1110.510 92.920 1380.390 93.060 ;
        RECT 1110.510 92.860 1110.830 92.920 ;
        RECT 1380.070 92.860 1380.390 92.920 ;
      LAYER via ;
        RECT 1110.540 92.860 1110.800 93.120 ;
        RECT 1380.100 92.860 1380.360 93.120 ;
      LAYER met2 ;
        RECT 1108.370 510.410 1108.650 514.000 ;
        RECT 1108.370 510.270 1110.740 510.410 ;
        RECT 1108.370 510.000 1108.650 510.270 ;
        RECT 1110.600 93.150 1110.740 510.270 ;
        RECT 1110.540 92.830 1110.800 93.150 ;
        RECT 1380.100 92.830 1380.360 93.150 ;
        RECT 1380.160 17.410 1380.300 92.830 ;
        RECT 1380.160 17.270 1382.600 17.410 ;
        RECT 1382.460 2.400 1382.600 17.270 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1124.770 499.020 1125.090 499.080 ;
        RECT 1131.210 499.020 1131.530 499.080 ;
        RECT 1124.770 498.880 1131.530 499.020 ;
        RECT 1124.770 498.820 1125.090 498.880 ;
        RECT 1131.210 498.820 1131.530 498.880 ;
        RECT 1131.210 107.340 1131.530 107.400 ;
        RECT 1394.330 107.340 1394.650 107.400 ;
        RECT 1131.210 107.200 1394.650 107.340 ;
        RECT 1131.210 107.140 1131.530 107.200 ;
        RECT 1394.330 107.140 1394.650 107.200 ;
        RECT 1394.330 17.920 1394.650 17.980 ;
        RECT 1400.310 17.920 1400.630 17.980 ;
        RECT 1394.330 17.780 1400.630 17.920 ;
        RECT 1394.330 17.720 1394.650 17.780 ;
        RECT 1400.310 17.720 1400.630 17.780 ;
      LAYER via ;
        RECT 1124.800 498.820 1125.060 499.080 ;
        RECT 1131.240 498.820 1131.500 499.080 ;
        RECT 1131.240 107.140 1131.500 107.400 ;
        RECT 1394.360 107.140 1394.620 107.400 ;
        RECT 1394.360 17.720 1394.620 17.980 ;
        RECT 1400.340 17.720 1400.600 17.980 ;
      LAYER met2 ;
        RECT 1124.930 510.340 1125.210 514.000 ;
        RECT 1124.860 510.000 1125.210 510.340 ;
        RECT 1124.860 499.110 1125.000 510.000 ;
        RECT 1124.800 498.790 1125.060 499.110 ;
        RECT 1131.240 498.790 1131.500 499.110 ;
        RECT 1131.300 107.430 1131.440 498.790 ;
        RECT 1131.240 107.110 1131.500 107.430 ;
        RECT 1394.360 107.110 1394.620 107.430 ;
        RECT 1394.420 18.010 1394.560 107.110 ;
        RECT 1394.360 17.690 1394.620 18.010 ;
        RECT 1400.340 17.690 1400.600 18.010 ;
        RECT 1400.400 2.400 1400.540 17.690 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1140.870 503.440 1141.190 503.500 ;
        RECT 1145.010 503.440 1145.330 503.500 ;
        RECT 1140.870 503.300 1145.330 503.440 ;
        RECT 1140.870 503.240 1141.190 503.300 ;
        RECT 1145.010 503.240 1145.330 503.300 ;
        RECT 1145.010 210.360 1145.330 210.420 ;
        RECT 1414.570 210.360 1414.890 210.420 ;
        RECT 1145.010 210.220 1414.890 210.360 ;
        RECT 1145.010 210.160 1145.330 210.220 ;
        RECT 1414.570 210.160 1414.890 210.220 ;
      LAYER via ;
        RECT 1140.900 503.240 1141.160 503.500 ;
        RECT 1145.040 503.240 1145.300 503.500 ;
        RECT 1145.040 210.160 1145.300 210.420 ;
        RECT 1414.600 210.160 1414.860 210.420 ;
      LAYER met2 ;
        RECT 1141.030 510.340 1141.310 514.000 ;
        RECT 1140.960 510.000 1141.310 510.340 ;
        RECT 1140.960 503.530 1141.100 510.000 ;
        RECT 1140.900 503.210 1141.160 503.530 ;
        RECT 1145.040 503.210 1145.300 503.530 ;
        RECT 1145.100 210.450 1145.240 503.210 ;
        RECT 1145.040 210.130 1145.300 210.450 ;
        RECT 1414.600 210.130 1414.860 210.450 ;
        RECT 1414.660 17.410 1414.800 210.130 ;
        RECT 1414.660 17.270 1418.480 17.410 ;
        RECT 1418.340 2.400 1418.480 17.270 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1157.430 500.040 1157.750 500.100 ;
        RECT 1436.190 500.040 1436.510 500.100 ;
        RECT 1157.430 499.900 1436.510 500.040 ;
        RECT 1157.430 499.840 1157.750 499.900 ;
        RECT 1436.190 499.840 1436.510 499.900 ;
      LAYER via ;
        RECT 1157.460 499.840 1157.720 500.100 ;
        RECT 1436.220 499.840 1436.480 500.100 ;
      LAYER met2 ;
        RECT 1157.590 510.340 1157.870 514.000 ;
        RECT 1157.520 510.000 1157.870 510.340 ;
        RECT 1157.520 500.130 1157.660 510.000 ;
        RECT 1157.460 499.810 1157.720 500.130 ;
        RECT 1436.220 499.810 1436.480 500.130 ;
        RECT 1436.280 7.210 1436.420 499.810 ;
        RECT 1435.820 7.070 1436.420 7.210 ;
        RECT 1435.820 2.400 1435.960 7.070 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.530 486.440 1173.850 486.500 ;
        RECT 1449.070 486.440 1449.390 486.500 ;
        RECT 1173.530 486.300 1449.390 486.440 ;
        RECT 1173.530 486.240 1173.850 486.300 ;
        RECT 1449.070 486.240 1449.390 486.300 ;
      LAYER via ;
        RECT 1173.560 486.240 1173.820 486.500 ;
        RECT 1449.100 486.240 1449.360 486.500 ;
      LAYER met2 ;
        RECT 1173.690 510.340 1173.970 514.000 ;
        RECT 1173.620 510.000 1173.970 510.340 ;
        RECT 1173.620 486.530 1173.760 510.000 ;
        RECT 1173.560 486.210 1173.820 486.530 ;
        RECT 1449.100 486.210 1449.360 486.530 ;
        RECT 1449.160 17.410 1449.300 486.210 ;
        RECT 1449.160 17.270 1453.900 17.410 ;
        RECT 1453.760 2.400 1453.900 17.270 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.310 37.980 1193.630 38.040 ;
        RECT 1471.610 37.980 1471.930 38.040 ;
        RECT 1193.310 37.840 1471.930 37.980 ;
        RECT 1193.310 37.780 1193.630 37.840 ;
        RECT 1471.610 37.780 1471.930 37.840 ;
      LAYER via ;
        RECT 1193.340 37.780 1193.600 38.040 ;
        RECT 1471.640 37.780 1471.900 38.040 ;
      LAYER met2 ;
        RECT 1190.250 510.410 1190.530 514.000 ;
        RECT 1190.250 510.270 1193.540 510.410 ;
        RECT 1190.250 510.000 1190.530 510.270 ;
        RECT 1193.400 38.070 1193.540 510.270 ;
        RECT 1193.340 37.750 1193.600 38.070 ;
        RECT 1471.640 37.750 1471.900 38.070 ;
        RECT 1471.700 2.400 1471.840 37.750 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 58.720 1207.430 58.780 ;
        RECT 1484.030 58.720 1484.350 58.780 ;
        RECT 1207.110 58.580 1484.350 58.720 ;
        RECT 1207.110 58.520 1207.430 58.580 ;
        RECT 1484.030 58.520 1484.350 58.580 ;
      LAYER via ;
        RECT 1207.140 58.520 1207.400 58.780 ;
        RECT 1484.060 58.520 1484.320 58.780 ;
      LAYER met2 ;
        RECT 1206.350 510.410 1206.630 514.000 ;
        RECT 1206.350 510.270 1207.340 510.410 ;
        RECT 1206.350 510.000 1206.630 510.270 ;
        RECT 1207.200 58.810 1207.340 510.270 ;
        RECT 1207.140 58.490 1207.400 58.810 ;
        RECT 1484.060 58.490 1484.320 58.810 ;
        RECT 1484.120 17.410 1484.260 58.490 ;
        RECT 1484.120 17.270 1489.780 17.410 ;
        RECT 1489.640 2.400 1489.780 17.270 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1222.750 496.980 1223.070 497.040 ;
        RECT 1227.810 496.980 1228.130 497.040 ;
        RECT 1222.750 496.840 1228.130 496.980 ;
        RECT 1222.750 496.780 1223.070 496.840 ;
        RECT 1227.810 496.780 1228.130 496.840 ;
        RECT 1227.810 44.780 1228.130 44.840 ;
        RECT 1507.030 44.780 1507.350 44.840 ;
        RECT 1227.810 44.640 1507.350 44.780 ;
        RECT 1227.810 44.580 1228.130 44.640 ;
        RECT 1507.030 44.580 1507.350 44.640 ;
      LAYER via ;
        RECT 1222.780 496.780 1223.040 497.040 ;
        RECT 1227.840 496.780 1228.100 497.040 ;
        RECT 1227.840 44.580 1228.100 44.840 ;
        RECT 1507.060 44.580 1507.320 44.840 ;
      LAYER met2 ;
        RECT 1222.910 510.340 1223.190 514.000 ;
        RECT 1222.840 510.000 1223.190 510.340 ;
        RECT 1222.840 497.070 1222.980 510.000 ;
        RECT 1222.780 496.750 1223.040 497.070 ;
        RECT 1227.840 496.750 1228.100 497.070 ;
        RECT 1227.900 44.870 1228.040 496.750 ;
        RECT 1227.840 44.550 1228.100 44.870 ;
        RECT 1507.060 44.550 1507.320 44.870 ;
        RECT 1507.120 2.400 1507.260 44.550 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.510 72.320 489.830 72.380 ;
        RECT 704.330 72.320 704.650 72.380 ;
        RECT 489.510 72.180 704.650 72.320 ;
        RECT 489.510 72.120 489.830 72.180 ;
        RECT 704.330 72.120 704.650 72.180 ;
      LAYER via ;
        RECT 489.540 72.120 489.800 72.380 ;
        RECT 704.360 72.120 704.620 72.380 ;
      LAYER met2 ;
        RECT 488.290 510.410 488.570 514.000 ;
        RECT 488.290 510.270 489.740 510.410 ;
        RECT 488.290 510.000 488.570 510.270 ;
        RECT 489.600 72.410 489.740 510.270 ;
        RECT 489.540 72.090 489.800 72.410 ;
        RECT 704.360 72.090 704.620 72.410 ;
        RECT 704.420 2.400 704.560 72.090 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 51.580 1241.930 51.640 ;
        RECT 1525.430 51.580 1525.750 51.640 ;
        RECT 1241.610 51.440 1525.750 51.580 ;
        RECT 1241.610 51.380 1241.930 51.440 ;
        RECT 1525.430 51.380 1525.750 51.440 ;
      LAYER via ;
        RECT 1241.640 51.380 1241.900 51.640 ;
        RECT 1525.460 51.380 1525.720 51.640 ;
      LAYER met2 ;
        RECT 1239.010 510.410 1239.290 514.000 ;
        RECT 1239.010 510.270 1241.840 510.410 ;
        RECT 1239.010 510.000 1239.290 510.270 ;
        RECT 1241.700 51.670 1241.840 510.270 ;
        RECT 1241.640 51.350 1241.900 51.670 ;
        RECT 1525.460 51.350 1525.720 51.670 ;
        RECT 1525.520 7.210 1525.660 51.350 ;
        RECT 1525.060 7.070 1525.660 7.210 ;
        RECT 1525.060 2.400 1525.200 7.070 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 182.820 1255.730 182.880 ;
        RECT 1538.770 182.820 1539.090 182.880 ;
        RECT 1255.410 182.680 1539.090 182.820 ;
        RECT 1255.410 182.620 1255.730 182.680 ;
        RECT 1538.770 182.620 1539.090 182.680 ;
      LAYER via ;
        RECT 1255.440 182.620 1255.700 182.880 ;
        RECT 1538.800 182.620 1539.060 182.880 ;
      LAYER met2 ;
        RECT 1255.570 510.340 1255.850 514.000 ;
        RECT 1255.500 510.000 1255.850 510.340 ;
        RECT 1255.500 182.910 1255.640 510.000 ;
        RECT 1255.440 182.590 1255.700 182.910 ;
        RECT 1538.800 182.590 1539.060 182.910 ;
        RECT 1538.860 17.410 1539.000 182.590 ;
        RECT 1538.860 17.270 1543.140 17.410 ;
        RECT 1543.000 2.400 1543.140 17.270 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1271.510 496.980 1271.830 497.040 ;
        RECT 1276.110 496.980 1276.430 497.040 ;
        RECT 1271.510 496.840 1276.430 496.980 ;
        RECT 1271.510 496.780 1271.830 496.840 ;
        RECT 1276.110 496.780 1276.430 496.840 ;
        RECT 1276.110 65.520 1276.430 65.580 ;
        RECT 1559.470 65.520 1559.790 65.580 ;
        RECT 1276.110 65.380 1559.790 65.520 ;
        RECT 1276.110 65.320 1276.430 65.380 ;
        RECT 1559.470 65.320 1559.790 65.380 ;
      LAYER via ;
        RECT 1271.540 496.780 1271.800 497.040 ;
        RECT 1276.140 496.780 1276.400 497.040 ;
        RECT 1276.140 65.320 1276.400 65.580 ;
        RECT 1559.500 65.320 1559.760 65.580 ;
      LAYER met2 ;
        RECT 1271.670 510.340 1271.950 514.000 ;
        RECT 1271.600 510.000 1271.950 510.340 ;
        RECT 1271.600 497.070 1271.740 510.000 ;
        RECT 1271.540 496.750 1271.800 497.070 ;
        RECT 1276.140 496.750 1276.400 497.070 ;
        RECT 1276.200 65.610 1276.340 496.750 ;
        RECT 1276.140 65.290 1276.400 65.610 ;
        RECT 1559.500 65.290 1559.760 65.610 ;
        RECT 1559.560 17.410 1559.700 65.290 ;
        RECT 1559.560 17.270 1561.080 17.410 ;
        RECT 1560.940 2.400 1561.080 17.270 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 72.320 1290.230 72.380 ;
        RECT 1573.270 72.320 1573.590 72.380 ;
        RECT 1289.910 72.180 1573.590 72.320 ;
        RECT 1289.910 72.120 1290.230 72.180 ;
        RECT 1573.270 72.120 1573.590 72.180 ;
      LAYER via ;
        RECT 1289.940 72.120 1290.200 72.380 ;
        RECT 1573.300 72.120 1573.560 72.380 ;
      LAYER met2 ;
        RECT 1288.230 510.410 1288.510 514.000 ;
        RECT 1288.230 510.270 1290.140 510.410 ;
        RECT 1288.230 510.000 1288.510 510.270 ;
        RECT 1290.000 72.410 1290.140 510.270 ;
        RECT 1289.940 72.090 1290.200 72.410 ;
        RECT 1573.300 72.090 1573.560 72.410 ;
        RECT 1573.360 17.410 1573.500 72.090 ;
        RECT 1573.360 17.270 1579.020 17.410 ;
        RECT 1578.880 2.400 1579.020 17.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 496.980 1304.490 497.040 ;
        RECT 1310.150 496.980 1310.470 497.040 ;
        RECT 1304.170 496.840 1310.470 496.980 ;
        RECT 1304.170 496.780 1304.490 496.840 ;
        RECT 1310.150 496.780 1310.470 496.840 ;
        RECT 1310.150 224.300 1310.470 224.360 ;
        RECT 1593.970 224.300 1594.290 224.360 ;
        RECT 1310.150 224.160 1594.290 224.300 ;
        RECT 1310.150 224.100 1310.470 224.160 ;
        RECT 1593.970 224.100 1594.290 224.160 ;
      LAYER via ;
        RECT 1304.200 496.780 1304.460 497.040 ;
        RECT 1310.180 496.780 1310.440 497.040 ;
        RECT 1310.180 224.100 1310.440 224.360 ;
        RECT 1594.000 224.100 1594.260 224.360 ;
      LAYER met2 ;
        RECT 1304.330 510.340 1304.610 514.000 ;
        RECT 1304.260 510.000 1304.610 510.340 ;
        RECT 1304.260 497.070 1304.400 510.000 ;
        RECT 1304.200 496.750 1304.460 497.070 ;
        RECT 1310.180 496.750 1310.440 497.070 ;
        RECT 1310.240 224.390 1310.380 496.750 ;
        RECT 1310.180 224.070 1310.440 224.390 ;
        RECT 1594.000 224.070 1594.260 224.390 ;
        RECT 1594.060 16.730 1594.200 224.070 ;
        RECT 1594.060 16.590 1596.500 16.730 ;
        RECT 1596.360 2.400 1596.500 16.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 24.040 1324.730 24.100 ;
        RECT 1614.210 24.040 1614.530 24.100 ;
        RECT 1324.410 23.900 1614.530 24.040 ;
        RECT 1324.410 23.840 1324.730 23.900 ;
        RECT 1614.210 23.840 1614.530 23.900 ;
      LAYER via ;
        RECT 1324.440 23.840 1324.700 24.100 ;
        RECT 1614.240 23.840 1614.500 24.100 ;
      LAYER met2 ;
        RECT 1320.890 510.410 1321.170 514.000 ;
        RECT 1320.890 510.270 1324.640 510.410 ;
        RECT 1320.890 510.000 1321.170 510.270 ;
        RECT 1324.500 24.130 1324.640 510.270 ;
        RECT 1324.440 23.810 1324.700 24.130 ;
        RECT 1614.240 23.810 1614.500 24.130 ;
        RECT 1614.300 2.400 1614.440 23.810 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 79.460 1338.530 79.520 ;
        RECT 1628.470 79.460 1628.790 79.520 ;
        RECT 1338.210 79.320 1628.790 79.460 ;
        RECT 1338.210 79.260 1338.530 79.320 ;
        RECT 1628.470 79.260 1628.790 79.320 ;
      LAYER via ;
        RECT 1338.240 79.260 1338.500 79.520 ;
        RECT 1628.500 79.260 1628.760 79.520 ;
      LAYER met2 ;
        RECT 1336.990 510.410 1337.270 514.000 ;
        RECT 1336.990 510.270 1338.440 510.410 ;
        RECT 1336.990 510.000 1337.270 510.270 ;
        RECT 1338.300 79.550 1338.440 510.270 ;
        RECT 1338.240 79.230 1338.500 79.550 ;
        RECT 1628.500 79.230 1628.760 79.550 ;
        RECT 1628.560 17.410 1628.700 79.230 ;
        RECT 1628.560 17.270 1632.380 17.410 ;
        RECT 1632.240 2.400 1632.380 17.270 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.930 493.240 1353.250 493.300 ;
        RECT 1649.170 493.240 1649.490 493.300 ;
        RECT 1352.930 493.100 1649.490 493.240 ;
        RECT 1352.930 493.040 1353.250 493.100 ;
        RECT 1649.170 493.040 1649.490 493.100 ;
      LAYER via ;
        RECT 1352.960 493.040 1353.220 493.300 ;
        RECT 1649.200 493.040 1649.460 493.300 ;
      LAYER met2 ;
        RECT 1353.090 510.340 1353.370 514.000 ;
        RECT 1353.020 510.000 1353.370 510.340 ;
        RECT 1353.020 493.330 1353.160 510.000 ;
        RECT 1352.960 493.010 1353.220 493.330 ;
        RECT 1649.200 493.010 1649.460 493.330 ;
        RECT 1649.260 17.410 1649.400 493.010 ;
        RECT 1649.260 17.270 1650.320 17.410 ;
        RECT 1650.180 2.400 1650.320 17.270 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.710 30.840 1373.030 30.900 ;
        RECT 1668.030 30.840 1668.350 30.900 ;
        RECT 1372.710 30.700 1668.350 30.840 ;
        RECT 1372.710 30.640 1373.030 30.700 ;
        RECT 1668.030 30.640 1668.350 30.700 ;
      LAYER via ;
        RECT 1372.740 30.640 1373.000 30.900 ;
        RECT 1668.060 30.640 1668.320 30.900 ;
      LAYER met2 ;
        RECT 1369.650 510.410 1369.930 514.000 ;
        RECT 1369.650 510.270 1372.940 510.410 ;
        RECT 1369.650 510.000 1369.930 510.270 ;
        RECT 1372.800 30.930 1372.940 510.270 ;
        RECT 1372.740 30.610 1373.000 30.930 ;
        RECT 1668.060 30.610 1668.320 30.930 ;
        RECT 1668.120 2.400 1668.260 30.610 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 168.880 1386.830 168.940 ;
        RECT 1683.670 168.880 1683.990 168.940 ;
        RECT 1386.510 168.740 1683.990 168.880 ;
        RECT 1386.510 168.680 1386.830 168.740 ;
        RECT 1683.670 168.680 1683.990 168.740 ;
      LAYER via ;
        RECT 1386.540 168.680 1386.800 168.940 ;
        RECT 1683.700 168.680 1683.960 168.940 ;
      LAYER met2 ;
        RECT 1385.750 510.410 1386.030 514.000 ;
        RECT 1385.750 510.270 1386.740 510.410 ;
        RECT 1385.750 510.000 1386.030 510.270 ;
        RECT 1386.600 168.970 1386.740 510.270 ;
        RECT 1386.540 168.650 1386.800 168.970 ;
        RECT 1683.700 168.650 1683.960 168.970 ;
        RECT 1683.760 17.410 1683.900 168.650 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 504.690 503.440 505.010 503.500 ;
        RECT 513.890 503.440 514.210 503.500 ;
        RECT 504.690 503.300 514.210 503.440 ;
        RECT 504.690 503.240 505.010 503.300 ;
        RECT 513.890 503.240 514.210 503.300 ;
        RECT 513.890 79.460 514.210 79.520 ;
        RECT 717.670 79.460 717.990 79.520 ;
        RECT 513.890 79.320 717.990 79.460 ;
        RECT 513.890 79.260 514.210 79.320 ;
        RECT 717.670 79.260 717.990 79.320 ;
      LAYER via ;
        RECT 504.720 503.240 504.980 503.500 ;
        RECT 513.920 503.240 514.180 503.500 ;
        RECT 513.920 79.260 514.180 79.520 ;
        RECT 717.700 79.260 717.960 79.520 ;
      LAYER met2 ;
        RECT 504.850 510.340 505.130 514.000 ;
        RECT 504.780 510.000 505.130 510.340 ;
        RECT 504.780 503.530 504.920 510.000 ;
        RECT 504.720 503.210 504.980 503.530 ;
        RECT 513.920 503.210 514.180 503.530 ;
        RECT 513.980 79.550 514.120 503.210 ;
        RECT 513.920 79.230 514.180 79.550 ;
        RECT 717.700 79.230 717.960 79.550 ;
        RECT 717.760 17.410 717.900 79.230 ;
        RECT 717.760 17.270 722.500 17.410 ;
        RECT 722.360 2.400 722.500 17.270 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1402.150 496.980 1402.470 497.040 ;
        RECT 1407.210 496.980 1407.530 497.040 ;
        RECT 1402.150 496.840 1407.530 496.980 ;
        RECT 1402.150 496.780 1402.470 496.840 ;
        RECT 1407.210 496.780 1407.530 496.840 ;
        RECT 1407.210 86.600 1407.530 86.660 ;
        RECT 1697.930 86.600 1698.250 86.660 ;
        RECT 1407.210 86.460 1698.250 86.600 ;
        RECT 1407.210 86.400 1407.530 86.460 ;
        RECT 1697.930 86.400 1698.250 86.460 ;
      LAYER via ;
        RECT 1402.180 496.780 1402.440 497.040 ;
        RECT 1407.240 496.780 1407.500 497.040 ;
        RECT 1407.240 86.400 1407.500 86.660 ;
        RECT 1697.960 86.400 1698.220 86.660 ;
      LAYER met2 ;
        RECT 1402.310 510.340 1402.590 514.000 ;
        RECT 1402.240 510.000 1402.590 510.340 ;
        RECT 1402.240 497.070 1402.380 510.000 ;
        RECT 1402.180 496.750 1402.440 497.070 ;
        RECT 1407.240 496.750 1407.500 497.070 ;
        RECT 1407.300 86.690 1407.440 496.750 ;
        RECT 1407.240 86.370 1407.500 86.690 ;
        RECT 1697.960 86.370 1698.220 86.690 ;
        RECT 1698.020 17.410 1698.160 86.370 ;
        RECT 1698.020 17.270 1703.680 17.410 ;
        RECT 1703.540 2.400 1703.680 17.270 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 93.060 1421.330 93.120 ;
        RECT 1718.170 93.060 1718.490 93.120 ;
        RECT 1421.010 92.920 1718.490 93.060 ;
        RECT 1421.010 92.860 1421.330 92.920 ;
        RECT 1718.170 92.860 1718.490 92.920 ;
      LAYER via ;
        RECT 1421.040 92.860 1421.300 93.120 ;
        RECT 1718.200 92.860 1718.460 93.120 ;
      LAYER met2 ;
        RECT 1418.410 510.410 1418.690 514.000 ;
        RECT 1418.410 510.270 1421.240 510.410 ;
        RECT 1418.410 510.000 1418.690 510.270 ;
        RECT 1421.100 93.150 1421.240 510.270 ;
        RECT 1421.040 92.830 1421.300 93.150 ;
        RECT 1718.200 92.830 1718.460 93.150 ;
        RECT 1718.260 17.410 1718.400 92.830 ;
        RECT 1718.260 17.270 1721.620 17.410 ;
        RECT 1721.480 2.400 1721.620 17.270 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 500.380 1435.130 500.440 ;
        RECT 1617.890 500.380 1618.210 500.440 ;
        RECT 1434.810 500.240 1618.210 500.380 ;
        RECT 1434.810 500.180 1435.130 500.240 ;
        RECT 1617.890 500.180 1618.210 500.240 ;
        RECT 1617.890 24.040 1618.210 24.100 ;
        RECT 1739.330 24.040 1739.650 24.100 ;
        RECT 1617.890 23.900 1739.650 24.040 ;
        RECT 1617.890 23.840 1618.210 23.900 ;
        RECT 1739.330 23.840 1739.650 23.900 ;
      LAYER via ;
        RECT 1434.840 500.180 1435.100 500.440 ;
        RECT 1617.920 500.180 1618.180 500.440 ;
        RECT 1617.920 23.840 1618.180 24.100 ;
        RECT 1739.360 23.840 1739.620 24.100 ;
      LAYER met2 ;
        RECT 1434.970 510.340 1435.250 514.000 ;
        RECT 1434.900 510.000 1435.250 510.340 ;
        RECT 1434.900 500.470 1435.040 510.000 ;
        RECT 1434.840 500.150 1435.100 500.470 ;
        RECT 1617.920 500.150 1618.180 500.470 ;
        RECT 1617.980 24.130 1618.120 500.150 ;
        RECT 1617.920 23.810 1618.180 24.130 ;
        RECT 1739.360 23.810 1739.620 24.130 ;
        RECT 1739.420 2.400 1739.560 23.810 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1450.910 496.980 1451.230 497.040 ;
        RECT 1455.510 496.980 1455.830 497.040 ;
        RECT 1450.910 496.840 1455.830 496.980 ;
        RECT 1450.910 496.780 1451.230 496.840 ;
        RECT 1455.510 496.780 1455.830 496.840 ;
        RECT 1455.510 196.760 1455.830 196.820 ;
        RECT 1752.670 196.760 1752.990 196.820 ;
        RECT 1455.510 196.620 1752.990 196.760 ;
        RECT 1455.510 196.560 1455.830 196.620 ;
        RECT 1752.670 196.560 1752.990 196.620 ;
        RECT 1752.670 62.120 1752.990 62.180 ;
        RECT 1756.810 62.120 1757.130 62.180 ;
        RECT 1752.670 61.980 1757.130 62.120 ;
        RECT 1752.670 61.920 1752.990 61.980 ;
        RECT 1756.810 61.920 1757.130 61.980 ;
      LAYER via ;
        RECT 1450.940 496.780 1451.200 497.040 ;
        RECT 1455.540 496.780 1455.800 497.040 ;
        RECT 1455.540 196.560 1455.800 196.820 ;
        RECT 1752.700 196.560 1752.960 196.820 ;
        RECT 1752.700 61.920 1752.960 62.180 ;
        RECT 1756.840 61.920 1757.100 62.180 ;
      LAYER met2 ;
        RECT 1451.070 510.340 1451.350 514.000 ;
        RECT 1451.000 510.000 1451.350 510.340 ;
        RECT 1451.000 497.070 1451.140 510.000 ;
        RECT 1450.940 496.750 1451.200 497.070 ;
        RECT 1455.540 496.750 1455.800 497.070 ;
        RECT 1455.600 196.850 1455.740 496.750 ;
        RECT 1455.540 196.530 1455.800 196.850 ;
        RECT 1752.700 196.530 1752.960 196.850 ;
        RECT 1752.760 62.210 1752.900 196.530 ;
        RECT 1752.700 61.890 1752.960 62.210 ;
        RECT 1756.840 61.890 1757.100 62.210 ;
        RECT 1756.900 2.400 1757.040 61.890 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 99.860 1469.630 99.920 ;
        RECT 1773.370 99.860 1773.690 99.920 ;
        RECT 1469.310 99.720 1773.690 99.860 ;
        RECT 1469.310 99.660 1469.630 99.720 ;
        RECT 1773.370 99.660 1773.690 99.720 ;
        RECT 1773.370 62.260 1773.690 62.520 ;
        RECT 1773.460 61.780 1773.600 62.260 ;
        RECT 1774.750 61.780 1775.070 61.840 ;
        RECT 1773.460 61.640 1775.070 61.780 ;
        RECT 1774.750 61.580 1775.070 61.640 ;
        RECT 1774.750 47.980 1775.070 48.240 ;
        RECT 1774.840 47.560 1774.980 47.980 ;
        RECT 1774.750 47.300 1775.070 47.560 ;
      LAYER via ;
        RECT 1469.340 99.660 1469.600 99.920 ;
        RECT 1773.400 99.660 1773.660 99.920 ;
        RECT 1773.400 62.260 1773.660 62.520 ;
        RECT 1774.780 61.580 1775.040 61.840 ;
        RECT 1774.780 47.980 1775.040 48.240 ;
        RECT 1774.780 47.300 1775.040 47.560 ;
      LAYER met2 ;
        RECT 1467.630 510.410 1467.910 514.000 ;
        RECT 1467.630 510.270 1469.540 510.410 ;
        RECT 1467.630 510.000 1467.910 510.270 ;
        RECT 1469.400 99.950 1469.540 510.270 ;
        RECT 1469.340 99.630 1469.600 99.950 ;
        RECT 1773.400 99.630 1773.660 99.950 ;
        RECT 1773.460 62.550 1773.600 99.630 ;
        RECT 1773.400 62.230 1773.660 62.550 ;
        RECT 1774.780 61.550 1775.040 61.870 ;
        RECT 1774.840 48.270 1774.980 61.550 ;
        RECT 1774.780 47.950 1775.040 48.270 ;
        RECT 1774.780 47.270 1775.040 47.590 ;
        RECT 1774.840 2.400 1774.980 47.270 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.570 498.000 1483.890 498.060 ;
        RECT 1490.010 498.000 1490.330 498.060 ;
        RECT 1483.570 497.860 1490.330 498.000 ;
        RECT 1483.570 497.800 1483.890 497.860 ;
        RECT 1490.010 497.800 1490.330 497.860 ;
        RECT 1490.010 37.980 1490.330 38.040 ;
        RECT 1490.010 37.840 1772.680 37.980 ;
        RECT 1490.010 37.780 1490.330 37.840 ;
        RECT 1772.540 37.640 1772.680 37.840 ;
        RECT 1792.690 37.640 1793.010 37.700 ;
        RECT 1772.540 37.500 1793.010 37.640 ;
        RECT 1792.690 37.440 1793.010 37.500 ;
      LAYER via ;
        RECT 1483.600 497.800 1483.860 498.060 ;
        RECT 1490.040 497.800 1490.300 498.060 ;
        RECT 1490.040 37.780 1490.300 38.040 ;
        RECT 1792.720 37.440 1792.980 37.700 ;
      LAYER met2 ;
        RECT 1483.730 510.340 1484.010 514.000 ;
        RECT 1483.660 510.000 1484.010 510.340 ;
        RECT 1483.660 498.090 1483.800 510.000 ;
        RECT 1483.600 497.770 1483.860 498.090 ;
        RECT 1490.040 497.770 1490.300 498.090 ;
        RECT 1490.100 38.070 1490.240 497.770 ;
        RECT 1490.040 37.750 1490.300 38.070 ;
        RECT 1792.720 37.410 1792.980 37.730 ;
        RECT 1792.780 2.400 1792.920 37.410 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1503.810 58.720 1504.130 58.780 ;
        RECT 1807.870 58.720 1808.190 58.780 ;
        RECT 1503.810 58.580 1808.190 58.720 ;
        RECT 1503.810 58.520 1504.130 58.580 ;
        RECT 1807.870 58.520 1808.190 58.580 ;
      LAYER via ;
        RECT 1503.840 58.520 1504.100 58.780 ;
        RECT 1807.900 58.520 1808.160 58.780 ;
      LAYER met2 ;
        RECT 1500.290 510.410 1500.570 514.000 ;
        RECT 1500.290 510.270 1504.040 510.410 ;
        RECT 1500.290 510.000 1500.570 510.270 ;
        RECT 1503.900 58.810 1504.040 510.270 ;
        RECT 1503.840 58.490 1504.100 58.810 ;
        RECT 1807.900 58.490 1808.160 58.810 ;
        RECT 1807.960 17.410 1808.100 58.490 ;
        RECT 1807.960 17.270 1810.860 17.410 ;
        RECT 1810.720 2.400 1810.860 17.270 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 44.780 1517.930 44.840 ;
        RECT 1829.030 44.780 1829.350 44.840 ;
        RECT 1517.610 44.640 1829.350 44.780 ;
        RECT 1517.610 44.580 1517.930 44.640 ;
        RECT 1829.030 44.580 1829.350 44.640 ;
      LAYER via ;
        RECT 1517.640 44.580 1517.900 44.840 ;
        RECT 1829.060 44.580 1829.320 44.840 ;
      LAYER met2 ;
        RECT 1516.390 510.410 1516.670 514.000 ;
        RECT 1516.390 510.270 1517.840 510.410 ;
        RECT 1516.390 510.000 1516.670 510.270 ;
        RECT 1517.700 44.870 1517.840 510.270 ;
        RECT 1517.640 44.550 1517.900 44.870 ;
        RECT 1829.060 44.550 1829.320 44.870 ;
        RECT 1829.120 17.410 1829.260 44.550 ;
        RECT 1828.660 17.270 1829.260 17.410 ;
        RECT 1828.660 2.400 1828.800 17.270 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1532.790 496.980 1533.110 497.040 ;
        RECT 1548.890 496.980 1549.210 497.040 ;
        RECT 1532.790 496.840 1549.210 496.980 ;
        RECT 1532.790 496.780 1533.110 496.840 ;
        RECT 1548.890 496.780 1549.210 496.840 ;
        RECT 1548.890 51.920 1549.210 51.980 ;
        RECT 1842.370 51.920 1842.690 51.980 ;
        RECT 1548.890 51.780 1842.690 51.920 ;
        RECT 1548.890 51.720 1549.210 51.780 ;
        RECT 1842.370 51.720 1842.690 51.780 ;
      LAYER via ;
        RECT 1532.820 496.780 1533.080 497.040 ;
        RECT 1548.920 496.780 1549.180 497.040 ;
        RECT 1548.920 51.720 1549.180 51.980 ;
        RECT 1842.400 51.720 1842.660 51.980 ;
      LAYER met2 ;
        RECT 1532.950 510.340 1533.230 514.000 ;
        RECT 1532.880 510.000 1533.230 510.340 ;
        RECT 1532.880 497.070 1533.020 510.000 ;
        RECT 1532.820 496.750 1533.080 497.070 ;
        RECT 1548.920 496.750 1549.180 497.070 ;
        RECT 1548.980 52.010 1549.120 496.750 ;
        RECT 1548.920 51.690 1549.180 52.010 ;
        RECT 1842.400 51.690 1842.660 52.010 ;
        RECT 1842.460 16.730 1842.600 51.690 ;
        RECT 1842.460 16.590 1846.280 16.730 ;
        RECT 1846.140 2.400 1846.280 16.590 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 148.140 1552.430 148.200 ;
        RECT 1863.070 148.140 1863.390 148.200 ;
        RECT 1552.110 148.000 1863.390 148.140 ;
        RECT 1552.110 147.940 1552.430 148.000 ;
        RECT 1863.070 147.940 1863.390 148.000 ;
        RECT 1863.070 62.260 1863.390 62.520 ;
        RECT 1863.160 61.780 1863.300 62.260 ;
        RECT 1863.990 61.780 1864.310 61.840 ;
        RECT 1863.160 61.640 1864.310 61.780 ;
        RECT 1863.990 61.580 1864.310 61.640 ;
      LAYER via ;
        RECT 1552.140 147.940 1552.400 148.200 ;
        RECT 1863.100 147.940 1863.360 148.200 ;
        RECT 1863.100 62.260 1863.360 62.520 ;
        RECT 1864.020 61.580 1864.280 61.840 ;
      LAYER met2 ;
        RECT 1549.050 510.410 1549.330 514.000 ;
        RECT 1549.050 510.270 1552.340 510.410 ;
        RECT 1549.050 510.000 1549.330 510.270 ;
        RECT 1552.200 148.230 1552.340 510.270 ;
        RECT 1552.140 147.910 1552.400 148.230 ;
        RECT 1863.100 147.910 1863.360 148.230 ;
        RECT 1863.160 62.550 1863.300 147.910 ;
        RECT 1863.100 62.230 1863.360 62.550 ;
        RECT 1864.020 61.550 1864.280 61.870 ;
        RECT 1864.080 2.400 1864.220 61.550 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.010 86.260 524.330 86.320 ;
        RECT 738.370 86.260 738.690 86.320 ;
        RECT 524.010 86.120 738.690 86.260 ;
        RECT 524.010 86.060 524.330 86.120 ;
        RECT 738.370 86.060 738.690 86.120 ;
      LAYER via ;
        RECT 524.040 86.060 524.300 86.320 ;
        RECT 738.400 86.060 738.660 86.320 ;
      LAYER met2 ;
        RECT 520.950 510.410 521.230 514.000 ;
        RECT 520.950 510.270 524.240 510.410 ;
        RECT 520.950 510.000 521.230 510.270 ;
        RECT 524.100 86.350 524.240 510.270 ;
        RECT 524.040 86.030 524.300 86.350 ;
        RECT 738.400 86.030 738.660 86.350 ;
        RECT 738.460 17.410 738.600 86.030 ;
        RECT 738.460 17.270 740.440 17.410 ;
        RECT 740.300 2.400 740.440 17.270 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 155.280 1566.230 155.340 ;
        RECT 1876.870 155.280 1877.190 155.340 ;
        RECT 1565.910 155.140 1877.190 155.280 ;
        RECT 1565.910 155.080 1566.230 155.140 ;
        RECT 1876.870 155.080 1877.190 155.140 ;
        RECT 1876.870 62.120 1877.190 62.180 ;
        RECT 1881.930 62.120 1882.250 62.180 ;
        RECT 1876.870 61.980 1882.250 62.120 ;
        RECT 1876.870 61.920 1877.190 61.980 ;
        RECT 1881.930 61.920 1882.250 61.980 ;
      LAYER via ;
        RECT 1565.940 155.080 1566.200 155.340 ;
        RECT 1876.900 155.080 1877.160 155.340 ;
        RECT 1876.900 61.920 1877.160 62.180 ;
        RECT 1881.960 61.920 1882.220 62.180 ;
      LAYER met2 ;
        RECT 1565.610 510.340 1565.890 514.000 ;
        RECT 1565.540 510.000 1565.890 510.340 ;
        RECT 1565.540 497.490 1565.680 510.000 ;
        RECT 1565.540 497.350 1566.140 497.490 ;
        RECT 1566.000 155.370 1566.140 497.350 ;
        RECT 1565.940 155.050 1566.200 155.370 ;
        RECT 1876.900 155.050 1877.160 155.370 ;
        RECT 1876.960 62.210 1877.100 155.050 ;
        RECT 1876.900 61.890 1877.160 62.210 ;
        RECT 1881.960 61.890 1882.220 62.210 ;
        RECT 1882.020 2.400 1882.160 61.890 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.550 496.980 1581.870 497.040 ;
        RECT 1586.610 496.980 1586.930 497.040 ;
        RECT 1581.550 496.840 1586.930 496.980 ;
        RECT 1581.550 496.780 1581.870 496.840 ;
        RECT 1586.610 496.780 1586.930 496.840 ;
        RECT 1586.610 65.520 1586.930 65.580 ;
        RECT 1897.570 65.520 1897.890 65.580 ;
        RECT 1586.610 65.380 1897.890 65.520 ;
        RECT 1586.610 65.320 1586.930 65.380 ;
        RECT 1897.570 65.320 1897.890 65.380 ;
      LAYER via ;
        RECT 1581.580 496.780 1581.840 497.040 ;
        RECT 1586.640 496.780 1586.900 497.040 ;
        RECT 1586.640 65.320 1586.900 65.580 ;
        RECT 1897.600 65.320 1897.860 65.580 ;
      LAYER met2 ;
        RECT 1581.710 510.340 1581.990 514.000 ;
        RECT 1581.640 510.000 1581.990 510.340 ;
        RECT 1581.640 497.070 1581.780 510.000 ;
        RECT 1581.580 496.750 1581.840 497.070 ;
        RECT 1586.640 496.750 1586.900 497.070 ;
        RECT 1586.700 65.610 1586.840 496.750 ;
        RECT 1586.640 65.290 1586.900 65.610 ;
        RECT 1897.600 65.290 1897.860 65.610 ;
        RECT 1897.660 16.730 1897.800 65.290 ;
        RECT 1897.660 16.590 1900.100 16.730 ;
        RECT 1899.960 2.400 1900.100 16.590 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 72.660 1600.730 72.720 ;
        RECT 1911.830 72.660 1912.150 72.720 ;
        RECT 1600.410 72.520 1912.150 72.660 ;
        RECT 1600.410 72.460 1600.730 72.520 ;
        RECT 1911.830 72.460 1912.150 72.520 ;
        RECT 1911.830 17.920 1912.150 17.980 ;
        RECT 1917.810 17.920 1918.130 17.980 ;
        RECT 1911.830 17.780 1918.130 17.920 ;
        RECT 1911.830 17.720 1912.150 17.780 ;
        RECT 1917.810 17.720 1918.130 17.780 ;
      LAYER via ;
        RECT 1600.440 72.460 1600.700 72.720 ;
        RECT 1911.860 72.460 1912.120 72.720 ;
        RECT 1911.860 17.720 1912.120 17.980 ;
        RECT 1917.840 17.720 1918.100 17.980 ;
      LAYER met2 ;
        RECT 1598.270 510.410 1598.550 514.000 ;
        RECT 1598.270 510.270 1600.640 510.410 ;
        RECT 1598.270 510.000 1598.550 510.270 ;
        RECT 1600.500 72.750 1600.640 510.270 ;
        RECT 1600.440 72.430 1600.700 72.750 ;
        RECT 1911.860 72.430 1912.120 72.750 ;
        RECT 1911.920 18.010 1912.060 72.430 ;
        RECT 1911.860 17.690 1912.120 18.010 ;
        RECT 1917.840 17.690 1918.100 18.010 ;
        RECT 1917.900 2.400 1918.040 17.690 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 107.340 1614.530 107.400 ;
        RECT 1932.070 107.340 1932.390 107.400 ;
        RECT 1614.210 107.200 1932.390 107.340 ;
        RECT 1614.210 107.140 1614.530 107.200 ;
        RECT 1932.070 107.140 1932.390 107.200 ;
      LAYER via ;
        RECT 1614.240 107.140 1614.500 107.400 ;
        RECT 1932.100 107.140 1932.360 107.400 ;
      LAYER met2 ;
        RECT 1614.370 510.340 1614.650 514.000 ;
        RECT 1614.300 510.000 1614.650 510.340 ;
        RECT 1614.300 107.430 1614.440 510.000 ;
        RECT 1614.240 107.110 1614.500 107.430 ;
        RECT 1932.100 107.110 1932.360 107.430 ;
        RECT 1932.160 16.730 1932.300 107.110 ;
        RECT 1932.160 16.590 1935.520 16.730 ;
        RECT 1935.380 2.400 1935.520 16.590 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1630.770 502.760 1631.090 502.820 ;
        RECT 1634.910 502.760 1635.230 502.820 ;
        RECT 1630.770 502.620 1635.230 502.760 ;
        RECT 1630.770 502.560 1631.090 502.620 ;
        RECT 1634.910 502.560 1635.230 502.620 ;
        RECT 1634.910 79.460 1635.230 79.520 ;
        RECT 1953.230 79.460 1953.550 79.520 ;
        RECT 1634.910 79.320 1953.550 79.460 ;
        RECT 1634.910 79.260 1635.230 79.320 ;
        RECT 1953.230 79.260 1953.550 79.320 ;
      LAYER via ;
        RECT 1630.800 502.560 1631.060 502.820 ;
        RECT 1634.940 502.560 1635.200 502.820 ;
        RECT 1634.940 79.260 1635.200 79.520 ;
        RECT 1953.260 79.260 1953.520 79.520 ;
      LAYER met2 ;
        RECT 1630.930 510.340 1631.210 514.000 ;
        RECT 1630.860 510.000 1631.210 510.340 ;
        RECT 1630.860 502.850 1631.000 510.000 ;
        RECT 1630.800 502.530 1631.060 502.850 ;
        RECT 1634.940 502.530 1635.200 502.850 ;
        RECT 1635.000 79.550 1635.140 502.530 ;
        RECT 1634.940 79.230 1635.200 79.550 ;
        RECT 1953.260 79.230 1953.520 79.550 ;
        RECT 1953.320 2.400 1953.460 79.230 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1646.870 500.040 1647.190 500.100 ;
        RECT 1967.030 500.040 1967.350 500.100 ;
        RECT 1646.870 499.900 1967.350 500.040 ;
        RECT 1646.870 499.840 1647.190 499.900 ;
        RECT 1967.030 499.840 1967.350 499.900 ;
        RECT 1967.030 62.120 1967.350 62.180 ;
        RECT 1971.170 62.120 1971.490 62.180 ;
        RECT 1967.030 61.980 1971.490 62.120 ;
        RECT 1967.030 61.920 1967.350 61.980 ;
        RECT 1971.170 61.920 1971.490 61.980 ;
      LAYER via ;
        RECT 1646.900 499.840 1647.160 500.100 ;
        RECT 1967.060 499.840 1967.320 500.100 ;
        RECT 1967.060 61.920 1967.320 62.180 ;
        RECT 1971.200 61.920 1971.460 62.180 ;
      LAYER met2 ;
        RECT 1647.030 510.340 1647.310 514.000 ;
        RECT 1646.960 510.000 1647.310 510.340 ;
        RECT 1646.960 500.130 1647.100 510.000 ;
        RECT 1646.900 499.810 1647.160 500.130 ;
        RECT 1967.060 499.810 1967.320 500.130 ;
        RECT 1967.120 62.210 1967.260 499.810 ;
        RECT 1967.060 61.890 1967.320 62.210 ;
        RECT 1971.200 61.890 1971.460 62.210 ;
        RECT 1971.260 2.400 1971.400 61.890 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1987.345 48.365 1987.515 96.475 ;
      LAYER mcon ;
        RECT 1987.345 96.305 1987.515 96.475 ;
      LAYER met1 ;
        RECT 1663.430 498.680 1663.750 498.740 ;
        RECT 1669.410 498.680 1669.730 498.740 ;
        RECT 1663.430 498.540 1669.730 498.680 ;
        RECT 1663.430 498.480 1663.750 498.540 ;
        RECT 1669.410 498.480 1669.730 498.540 ;
        RECT 1669.410 113.800 1669.730 113.860 ;
        RECT 1987.730 113.800 1988.050 113.860 ;
        RECT 1669.410 113.660 1988.050 113.800 ;
        RECT 1669.410 113.600 1669.730 113.660 ;
        RECT 1987.730 113.600 1988.050 113.660 ;
        RECT 1987.270 96.460 1987.590 96.520 ;
        RECT 1987.075 96.320 1987.590 96.460 ;
        RECT 1987.270 96.260 1987.590 96.320 ;
        RECT 1987.285 48.520 1987.575 48.565 ;
        RECT 1989.110 48.520 1989.430 48.580 ;
        RECT 1987.285 48.380 1989.430 48.520 ;
        RECT 1987.285 48.335 1987.575 48.380 ;
        RECT 1989.110 48.320 1989.430 48.380 ;
      LAYER via ;
        RECT 1663.460 498.480 1663.720 498.740 ;
        RECT 1669.440 498.480 1669.700 498.740 ;
        RECT 1669.440 113.600 1669.700 113.860 ;
        RECT 1987.760 113.600 1988.020 113.860 ;
        RECT 1987.300 96.260 1987.560 96.520 ;
        RECT 1989.140 48.320 1989.400 48.580 ;
      LAYER met2 ;
        RECT 1663.590 510.340 1663.870 514.000 ;
        RECT 1663.520 510.000 1663.870 510.340 ;
        RECT 1663.520 498.770 1663.660 510.000 ;
        RECT 1663.460 498.450 1663.720 498.770 ;
        RECT 1669.440 498.450 1669.700 498.770 ;
        RECT 1669.500 113.890 1669.640 498.450 ;
        RECT 1669.440 113.570 1669.700 113.890 ;
        RECT 1987.760 113.570 1988.020 113.890 ;
        RECT 1987.820 96.970 1987.960 113.570 ;
        RECT 1987.360 96.830 1987.960 96.970 ;
        RECT 1987.360 96.550 1987.500 96.830 ;
        RECT 1987.300 96.230 1987.560 96.550 ;
        RECT 1989.140 48.290 1989.400 48.610 ;
        RECT 1989.200 2.400 1989.340 48.290 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 30.840 1683.530 30.900 ;
        RECT 2006.590 30.840 2006.910 30.900 ;
        RECT 1683.210 30.700 2006.910 30.840 ;
        RECT 1683.210 30.640 1683.530 30.700 ;
        RECT 2006.590 30.640 2006.910 30.700 ;
      LAYER via ;
        RECT 1683.240 30.640 1683.500 30.900 ;
        RECT 2006.620 30.640 2006.880 30.900 ;
      LAYER met2 ;
        RECT 1679.690 510.410 1679.970 514.000 ;
        RECT 1679.690 510.270 1683.440 510.410 ;
        RECT 1679.690 510.000 1679.970 510.270 ;
        RECT 1683.300 30.930 1683.440 510.270 ;
        RECT 1683.240 30.610 1683.500 30.930 ;
        RECT 2006.620 30.610 2006.880 30.930 ;
        RECT 2006.680 2.400 2006.820 30.610 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.010 86.260 1697.330 86.320 ;
        RECT 2021.770 86.260 2022.090 86.320 ;
        RECT 1697.010 86.120 2022.090 86.260 ;
        RECT 1697.010 86.060 1697.330 86.120 ;
        RECT 2021.770 86.060 2022.090 86.120 ;
      LAYER via ;
        RECT 1697.040 86.060 1697.300 86.320 ;
        RECT 2021.800 86.060 2022.060 86.320 ;
      LAYER met2 ;
        RECT 1696.250 510.410 1696.530 514.000 ;
        RECT 1696.250 510.270 1697.240 510.410 ;
        RECT 1696.250 510.000 1696.530 510.270 ;
        RECT 1697.100 86.350 1697.240 510.270 ;
        RECT 1697.040 86.030 1697.300 86.350 ;
        RECT 2021.800 86.030 2022.060 86.350 ;
        RECT 2021.860 17.410 2022.000 86.030 ;
        RECT 2021.860 17.270 2024.760 17.410 ;
        RECT 2024.620 2.400 2024.760 17.270 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1712.190 493.240 1712.510 493.300 ;
        RECT 2042.470 493.240 2042.790 493.300 ;
        RECT 1712.190 493.100 2042.790 493.240 ;
        RECT 1712.190 493.040 1712.510 493.100 ;
        RECT 2042.470 493.040 2042.790 493.100 ;
      LAYER via ;
        RECT 1712.220 493.040 1712.480 493.300 ;
        RECT 2042.500 493.040 2042.760 493.300 ;
      LAYER met2 ;
        RECT 1712.350 510.340 1712.630 514.000 ;
        RECT 1712.280 510.000 1712.630 510.340 ;
        RECT 1712.280 493.330 1712.420 510.000 ;
        RECT 1712.220 493.010 1712.480 493.330 ;
        RECT 2042.500 493.010 2042.760 493.330 ;
        RECT 2042.560 2.400 2042.700 493.010 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 497.320 537.670 497.380 ;
        RECT 569.090 497.320 569.410 497.380 ;
        RECT 537.350 497.180 569.410 497.320 ;
        RECT 537.350 497.120 537.670 497.180 ;
        RECT 569.090 497.120 569.410 497.180 ;
        RECT 569.090 93.060 569.410 93.120 ;
        RECT 752.630 93.060 752.950 93.120 ;
        RECT 569.090 92.920 752.950 93.060 ;
        RECT 569.090 92.860 569.410 92.920 ;
        RECT 752.630 92.860 752.950 92.920 ;
      LAYER via ;
        RECT 537.380 497.120 537.640 497.380 ;
        RECT 569.120 497.120 569.380 497.380 ;
        RECT 569.120 92.860 569.380 93.120 ;
        RECT 752.660 92.860 752.920 93.120 ;
      LAYER met2 ;
        RECT 537.510 510.340 537.790 514.000 ;
        RECT 537.440 510.000 537.790 510.340 ;
        RECT 537.440 497.410 537.580 510.000 ;
        RECT 537.380 497.090 537.640 497.410 ;
        RECT 569.120 497.090 569.380 497.410 ;
        RECT 569.180 93.150 569.320 497.090 ;
        RECT 569.120 92.830 569.380 93.150 ;
        RECT 752.660 92.830 752.920 93.150 ;
        RECT 752.720 17.410 752.860 92.830 ;
        RECT 752.720 17.270 757.920 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.510 93.060 1731.830 93.120 ;
        RECT 1731.510 92.920 2039.020 93.060 ;
        RECT 1731.510 92.860 1731.830 92.920 ;
        RECT 2038.880 92.720 2039.020 92.920 ;
        RECT 2060.410 92.720 2060.730 92.780 ;
        RECT 2038.880 92.580 2060.730 92.720 ;
        RECT 2060.410 92.520 2060.730 92.580 ;
      LAYER via ;
        RECT 1731.540 92.860 1731.800 93.120 ;
        RECT 2060.440 92.520 2060.700 92.780 ;
      LAYER met2 ;
        RECT 1728.450 510.410 1728.730 514.000 ;
        RECT 1728.450 510.270 1731.740 510.410 ;
        RECT 1728.450 510.000 1728.730 510.270 ;
        RECT 1731.600 93.150 1731.740 510.270 ;
        RECT 1731.540 92.830 1731.800 93.150 ;
        RECT 2060.440 92.490 2060.700 92.810 ;
        RECT 2060.500 2.400 2060.640 92.490 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2077.045 48.365 2077.215 96.475 ;
      LAYER mcon ;
        RECT 2077.045 96.305 2077.215 96.475 ;
      LAYER met1 ;
        RECT 1745.310 120.600 1745.630 120.660 ;
        RECT 2076.970 120.600 2077.290 120.660 ;
        RECT 1745.310 120.460 2077.290 120.600 ;
        RECT 1745.310 120.400 1745.630 120.460 ;
        RECT 2076.970 120.400 2077.290 120.460 ;
        RECT 2076.970 96.460 2077.290 96.520 ;
        RECT 2076.970 96.320 2077.485 96.460 ;
        RECT 2076.970 96.260 2077.290 96.320 ;
        RECT 2076.985 48.520 2077.275 48.565 ;
        RECT 2078.350 48.520 2078.670 48.580 ;
        RECT 2076.985 48.380 2078.670 48.520 ;
        RECT 2076.985 48.335 2077.275 48.380 ;
        RECT 2078.350 48.320 2078.670 48.380 ;
      LAYER via ;
        RECT 1745.340 120.400 1745.600 120.660 ;
        RECT 2077.000 120.400 2077.260 120.660 ;
        RECT 2077.000 96.260 2077.260 96.520 ;
        RECT 2078.380 48.320 2078.640 48.580 ;
      LAYER met2 ;
        RECT 1745.010 510.340 1745.290 514.000 ;
        RECT 1744.940 510.000 1745.290 510.340 ;
        RECT 1744.940 497.490 1745.080 510.000 ;
        RECT 1744.940 497.350 1745.540 497.490 ;
        RECT 1745.400 120.690 1745.540 497.350 ;
        RECT 1745.340 120.370 1745.600 120.690 ;
        RECT 2077.000 120.370 2077.260 120.690 ;
        RECT 2077.060 96.550 2077.200 120.370 ;
        RECT 2077.000 96.230 2077.260 96.550 ;
        RECT 2078.380 48.290 2078.640 48.610 ;
        RECT 2078.440 2.400 2078.580 48.290 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1780.345 24.225 1780.515 25.075 ;
        RECT 1828.185 23.885 1828.355 25.075 ;
        RECT 1828.645 24.225 1828.815 25.075 ;
        RECT 1852.565 24.225 1852.735 25.075 ;
        RECT 1883.845 23.885 1884.475 24.055 ;
      LAYER mcon ;
        RECT 1780.345 24.905 1780.515 25.075 ;
        RECT 1828.185 24.905 1828.355 25.075 ;
        RECT 1828.645 24.905 1828.815 25.075 ;
        RECT 1852.565 24.905 1852.735 25.075 ;
        RECT 1884.305 23.885 1884.475 24.055 ;
      LAYER met1 ;
        RECT 1760.950 496.980 1761.270 497.040 ;
        RECT 1766.010 496.980 1766.330 497.040 ;
        RECT 1760.950 496.840 1766.330 496.980 ;
        RECT 1760.950 496.780 1761.270 496.840 ;
        RECT 1766.010 496.780 1766.330 496.840 ;
        RECT 1780.285 25.060 1780.575 25.105 ;
        RECT 1828.125 25.060 1828.415 25.105 ;
        RECT 1780.285 24.920 1828.415 25.060 ;
        RECT 1780.285 24.875 1780.575 24.920 ;
        RECT 1828.125 24.875 1828.415 24.920 ;
        RECT 1828.585 25.060 1828.875 25.105 ;
        RECT 1852.505 25.060 1852.795 25.105 ;
        RECT 1828.585 24.920 1852.795 25.060 ;
        RECT 1828.585 24.875 1828.875 24.920 ;
        RECT 1852.505 24.875 1852.795 24.920 ;
        RECT 1766.010 24.380 1766.330 24.440 ;
        RECT 1780.285 24.380 1780.575 24.425 ;
        RECT 1766.010 24.240 1780.575 24.380 ;
        RECT 1766.010 24.180 1766.330 24.240 ;
        RECT 1780.285 24.195 1780.575 24.240 ;
        RECT 1828.585 24.195 1828.875 24.425 ;
        RECT 1852.505 24.380 1852.795 24.425 ;
        RECT 2095.830 24.380 2096.150 24.440 ;
        RECT 1852.505 24.240 1884.000 24.380 ;
        RECT 1852.505 24.195 1852.795 24.240 ;
        RECT 1828.125 24.040 1828.415 24.085 ;
        RECT 1828.660 24.040 1828.800 24.195 ;
        RECT 1883.860 24.085 1884.000 24.240 ;
        RECT 1956.080 24.240 2096.150 24.380 ;
        RECT 1828.125 23.900 1828.800 24.040 ;
        RECT 1828.125 23.855 1828.415 23.900 ;
        RECT 1883.785 23.855 1884.075 24.085 ;
        RECT 1884.245 24.040 1884.535 24.085 ;
        RECT 1956.080 24.040 1956.220 24.240 ;
        RECT 2095.830 24.180 2096.150 24.240 ;
        RECT 1884.245 23.900 1956.220 24.040 ;
        RECT 1884.245 23.855 1884.535 23.900 ;
      LAYER via ;
        RECT 1760.980 496.780 1761.240 497.040 ;
        RECT 1766.040 496.780 1766.300 497.040 ;
        RECT 1766.040 24.180 1766.300 24.440 ;
        RECT 2095.860 24.180 2096.120 24.440 ;
      LAYER met2 ;
        RECT 1761.110 510.340 1761.390 514.000 ;
        RECT 1761.040 510.000 1761.390 510.340 ;
        RECT 1761.040 497.070 1761.180 510.000 ;
        RECT 1760.980 496.750 1761.240 497.070 ;
        RECT 1766.040 496.750 1766.300 497.070 ;
        RECT 1766.100 24.470 1766.240 496.750 ;
        RECT 1766.040 24.150 1766.300 24.470 ;
        RECT 2095.860 24.150 2096.120 24.470 ;
        RECT 2095.920 2.400 2096.060 24.150 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 99.860 1780.130 99.920 ;
        RECT 2111.470 99.860 2111.790 99.920 ;
        RECT 1779.810 99.720 2111.790 99.860 ;
        RECT 1779.810 99.660 1780.130 99.720 ;
        RECT 2111.470 99.660 2111.790 99.720 ;
      LAYER via ;
        RECT 1779.840 99.660 1780.100 99.920 ;
        RECT 2111.500 99.660 2111.760 99.920 ;
      LAYER met2 ;
        RECT 1777.670 510.410 1777.950 514.000 ;
        RECT 1777.670 510.270 1780.040 510.410 ;
        RECT 1777.670 510.000 1777.950 510.270 ;
        RECT 1779.900 99.950 1780.040 510.270 ;
        RECT 1779.840 99.630 1780.100 99.950 ;
        RECT 2111.500 99.630 2111.760 99.950 ;
        RECT 2111.560 17.410 2111.700 99.630 ;
        RECT 2111.560 17.270 2114.000 17.410 ;
        RECT 2113.860 2.400 2114.000 17.270 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 38.320 1793.930 38.380 ;
        RECT 2131.710 38.320 2132.030 38.380 ;
        RECT 1793.610 38.180 2132.030 38.320 ;
        RECT 1793.610 38.120 1793.930 38.180 ;
        RECT 2131.710 38.120 2132.030 38.180 ;
      LAYER via ;
        RECT 1793.640 38.120 1793.900 38.380 ;
        RECT 2131.740 38.120 2132.000 38.380 ;
      LAYER met2 ;
        RECT 1793.770 510.340 1794.050 514.000 ;
        RECT 1793.700 510.000 1794.050 510.340 ;
        RECT 1793.700 38.410 1793.840 510.000 ;
        RECT 1793.640 38.090 1793.900 38.410 ;
        RECT 2131.740 38.090 2132.000 38.410 ;
        RECT 2131.800 2.400 2131.940 38.090 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1810.170 496.980 1810.490 497.040 ;
        RECT 1814.310 496.980 1814.630 497.040 ;
        RECT 1810.170 496.840 1814.630 496.980 ;
        RECT 1810.170 496.780 1810.490 496.840 ;
        RECT 1814.310 496.780 1814.630 496.840 ;
        RECT 1814.310 127.740 1814.630 127.800 ;
        RECT 2145.970 127.740 2146.290 127.800 ;
        RECT 1814.310 127.600 2146.290 127.740 ;
        RECT 1814.310 127.540 1814.630 127.600 ;
        RECT 2145.970 127.540 2146.290 127.600 ;
      LAYER via ;
        RECT 1810.200 496.780 1810.460 497.040 ;
        RECT 1814.340 496.780 1814.600 497.040 ;
        RECT 1814.340 127.540 1814.600 127.800 ;
        RECT 2146.000 127.540 2146.260 127.800 ;
      LAYER met2 ;
        RECT 1810.330 510.340 1810.610 514.000 ;
        RECT 1810.260 510.000 1810.610 510.340 ;
        RECT 1810.260 497.070 1810.400 510.000 ;
        RECT 1810.200 496.750 1810.460 497.070 ;
        RECT 1814.340 496.750 1814.600 497.070 ;
        RECT 1814.400 127.830 1814.540 496.750 ;
        RECT 1814.340 127.510 1814.600 127.830 ;
        RECT 2146.000 127.510 2146.260 127.830 ;
        RECT 2146.060 17.410 2146.200 127.510 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 196.760 1828.430 196.820 ;
        RECT 2167.130 196.760 2167.450 196.820 ;
        RECT 1828.110 196.620 2167.450 196.760 ;
        RECT 1828.110 196.560 1828.430 196.620 ;
        RECT 2167.130 196.560 2167.450 196.620 ;
      LAYER via ;
        RECT 1828.140 196.560 1828.400 196.820 ;
        RECT 2167.160 196.560 2167.420 196.820 ;
      LAYER met2 ;
        RECT 1826.430 510.410 1826.710 514.000 ;
        RECT 1826.430 510.270 1828.340 510.410 ;
        RECT 1826.430 510.000 1826.710 510.270 ;
        RECT 1828.200 196.850 1828.340 510.270 ;
        RECT 1828.140 196.530 1828.400 196.850 ;
        RECT 2167.160 196.530 2167.420 196.850 ;
        RECT 2167.220 17.410 2167.360 196.530 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1842.830 496.980 1843.150 497.040 ;
        RECT 1848.810 496.980 1849.130 497.040 ;
        RECT 1842.830 496.840 1849.130 496.980 ;
        RECT 1842.830 496.780 1843.150 496.840 ;
        RECT 1848.810 496.780 1849.130 496.840 ;
        RECT 1848.810 44.780 1849.130 44.840 ;
        RECT 2185.070 44.780 2185.390 44.840 ;
        RECT 1848.810 44.640 2185.390 44.780 ;
        RECT 1848.810 44.580 1849.130 44.640 ;
        RECT 2185.070 44.580 2185.390 44.640 ;
      LAYER via ;
        RECT 1842.860 496.780 1843.120 497.040 ;
        RECT 1848.840 496.780 1849.100 497.040 ;
        RECT 1848.840 44.580 1849.100 44.840 ;
        RECT 2185.100 44.580 2185.360 44.840 ;
      LAYER met2 ;
        RECT 1842.990 510.340 1843.270 514.000 ;
        RECT 1842.920 510.000 1843.270 510.340 ;
        RECT 1842.920 497.070 1843.060 510.000 ;
        RECT 1842.860 496.750 1843.120 497.070 ;
        RECT 1848.840 496.750 1849.100 497.070 ;
        RECT 1848.900 44.870 1849.040 496.750 ;
        RECT 1848.840 44.550 1849.100 44.870 ;
        RECT 2185.100 44.550 2185.360 44.870 ;
        RECT 2185.160 2.400 2185.300 44.550 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 134.540 1862.930 134.600 ;
        RECT 2201.170 134.540 2201.490 134.600 ;
        RECT 1862.610 134.400 2201.490 134.540 ;
        RECT 1862.610 134.340 1862.930 134.400 ;
        RECT 2201.170 134.340 2201.490 134.400 ;
      LAYER via ;
        RECT 1862.640 134.340 1862.900 134.600 ;
        RECT 2201.200 134.340 2201.460 134.600 ;
      LAYER met2 ;
        RECT 1859.090 510.410 1859.370 514.000 ;
        RECT 1859.090 510.270 1862.840 510.410 ;
        RECT 1859.090 510.000 1859.370 510.270 ;
        RECT 1862.700 134.630 1862.840 510.270 ;
        RECT 1862.640 134.310 1862.900 134.630 ;
        RECT 2201.200 134.310 2201.460 134.630 ;
        RECT 2201.260 17.410 2201.400 134.310 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 141.340 1876.730 141.400 ;
        RECT 2215.430 141.340 2215.750 141.400 ;
        RECT 1876.410 141.200 2215.750 141.340 ;
        RECT 1876.410 141.140 1876.730 141.200 ;
        RECT 2215.430 141.140 2215.750 141.200 ;
      LAYER via ;
        RECT 1876.440 141.140 1876.700 141.400 ;
        RECT 2215.460 141.140 2215.720 141.400 ;
      LAYER met2 ;
        RECT 1875.650 510.410 1875.930 514.000 ;
        RECT 1875.650 510.270 1876.640 510.410 ;
        RECT 1875.650 510.000 1875.930 510.270 ;
        RECT 1876.500 141.430 1876.640 510.270 ;
        RECT 1876.440 141.110 1876.700 141.430 ;
        RECT 2215.460 141.110 2215.720 141.430 ;
        RECT 2215.520 17.410 2215.660 141.110 ;
        RECT 2215.520 17.270 2221.180 17.410 ;
        RECT 2221.040 2.400 2221.180 17.270 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 553.450 496.980 553.770 497.040 ;
        RECT 558.510 496.980 558.830 497.040 ;
        RECT 553.450 496.840 558.830 496.980 ;
        RECT 553.450 496.780 553.770 496.840 ;
        RECT 558.510 496.780 558.830 496.840 ;
        RECT 558.510 99.860 558.830 99.920 ;
        RECT 772.870 99.860 773.190 99.920 ;
        RECT 558.510 99.720 773.190 99.860 ;
        RECT 558.510 99.660 558.830 99.720 ;
        RECT 772.870 99.660 773.190 99.720 ;
      LAYER via ;
        RECT 553.480 496.780 553.740 497.040 ;
        RECT 558.540 496.780 558.800 497.040 ;
        RECT 558.540 99.660 558.800 99.920 ;
        RECT 772.900 99.660 773.160 99.920 ;
      LAYER met2 ;
        RECT 553.610 510.340 553.890 514.000 ;
        RECT 553.540 510.000 553.890 510.340 ;
        RECT 553.540 497.070 553.680 510.000 ;
        RECT 553.480 496.750 553.740 497.070 ;
        RECT 558.540 496.750 558.800 497.070 ;
        RECT 558.600 99.950 558.740 496.750 ;
        RECT 558.540 99.630 558.800 99.950 ;
        RECT 772.900 99.630 773.160 99.950 ;
        RECT 772.960 16.730 773.100 99.630 ;
        RECT 772.960 16.590 775.860 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.590 496.980 1891.910 497.040 ;
        RECT 1900.790 496.980 1901.110 497.040 ;
        RECT 1891.590 496.840 1901.110 496.980 ;
        RECT 1891.590 496.780 1891.910 496.840 ;
        RECT 1900.790 496.780 1901.110 496.840 ;
        RECT 1900.790 148.140 1901.110 148.200 ;
        RECT 2235.670 148.140 2235.990 148.200 ;
        RECT 1900.790 148.000 2235.990 148.140 ;
        RECT 1900.790 147.940 1901.110 148.000 ;
        RECT 2235.670 147.940 2235.990 148.000 ;
      LAYER via ;
        RECT 1891.620 496.780 1891.880 497.040 ;
        RECT 1900.820 496.780 1901.080 497.040 ;
        RECT 1900.820 147.940 1901.080 148.200 ;
        RECT 2235.700 147.940 2235.960 148.200 ;
      LAYER met2 ;
        RECT 1891.750 510.340 1892.030 514.000 ;
        RECT 1891.680 510.000 1892.030 510.340 ;
        RECT 1891.680 497.070 1891.820 510.000 ;
        RECT 1891.620 496.750 1891.880 497.070 ;
        RECT 1900.820 496.750 1901.080 497.070 ;
        RECT 1900.880 148.230 1901.020 496.750 ;
        RECT 1900.820 147.910 1901.080 148.230 ;
        RECT 2235.700 147.910 2235.960 148.230 ;
        RECT 2235.760 17.410 2235.900 147.910 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.910 72.320 1911.230 72.380 ;
        RECT 2256.830 72.320 2257.150 72.380 ;
        RECT 1910.910 72.180 2257.150 72.320 ;
        RECT 1910.910 72.120 1911.230 72.180 ;
        RECT 2256.830 72.120 2257.150 72.180 ;
      LAYER via ;
        RECT 1910.940 72.120 1911.200 72.380 ;
        RECT 2256.860 72.120 2257.120 72.380 ;
      LAYER met2 ;
        RECT 1908.310 510.410 1908.590 514.000 ;
        RECT 1908.310 510.270 1911.140 510.410 ;
        RECT 1908.310 510.000 1908.590 510.270 ;
        RECT 1911.000 72.410 1911.140 510.270 ;
        RECT 1910.940 72.090 1911.200 72.410 ;
        RECT 2256.860 72.090 2257.120 72.410 ;
        RECT 2256.920 7.210 2257.060 72.090 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.250 107.000 1924.570 107.060 ;
        RECT 2270.170 107.000 2270.490 107.060 ;
        RECT 1924.250 106.860 2270.490 107.000 ;
        RECT 1924.250 106.800 1924.570 106.860 ;
        RECT 2270.170 106.800 2270.490 106.860 ;
      LAYER via ;
        RECT 1924.280 106.800 1924.540 107.060 ;
        RECT 2270.200 106.800 2270.460 107.060 ;
      LAYER met2 ;
        RECT 1924.410 510.340 1924.690 514.000 ;
        RECT 1924.340 510.000 1924.690 510.340 ;
        RECT 1924.340 107.090 1924.480 510.000 ;
        RECT 1924.280 106.770 1924.540 107.090 ;
        RECT 2270.200 106.770 2270.460 107.090 ;
        RECT 2270.260 17.410 2270.400 106.770 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1940.810 496.980 1941.130 497.040 ;
        RECT 1945.410 496.980 1945.730 497.040 ;
        RECT 1940.810 496.840 1945.730 496.980 ;
        RECT 1940.810 496.780 1941.130 496.840 ;
        RECT 1945.410 496.780 1945.730 496.840 ;
        RECT 1945.410 155.280 1945.730 155.340 ;
        RECT 2290.870 155.280 2291.190 155.340 ;
        RECT 1945.410 155.140 2291.190 155.280 ;
        RECT 1945.410 155.080 1945.730 155.140 ;
        RECT 2290.870 155.080 2291.190 155.140 ;
      LAYER via ;
        RECT 1940.840 496.780 1941.100 497.040 ;
        RECT 1945.440 496.780 1945.700 497.040 ;
        RECT 1945.440 155.080 1945.700 155.340 ;
        RECT 2290.900 155.080 2291.160 155.340 ;
      LAYER met2 ;
        RECT 1940.970 510.340 1941.250 514.000 ;
        RECT 1940.900 510.000 1941.250 510.340 ;
        RECT 1940.900 497.070 1941.040 510.000 ;
        RECT 1940.840 496.750 1941.100 497.070 ;
        RECT 1945.440 496.750 1945.700 497.070 ;
        RECT 1945.500 155.370 1945.640 496.750 ;
        RECT 1945.440 155.050 1945.700 155.370 ;
        RECT 2290.900 155.050 2291.160 155.370 ;
        RECT 2290.960 17.410 2291.100 155.050 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1959.210 162.080 1959.530 162.140 ;
        RECT 2304.670 162.080 2304.990 162.140 ;
        RECT 1959.210 161.940 2304.990 162.080 ;
        RECT 1959.210 161.880 1959.530 161.940 ;
        RECT 2304.670 161.880 2304.990 161.940 ;
      LAYER via ;
        RECT 1959.240 161.880 1959.500 162.140 ;
        RECT 2304.700 161.880 2304.960 162.140 ;
      LAYER met2 ;
        RECT 1957.070 510.410 1957.350 514.000 ;
        RECT 1957.070 510.270 1959.440 510.410 ;
        RECT 1957.070 510.000 1957.350 510.270 ;
        RECT 1959.300 162.170 1959.440 510.270 ;
        RECT 1959.240 161.850 1959.500 162.170 ;
        RECT 2304.700 161.850 2304.960 162.170 ;
        RECT 2304.760 17.410 2304.900 161.850 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.470 498.000 1973.790 498.060 ;
        RECT 1979.910 498.000 1980.230 498.060 ;
        RECT 1973.470 497.860 1980.230 498.000 ;
        RECT 1973.470 497.800 1973.790 497.860 ;
        RECT 1979.910 497.800 1980.230 497.860 ;
        RECT 1979.910 168.880 1980.230 168.940 ;
        RECT 2325.370 168.880 2325.690 168.940 ;
        RECT 1979.910 168.740 2325.690 168.880 ;
        RECT 1979.910 168.680 1980.230 168.740 ;
        RECT 2325.370 168.680 2325.690 168.740 ;
      LAYER via ;
        RECT 1973.500 497.800 1973.760 498.060 ;
        RECT 1979.940 497.800 1980.200 498.060 ;
        RECT 1979.940 168.680 1980.200 168.940 ;
        RECT 2325.400 168.680 2325.660 168.940 ;
      LAYER met2 ;
        RECT 1973.630 510.340 1973.910 514.000 ;
        RECT 1973.560 510.000 1973.910 510.340 ;
        RECT 1973.560 498.090 1973.700 510.000 ;
        RECT 1973.500 497.770 1973.760 498.090 ;
        RECT 1979.940 497.770 1980.200 498.090 ;
        RECT 1980.000 168.970 1980.140 497.770 ;
        RECT 1979.940 168.650 1980.200 168.970 ;
        RECT 2325.400 168.650 2325.660 168.970 ;
        RECT 2325.460 17.410 2325.600 168.650 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1989.570 503.440 1989.890 503.500 ;
        RECT 1993.710 503.440 1994.030 503.500 ;
        RECT 1989.570 503.300 1994.030 503.440 ;
        RECT 1989.570 503.240 1989.890 503.300 ;
        RECT 1993.710 503.240 1994.030 503.300 ;
        RECT 1993.710 176.020 1994.030 176.080 ;
        RECT 2339.630 176.020 2339.950 176.080 ;
        RECT 1993.710 175.880 2339.950 176.020 ;
        RECT 1993.710 175.820 1994.030 175.880 ;
        RECT 2339.630 175.820 2339.950 175.880 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.610 16.900 2345.930 16.960 ;
        RECT 2339.630 16.760 2345.930 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.610 16.700 2345.930 16.760 ;
      LAYER via ;
        RECT 1989.600 503.240 1989.860 503.500 ;
        RECT 1993.740 503.240 1994.000 503.500 ;
        RECT 1993.740 175.820 1994.000 176.080 ;
        RECT 2339.660 175.820 2339.920 176.080 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.640 16.700 2345.900 16.960 ;
      LAYER met2 ;
        RECT 1989.730 510.340 1990.010 514.000 ;
        RECT 1989.660 510.000 1990.010 510.340 ;
        RECT 1989.660 503.530 1989.800 510.000 ;
        RECT 1989.600 503.210 1989.860 503.530 ;
        RECT 1993.740 503.210 1994.000 503.530 ;
        RECT 1993.800 176.110 1993.940 503.210 ;
        RECT 1993.740 175.790 1994.000 176.110 ;
        RECT 2339.660 175.790 2339.920 176.110 ;
        RECT 2339.720 16.990 2339.860 175.790 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.640 16.670 2345.900 16.990 ;
        RECT 2345.700 2.400 2345.840 16.670 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 182.820 2007.830 182.880 ;
        RECT 2359.870 182.820 2360.190 182.880 ;
        RECT 2007.510 182.680 2360.190 182.820 ;
        RECT 2007.510 182.620 2007.830 182.680 ;
        RECT 2359.870 182.620 2360.190 182.680 ;
      LAYER via ;
        RECT 2007.540 182.620 2007.800 182.880 ;
        RECT 2359.900 182.620 2360.160 182.880 ;
      LAYER met2 ;
        RECT 2006.290 510.410 2006.570 514.000 ;
        RECT 2006.290 510.270 2007.740 510.410 ;
        RECT 2006.290 510.000 2006.570 510.270 ;
        RECT 2007.600 182.910 2007.740 510.270 ;
        RECT 2007.540 182.590 2007.800 182.910 ;
        RECT 2359.900 182.590 2360.160 182.910 ;
        RECT 2359.960 16.730 2360.100 182.590 ;
        RECT 2359.960 16.590 2363.780 16.730 ;
        RECT 2363.640 2.400 2363.780 16.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2022.230 496.980 2022.550 497.040 ;
        RECT 2028.210 496.980 2028.530 497.040 ;
        RECT 2022.230 496.840 2028.530 496.980 ;
        RECT 2022.230 496.780 2022.550 496.840 ;
        RECT 2028.210 496.780 2028.530 496.840 ;
        RECT 2028.210 189.620 2028.530 189.680 ;
        RECT 2380.570 189.620 2380.890 189.680 ;
        RECT 2028.210 189.480 2380.890 189.620 ;
        RECT 2028.210 189.420 2028.530 189.480 ;
        RECT 2380.570 189.420 2380.890 189.480 ;
      LAYER via ;
        RECT 2022.260 496.780 2022.520 497.040 ;
        RECT 2028.240 496.780 2028.500 497.040 ;
        RECT 2028.240 189.420 2028.500 189.680 ;
        RECT 2380.600 189.420 2380.860 189.680 ;
      LAYER met2 ;
        RECT 2022.390 510.340 2022.670 514.000 ;
        RECT 2022.320 510.000 2022.670 510.340 ;
        RECT 2022.320 497.070 2022.460 510.000 ;
        RECT 2022.260 496.750 2022.520 497.070 ;
        RECT 2028.240 496.750 2028.500 497.070 ;
        RECT 2028.300 189.710 2028.440 496.750 ;
        RECT 2028.240 189.390 2028.500 189.710 ;
        RECT 2380.600 189.390 2380.860 189.710 ;
        RECT 2380.660 16.730 2380.800 189.390 ;
        RECT 2380.660 16.590 2381.720 16.730 ;
        RECT 2381.580 2.400 2381.720 16.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 203.560 2042.330 203.620 ;
        RECT 2394.370 203.560 2394.690 203.620 ;
        RECT 2042.010 203.420 2394.690 203.560 ;
        RECT 2042.010 203.360 2042.330 203.420 ;
        RECT 2394.370 203.360 2394.690 203.420 ;
      LAYER via ;
        RECT 2042.040 203.360 2042.300 203.620 ;
        RECT 2394.400 203.360 2394.660 203.620 ;
      LAYER met2 ;
        RECT 2038.950 510.410 2039.230 514.000 ;
        RECT 2038.950 510.270 2042.240 510.410 ;
        RECT 2038.950 510.000 2039.230 510.270 ;
        RECT 2042.100 203.650 2042.240 510.270 ;
        RECT 2042.040 203.330 2042.300 203.650 ;
        RECT 2394.400 203.330 2394.660 203.650 ;
        RECT 2394.460 16.730 2394.600 203.330 ;
        RECT 2394.460 16.590 2399.660 16.730 ;
        RECT 2399.520 2.400 2399.660 16.590 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 107.000 572.630 107.060 ;
        RECT 794.030 107.000 794.350 107.060 ;
        RECT 572.310 106.860 794.350 107.000 ;
        RECT 572.310 106.800 572.630 106.860 ;
        RECT 794.030 106.800 794.350 106.860 ;
      LAYER via ;
        RECT 572.340 106.800 572.600 107.060 ;
        RECT 794.060 106.800 794.320 107.060 ;
      LAYER met2 ;
        RECT 569.710 510.410 569.990 514.000 ;
        RECT 569.710 510.270 572.540 510.410 ;
        RECT 569.710 510.000 569.990 510.270 ;
        RECT 572.400 107.090 572.540 510.270 ;
        RECT 572.340 106.770 572.600 107.090 ;
        RECT 794.060 106.770 794.320 107.090 ;
        RECT 794.120 7.210 794.260 106.770 ;
        RECT 793.660 7.070 794.260 7.210 ;
        RECT 793.660 2.400 793.800 7.070 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 428.330 500.040 428.650 500.100 ;
        RECT 486.290 500.040 486.610 500.100 ;
        RECT 428.330 499.900 486.610 500.040 ;
        RECT 428.330 499.840 428.650 499.900 ;
        RECT 486.290 499.840 486.610 499.900 ;
        RECT 486.290 65.520 486.610 65.580 ;
        RECT 634.870 65.520 635.190 65.580 ;
        RECT 486.290 65.380 635.190 65.520 ;
        RECT 486.290 65.320 486.610 65.380 ;
        RECT 634.870 65.320 635.190 65.380 ;
        RECT 634.870 2.960 635.190 3.020 ;
        RECT 639.010 2.960 639.330 3.020 ;
        RECT 634.870 2.820 639.330 2.960 ;
        RECT 634.870 2.760 635.190 2.820 ;
        RECT 639.010 2.760 639.330 2.820 ;
      LAYER via ;
        RECT 428.360 499.840 428.620 500.100 ;
        RECT 486.320 499.840 486.580 500.100 ;
        RECT 486.320 65.320 486.580 65.580 ;
        RECT 634.900 65.320 635.160 65.580 ;
        RECT 634.900 2.760 635.160 3.020 ;
        RECT 639.040 2.760 639.300 3.020 ;
      LAYER met2 ;
        RECT 428.490 510.340 428.770 514.000 ;
        RECT 428.420 510.000 428.770 510.340 ;
        RECT 428.420 500.130 428.560 510.000 ;
        RECT 428.360 499.810 428.620 500.130 ;
        RECT 486.320 499.810 486.580 500.130 ;
        RECT 486.380 65.610 486.520 499.810 ;
        RECT 486.320 65.290 486.580 65.610 ;
        RECT 634.900 65.290 635.160 65.610 ;
        RECT 634.960 3.050 635.100 65.290 ;
        RECT 634.900 2.730 635.160 3.050 ;
        RECT 639.040 2.730 639.300 3.050 ;
        RECT 639.100 2.400 639.240 2.730 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.710 210.360 2063.030 210.420 ;
        RECT 2421.970 210.360 2422.290 210.420 ;
        RECT 2062.710 210.220 2422.290 210.360 ;
        RECT 2062.710 210.160 2063.030 210.220 ;
        RECT 2421.970 210.160 2422.290 210.220 ;
      LAYER via ;
        RECT 2062.740 210.160 2063.000 210.420 ;
        RECT 2422.000 210.160 2422.260 210.420 ;
      LAYER met2 ;
        RECT 2060.570 510.410 2060.850 514.000 ;
        RECT 2060.570 510.270 2062.940 510.410 ;
        RECT 2060.570 510.000 2060.850 510.270 ;
        RECT 2062.800 210.450 2062.940 510.270 ;
        RECT 2062.740 210.130 2063.000 210.450 ;
        RECT 2422.000 210.130 2422.260 210.450 ;
        RECT 2422.060 17.410 2422.200 210.130 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2076.510 217.160 2076.830 217.220 ;
        RECT 2435.770 217.160 2436.090 217.220 ;
        RECT 2076.510 217.020 2436.090 217.160 ;
        RECT 2076.510 216.960 2076.830 217.020 ;
        RECT 2435.770 216.960 2436.090 217.020 ;
      LAYER via ;
        RECT 2076.540 216.960 2076.800 217.220 ;
        RECT 2435.800 216.960 2436.060 217.220 ;
      LAYER met2 ;
        RECT 2076.670 510.340 2076.950 514.000 ;
        RECT 2076.600 510.000 2076.950 510.340 ;
        RECT 2076.600 217.250 2076.740 510.000 ;
        RECT 2076.540 216.930 2076.800 217.250 ;
        RECT 2435.800 216.930 2436.060 217.250 ;
        RECT 2435.860 17.410 2436.000 216.930 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2093.070 503.440 2093.390 503.500 ;
        RECT 2097.210 503.440 2097.530 503.500 ;
        RECT 2093.070 503.300 2097.530 503.440 ;
        RECT 2093.070 503.240 2093.390 503.300 ;
        RECT 2097.210 503.240 2097.530 503.300 ;
        RECT 2097.210 444.960 2097.530 445.020 ;
        RECT 2456.470 444.960 2456.790 445.020 ;
        RECT 2097.210 444.820 2456.790 444.960 ;
        RECT 2097.210 444.760 2097.530 444.820 ;
        RECT 2456.470 444.760 2456.790 444.820 ;
      LAYER via ;
        RECT 2093.100 503.240 2093.360 503.500 ;
        RECT 2097.240 503.240 2097.500 503.500 ;
        RECT 2097.240 444.760 2097.500 445.020 ;
        RECT 2456.500 444.760 2456.760 445.020 ;
      LAYER met2 ;
        RECT 2093.230 510.340 2093.510 514.000 ;
        RECT 2093.160 510.000 2093.510 510.340 ;
        RECT 2093.160 503.530 2093.300 510.000 ;
        RECT 2093.100 503.210 2093.360 503.530 ;
        RECT 2097.240 503.210 2097.500 503.530 ;
        RECT 2097.300 445.050 2097.440 503.210 ;
        RECT 2097.240 444.730 2097.500 445.050 ;
        RECT 2456.500 444.730 2456.760 445.050 ;
        RECT 2456.560 18.090 2456.700 444.730 ;
        RECT 2456.560 17.950 2459.000 18.090 ;
        RECT 2458.860 2.400 2459.000 17.950 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2111.010 224.300 2111.330 224.360 ;
        RECT 2470.270 224.300 2470.590 224.360 ;
        RECT 2111.010 224.160 2470.590 224.300 ;
        RECT 2111.010 224.100 2111.330 224.160 ;
        RECT 2470.270 224.100 2470.590 224.160 ;
        RECT 2470.270 17.580 2470.590 17.640 ;
        RECT 2476.710 17.580 2477.030 17.640 ;
        RECT 2470.270 17.440 2477.030 17.580 ;
        RECT 2470.270 17.380 2470.590 17.440 ;
        RECT 2476.710 17.380 2477.030 17.440 ;
      LAYER via ;
        RECT 2111.040 224.100 2111.300 224.360 ;
        RECT 2470.300 224.100 2470.560 224.360 ;
        RECT 2470.300 17.380 2470.560 17.640 ;
        RECT 2476.740 17.380 2477.000 17.640 ;
      LAYER met2 ;
        RECT 2109.330 510.410 2109.610 514.000 ;
        RECT 2109.330 510.270 2111.240 510.410 ;
        RECT 2109.330 510.000 2109.610 510.270 ;
        RECT 2111.100 224.390 2111.240 510.270 ;
        RECT 2111.040 224.070 2111.300 224.390 ;
        RECT 2470.300 224.070 2470.560 224.390 ;
        RECT 2470.360 17.670 2470.500 224.070 ;
        RECT 2470.300 17.350 2470.560 17.670 ;
        RECT 2476.740 17.350 2477.000 17.670 ;
        RECT 2476.800 2.400 2476.940 17.350 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2125.730 503.440 2126.050 503.500 ;
        RECT 2135.390 503.440 2135.710 503.500 ;
        RECT 2125.730 503.300 2135.710 503.440 ;
        RECT 2125.730 503.240 2126.050 503.300 ;
        RECT 2135.390 503.240 2135.710 503.300 ;
        RECT 2135.390 245.040 2135.710 245.100 ;
        RECT 2490.970 245.040 2491.290 245.100 ;
        RECT 2135.390 244.900 2491.290 245.040 ;
        RECT 2135.390 244.840 2135.710 244.900 ;
        RECT 2490.970 244.840 2491.290 244.900 ;
        RECT 2490.970 14.180 2491.290 14.240 ;
        RECT 2490.970 14.040 2494.880 14.180 ;
        RECT 2490.970 13.980 2491.290 14.040 ;
        RECT 2494.740 13.900 2494.880 14.040 ;
        RECT 2494.650 13.640 2494.970 13.900 ;
      LAYER via ;
        RECT 2125.760 503.240 2126.020 503.500 ;
        RECT 2135.420 503.240 2135.680 503.500 ;
        RECT 2135.420 244.840 2135.680 245.100 ;
        RECT 2491.000 244.840 2491.260 245.100 ;
        RECT 2491.000 13.980 2491.260 14.240 ;
        RECT 2494.680 13.640 2494.940 13.900 ;
      LAYER met2 ;
        RECT 2125.890 510.340 2126.170 514.000 ;
        RECT 2125.820 510.000 2126.170 510.340 ;
        RECT 2125.820 503.530 2125.960 510.000 ;
        RECT 2125.760 503.210 2126.020 503.530 ;
        RECT 2135.420 503.210 2135.680 503.530 ;
        RECT 2135.480 245.130 2135.620 503.210 ;
        RECT 2135.420 244.810 2135.680 245.130 ;
        RECT 2491.000 244.810 2491.260 245.130 ;
        RECT 2491.060 14.270 2491.200 244.810 ;
        RECT 2491.000 13.950 2491.260 14.270 ;
        RECT 2494.680 13.610 2494.940 13.930 ;
        RECT 2494.740 2.400 2494.880 13.610 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2141.830 496.980 2142.150 497.040 ;
        RECT 2145.510 496.980 2145.830 497.040 ;
        RECT 2141.830 496.840 2145.830 496.980 ;
        RECT 2141.830 496.780 2142.150 496.840 ;
        RECT 2145.510 496.780 2145.830 496.840 ;
        RECT 2145.510 231.100 2145.830 231.160 ;
        RECT 2512.130 231.100 2512.450 231.160 ;
        RECT 2145.510 230.960 2512.450 231.100 ;
        RECT 2145.510 230.900 2145.830 230.960 ;
        RECT 2512.130 230.900 2512.450 230.960 ;
      LAYER via ;
        RECT 2141.860 496.780 2142.120 497.040 ;
        RECT 2145.540 496.780 2145.800 497.040 ;
        RECT 2145.540 230.900 2145.800 231.160 ;
        RECT 2512.160 230.900 2512.420 231.160 ;
      LAYER met2 ;
        RECT 2141.990 510.340 2142.270 514.000 ;
        RECT 2141.920 510.000 2142.270 510.340 ;
        RECT 2141.920 497.070 2142.060 510.000 ;
        RECT 2141.860 496.750 2142.120 497.070 ;
        RECT 2145.540 496.750 2145.800 497.070 ;
        RECT 2145.600 231.190 2145.740 496.750 ;
        RECT 2145.540 230.870 2145.800 231.190 ;
        RECT 2512.160 230.870 2512.420 231.190 ;
        RECT 2512.220 2.400 2512.360 230.870 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2159.310 251.840 2159.630 251.900 ;
        RECT 2525.470 251.840 2525.790 251.900 ;
        RECT 2159.310 251.700 2525.790 251.840 ;
        RECT 2159.310 251.640 2159.630 251.700 ;
        RECT 2525.470 251.640 2525.790 251.700 ;
      LAYER via ;
        RECT 2159.340 251.640 2159.600 251.900 ;
        RECT 2525.500 251.640 2525.760 251.900 ;
      LAYER met2 ;
        RECT 2158.550 510.410 2158.830 514.000 ;
        RECT 2158.550 510.270 2159.540 510.410 ;
        RECT 2158.550 510.000 2158.830 510.270 ;
        RECT 2159.400 251.930 2159.540 510.270 ;
        RECT 2159.340 251.610 2159.600 251.930 ;
        RECT 2525.500 251.610 2525.760 251.930 ;
        RECT 2525.560 17.410 2525.700 251.610 ;
        RECT 2525.560 17.270 2530.300 17.410 ;
        RECT 2530.160 2.400 2530.300 17.270 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2174.490 496.980 2174.810 497.040 ;
        RECT 2179.550 496.980 2179.870 497.040 ;
        RECT 2174.490 496.840 2179.870 496.980 ;
        RECT 2174.490 496.780 2174.810 496.840 ;
        RECT 2179.550 496.780 2179.870 496.840 ;
        RECT 2179.550 458.900 2179.870 458.960 ;
        RECT 2546.170 458.900 2546.490 458.960 ;
        RECT 2179.550 458.760 2546.490 458.900 ;
        RECT 2179.550 458.700 2179.870 458.760 ;
        RECT 2546.170 458.700 2546.490 458.760 ;
      LAYER via ;
        RECT 2174.520 496.780 2174.780 497.040 ;
        RECT 2179.580 496.780 2179.840 497.040 ;
        RECT 2179.580 458.700 2179.840 458.960 ;
        RECT 2546.200 458.700 2546.460 458.960 ;
      LAYER met2 ;
        RECT 2174.650 510.340 2174.930 514.000 ;
        RECT 2174.580 510.000 2174.930 510.340 ;
        RECT 2174.580 497.070 2174.720 510.000 ;
        RECT 2174.520 496.750 2174.780 497.070 ;
        RECT 2179.580 496.750 2179.840 497.070 ;
        RECT 2179.640 458.990 2179.780 496.750 ;
        RECT 2179.580 458.670 2179.840 458.990 ;
        RECT 2546.200 458.670 2546.460 458.990 ;
        RECT 2546.260 17.410 2546.400 458.670 ;
        RECT 2546.260 17.270 2548.240 17.410 ;
        RECT 2548.100 2.400 2548.240 17.270 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2193.810 196.760 2194.130 196.820 ;
        RECT 2559.970 196.760 2560.290 196.820 ;
        RECT 2193.810 196.620 2560.290 196.760 ;
        RECT 2193.810 196.560 2194.130 196.620 ;
        RECT 2559.970 196.560 2560.290 196.620 ;
        RECT 2559.970 16.900 2560.290 16.960 ;
        RECT 2565.950 16.900 2566.270 16.960 ;
        RECT 2559.970 16.760 2566.270 16.900 ;
        RECT 2559.970 16.700 2560.290 16.760 ;
        RECT 2565.950 16.700 2566.270 16.760 ;
      LAYER via ;
        RECT 2193.840 196.560 2194.100 196.820 ;
        RECT 2560.000 196.560 2560.260 196.820 ;
        RECT 2560.000 16.700 2560.260 16.960 ;
        RECT 2565.980 16.700 2566.240 16.960 ;
      LAYER met2 ;
        RECT 2191.210 510.410 2191.490 514.000 ;
        RECT 2191.210 510.270 2194.040 510.410 ;
        RECT 2191.210 510.000 2191.490 510.270 ;
        RECT 2193.900 196.850 2194.040 510.270 ;
        RECT 2193.840 196.530 2194.100 196.850 ;
        RECT 2560.000 196.530 2560.260 196.850 ;
        RECT 2560.060 16.990 2560.200 196.530 ;
        RECT 2560.000 16.670 2560.260 16.990 ;
        RECT 2565.980 16.670 2566.240 16.990 ;
        RECT 2566.040 2.400 2566.180 16.670 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.150 451.760 2207.470 451.820 ;
        RECT 2580.670 451.760 2580.990 451.820 ;
        RECT 2207.150 451.620 2580.990 451.760 ;
        RECT 2207.150 451.560 2207.470 451.620 ;
        RECT 2580.670 451.560 2580.990 451.620 ;
      LAYER via ;
        RECT 2207.180 451.560 2207.440 451.820 ;
        RECT 2580.700 451.560 2580.960 451.820 ;
      LAYER met2 ;
        RECT 2207.310 510.340 2207.590 514.000 ;
        RECT 2207.240 510.000 2207.590 510.340 ;
        RECT 2207.240 451.850 2207.380 510.000 ;
        RECT 2207.180 451.530 2207.440 451.850 ;
        RECT 2580.700 451.530 2580.960 451.850 ;
        RECT 2580.760 17.410 2580.900 451.530 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 113.800 593.330 113.860 ;
        RECT 814.270 113.800 814.590 113.860 ;
        RECT 593.010 113.660 814.590 113.800 ;
        RECT 593.010 113.600 593.330 113.660 ;
        RECT 814.270 113.600 814.590 113.660 ;
      LAYER via ;
        RECT 593.040 113.600 593.300 113.860 ;
        RECT 814.300 113.600 814.560 113.860 ;
      LAYER met2 ;
        RECT 591.790 510.410 592.070 514.000 ;
        RECT 591.790 510.270 593.240 510.410 ;
        RECT 591.790 510.000 592.070 510.270 ;
        RECT 593.100 113.890 593.240 510.270 ;
        RECT 593.040 113.570 593.300 113.890 ;
        RECT 814.300 113.570 814.560 113.890 ;
        RECT 814.360 17.410 814.500 113.570 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2223.710 496.980 2224.030 497.040 ;
        RECT 2228.310 496.980 2228.630 497.040 ;
        RECT 2223.710 496.840 2228.630 496.980 ;
        RECT 2223.710 496.780 2224.030 496.840 ;
        RECT 2228.310 496.780 2228.630 496.840 ;
        RECT 2228.310 134.540 2228.630 134.600 ;
        RECT 2601.830 134.540 2602.150 134.600 ;
        RECT 2228.310 134.400 2602.150 134.540 ;
        RECT 2228.310 134.340 2228.630 134.400 ;
        RECT 2601.830 134.340 2602.150 134.400 ;
      LAYER via ;
        RECT 2223.740 496.780 2224.000 497.040 ;
        RECT 2228.340 496.780 2228.600 497.040 ;
        RECT 2228.340 134.340 2228.600 134.600 ;
        RECT 2601.860 134.340 2602.120 134.600 ;
      LAYER met2 ;
        RECT 2223.870 510.340 2224.150 514.000 ;
        RECT 2223.800 510.000 2224.150 510.340 ;
        RECT 2223.800 497.070 2223.940 510.000 ;
        RECT 2223.740 496.750 2224.000 497.070 ;
        RECT 2228.340 496.750 2228.600 497.070 ;
        RECT 2228.400 134.630 2228.540 496.750 ;
        RECT 2228.340 134.310 2228.600 134.630 ;
        RECT 2601.860 134.310 2602.120 134.630 ;
        RECT 2601.920 17.410 2602.060 134.310 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2242.110 141.340 2242.430 141.400 ;
        RECT 2615.170 141.340 2615.490 141.400 ;
        RECT 2242.110 141.200 2615.490 141.340 ;
        RECT 2242.110 141.140 2242.430 141.200 ;
        RECT 2615.170 141.140 2615.490 141.200 ;
      LAYER via ;
        RECT 2242.140 141.140 2242.400 141.400 ;
        RECT 2615.200 141.140 2615.460 141.400 ;
      LAYER met2 ;
        RECT 2239.970 510.410 2240.250 514.000 ;
        RECT 2239.970 510.270 2242.340 510.410 ;
        RECT 2239.970 510.000 2240.250 510.270 ;
        RECT 2242.200 141.430 2242.340 510.270 ;
        RECT 2242.140 141.110 2242.400 141.430 ;
        RECT 2615.200 141.110 2615.460 141.430 ;
        RECT 2615.260 17.410 2615.400 141.110 ;
        RECT 2615.260 17.270 2619.540 17.410 ;
        RECT 2619.400 2.400 2619.540 17.270 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2256.370 496.980 2256.690 497.040 ;
        RECT 2262.810 496.980 2263.130 497.040 ;
        RECT 2256.370 496.840 2263.130 496.980 ;
        RECT 2256.370 496.780 2256.690 496.840 ;
        RECT 2262.810 496.780 2263.130 496.840 ;
        RECT 2262.810 320.860 2263.130 320.920 ;
        RECT 2635.870 320.860 2636.190 320.920 ;
        RECT 2262.810 320.720 2636.190 320.860 ;
        RECT 2262.810 320.660 2263.130 320.720 ;
        RECT 2635.870 320.660 2636.190 320.720 ;
      LAYER via ;
        RECT 2256.400 496.780 2256.660 497.040 ;
        RECT 2262.840 496.780 2263.100 497.040 ;
        RECT 2262.840 320.660 2263.100 320.920 ;
        RECT 2635.900 320.660 2636.160 320.920 ;
      LAYER met2 ;
        RECT 2256.530 510.340 2256.810 514.000 ;
        RECT 2256.460 510.000 2256.810 510.340 ;
        RECT 2256.460 497.070 2256.600 510.000 ;
        RECT 2256.400 496.750 2256.660 497.070 ;
        RECT 2262.840 496.750 2263.100 497.070 ;
        RECT 2262.900 320.950 2263.040 496.750 ;
        RECT 2262.840 320.630 2263.100 320.950 ;
        RECT 2635.900 320.630 2636.160 320.950 ;
        RECT 2635.960 17.410 2636.100 320.630 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2272.470 496.980 2272.790 497.040 ;
        RECT 2276.610 496.980 2276.930 497.040 ;
        RECT 2272.470 496.840 2276.930 496.980 ;
        RECT 2272.470 496.780 2272.790 496.840 ;
        RECT 2276.610 496.780 2276.930 496.840 ;
        RECT 2276.610 258.640 2276.930 258.700 ;
        RECT 2649.670 258.640 2649.990 258.700 ;
        RECT 2276.610 258.500 2649.990 258.640 ;
        RECT 2276.610 258.440 2276.930 258.500 ;
        RECT 2649.670 258.440 2649.990 258.500 ;
      LAYER via ;
        RECT 2272.500 496.780 2272.760 497.040 ;
        RECT 2276.640 496.780 2276.900 497.040 ;
        RECT 2276.640 258.440 2276.900 258.700 ;
        RECT 2649.700 258.440 2649.960 258.700 ;
      LAYER met2 ;
        RECT 2272.630 510.340 2272.910 514.000 ;
        RECT 2272.560 510.000 2272.910 510.340 ;
        RECT 2272.560 497.070 2272.700 510.000 ;
        RECT 2272.500 496.750 2272.760 497.070 ;
        RECT 2276.640 496.750 2276.900 497.070 ;
        RECT 2276.700 258.730 2276.840 496.750 ;
        RECT 2276.640 258.410 2276.900 258.730 ;
        RECT 2649.700 258.410 2649.960 258.730 ;
        RECT 2649.760 17.410 2649.900 258.410 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2290.410 265.440 2290.730 265.500 ;
        RECT 2670.370 265.440 2670.690 265.500 ;
        RECT 2290.410 265.300 2670.690 265.440 ;
        RECT 2290.410 265.240 2290.730 265.300 ;
        RECT 2670.370 265.240 2670.690 265.300 ;
      LAYER via ;
        RECT 2290.440 265.240 2290.700 265.500 ;
        RECT 2670.400 265.240 2670.660 265.500 ;
      LAYER met2 ;
        RECT 2289.190 510.410 2289.470 514.000 ;
        RECT 2289.190 510.270 2290.640 510.410 ;
        RECT 2289.190 510.000 2289.470 510.270 ;
        RECT 2290.500 265.530 2290.640 510.270 ;
        RECT 2290.440 265.210 2290.700 265.530 ;
        RECT 2670.400 265.210 2670.660 265.530 ;
        RECT 2670.460 17.410 2670.600 265.210 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2305.130 503.440 2305.450 503.500 ;
        RECT 2314.790 503.440 2315.110 503.500 ;
        RECT 2305.130 503.300 2315.110 503.440 ;
        RECT 2305.130 503.240 2305.450 503.300 ;
        RECT 2314.790 503.240 2315.110 503.300 ;
        RECT 2314.790 431.360 2315.110 431.420 ;
        RECT 2684.170 431.360 2684.490 431.420 ;
        RECT 2314.790 431.220 2684.490 431.360 ;
        RECT 2314.790 431.160 2315.110 431.220 ;
        RECT 2684.170 431.160 2684.490 431.220 ;
        RECT 2684.170 16.900 2684.490 16.960 ;
        RECT 2690.610 16.900 2690.930 16.960 ;
        RECT 2684.170 16.760 2690.930 16.900 ;
        RECT 2684.170 16.700 2684.490 16.760 ;
        RECT 2690.610 16.700 2690.930 16.760 ;
      LAYER via ;
        RECT 2305.160 503.240 2305.420 503.500 ;
        RECT 2314.820 503.240 2315.080 503.500 ;
        RECT 2314.820 431.160 2315.080 431.420 ;
        RECT 2684.200 431.160 2684.460 431.420 ;
        RECT 2684.200 16.700 2684.460 16.960 ;
        RECT 2690.640 16.700 2690.900 16.960 ;
      LAYER met2 ;
        RECT 2305.290 510.340 2305.570 514.000 ;
        RECT 2305.220 510.000 2305.570 510.340 ;
        RECT 2305.220 503.530 2305.360 510.000 ;
        RECT 2305.160 503.210 2305.420 503.530 ;
        RECT 2314.820 503.210 2315.080 503.530 ;
        RECT 2314.880 431.450 2315.020 503.210 ;
        RECT 2314.820 431.130 2315.080 431.450 ;
        RECT 2684.200 431.130 2684.460 431.450 ;
        RECT 2684.260 16.990 2684.400 431.130 ;
        RECT 2684.200 16.670 2684.460 16.990 ;
        RECT 2690.640 16.670 2690.900 16.990 ;
        RECT 2690.700 2.400 2690.840 16.670 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2324.910 155.280 2325.230 155.340 ;
        RECT 2704.870 155.280 2705.190 155.340 ;
        RECT 2324.910 155.140 2705.190 155.280 ;
        RECT 2324.910 155.080 2325.230 155.140 ;
        RECT 2704.870 155.080 2705.190 155.140 ;
      LAYER via ;
        RECT 2324.940 155.080 2325.200 155.340 ;
        RECT 2704.900 155.080 2705.160 155.340 ;
      LAYER met2 ;
        RECT 2321.850 510.410 2322.130 514.000 ;
        RECT 2321.850 510.270 2325.140 510.410 ;
        RECT 2321.850 510.000 2322.130 510.270 ;
        RECT 2325.000 155.370 2325.140 510.270 ;
        RECT 2324.940 155.050 2325.200 155.370 ;
        RECT 2704.900 155.050 2705.160 155.370 ;
        RECT 2704.960 17.410 2705.100 155.050 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2337.790 424.220 2338.110 424.280 ;
        RECT 2725.570 424.220 2725.890 424.280 ;
        RECT 2337.790 424.080 2725.890 424.220 ;
        RECT 2337.790 424.020 2338.110 424.080 ;
        RECT 2725.570 424.020 2725.890 424.080 ;
      LAYER via ;
        RECT 2337.820 424.020 2338.080 424.280 ;
        RECT 2725.600 424.020 2725.860 424.280 ;
      LAYER met2 ;
        RECT 2337.950 510.340 2338.230 514.000 ;
        RECT 2337.880 510.000 2338.230 510.340 ;
        RECT 2337.880 424.310 2338.020 510.000 ;
        RECT 2337.820 423.990 2338.080 424.310 ;
        RECT 2725.600 423.990 2725.860 424.310 ;
        RECT 2725.660 17.410 2725.800 423.990 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2354.350 496.980 2354.670 497.040 ;
        RECT 2358.950 496.980 2359.270 497.040 ;
        RECT 2354.350 496.840 2359.270 496.980 ;
        RECT 2354.350 496.780 2354.670 496.840 ;
        RECT 2358.950 496.780 2359.270 496.840 ;
        RECT 2358.950 162.080 2359.270 162.140 ;
        RECT 2739.370 162.080 2739.690 162.140 ;
        RECT 2358.950 161.940 2739.690 162.080 ;
        RECT 2358.950 161.880 2359.270 161.940 ;
        RECT 2739.370 161.880 2739.690 161.940 ;
      LAYER via ;
        RECT 2354.380 496.780 2354.640 497.040 ;
        RECT 2358.980 496.780 2359.240 497.040 ;
        RECT 2358.980 161.880 2359.240 162.140 ;
        RECT 2739.400 161.880 2739.660 162.140 ;
      LAYER met2 ;
        RECT 2354.510 510.340 2354.790 514.000 ;
        RECT 2354.440 510.000 2354.790 510.340 ;
        RECT 2354.440 497.070 2354.580 510.000 ;
        RECT 2354.380 496.750 2354.640 497.070 ;
        RECT 2358.980 496.750 2359.240 497.070 ;
        RECT 2359.040 162.170 2359.180 496.750 ;
        RECT 2358.980 161.850 2359.240 162.170 ;
        RECT 2739.400 161.850 2739.660 162.170 ;
        RECT 2739.460 17.410 2739.600 161.850 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2373.210 168.880 2373.530 168.940 ;
        RECT 2760.070 168.880 2760.390 168.940 ;
        RECT 2373.210 168.740 2760.390 168.880 ;
        RECT 2373.210 168.680 2373.530 168.740 ;
        RECT 2760.070 168.680 2760.390 168.740 ;
      LAYER via ;
        RECT 2373.240 168.680 2373.500 168.940 ;
        RECT 2760.100 168.680 2760.360 168.940 ;
      LAYER met2 ;
        RECT 2370.610 510.410 2370.890 514.000 ;
        RECT 2370.610 510.270 2373.440 510.410 ;
        RECT 2370.610 510.000 2370.890 510.270 ;
        RECT 2373.300 168.970 2373.440 510.270 ;
        RECT 2373.240 168.650 2373.500 168.970 ;
        RECT 2760.100 168.650 2760.360 168.970 ;
        RECT 2760.160 17.410 2760.300 168.650 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 607.730 496.980 608.050 497.040 ;
        RECT 613.710 496.980 614.030 497.040 ;
        RECT 607.730 496.840 614.030 496.980 ;
        RECT 607.730 496.780 608.050 496.840 ;
        RECT 613.710 496.780 614.030 496.840 ;
        RECT 613.710 120.600 614.030 120.660 ;
        RECT 835.430 120.600 835.750 120.660 ;
        RECT 613.710 120.460 835.750 120.600 ;
        RECT 613.710 120.400 614.030 120.460 ;
        RECT 835.430 120.400 835.750 120.460 ;
      LAYER via ;
        RECT 607.760 496.780 608.020 497.040 ;
        RECT 613.740 496.780 614.000 497.040 ;
        RECT 613.740 120.400 614.000 120.660 ;
        RECT 835.460 120.400 835.720 120.660 ;
      LAYER met2 ;
        RECT 607.890 510.340 608.170 514.000 ;
        RECT 607.820 510.000 608.170 510.340 ;
        RECT 607.820 497.070 607.960 510.000 ;
        RECT 607.760 496.750 608.020 497.070 ;
        RECT 613.740 496.750 614.000 497.070 ;
        RECT 613.800 120.690 613.940 496.750 ;
        RECT 613.740 120.370 614.000 120.690 ;
        RECT 835.460 120.370 835.720 120.690 ;
        RECT 835.520 2.400 835.660 120.370 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.010 189.620 2387.330 189.680 ;
        RECT 2774.330 189.620 2774.650 189.680 ;
        RECT 2387.010 189.480 2774.650 189.620 ;
        RECT 2387.010 189.420 2387.330 189.480 ;
        RECT 2774.330 189.420 2774.650 189.480 ;
        RECT 2774.330 62.120 2774.650 62.180 ;
        RECT 2779.850 62.120 2780.170 62.180 ;
        RECT 2774.330 61.980 2780.170 62.120 ;
        RECT 2774.330 61.920 2774.650 61.980 ;
        RECT 2779.850 61.920 2780.170 61.980 ;
      LAYER via ;
        RECT 2387.040 189.420 2387.300 189.680 ;
        RECT 2774.360 189.420 2774.620 189.680 ;
        RECT 2774.360 61.920 2774.620 62.180 ;
        RECT 2779.880 61.920 2780.140 62.180 ;
      LAYER met2 ;
        RECT 2386.710 511.090 2386.990 514.000 ;
        RECT 2386.710 510.950 2387.700 511.090 ;
        RECT 2386.710 510.000 2386.990 510.950 ;
        RECT 2387.560 483.210 2387.700 510.950 ;
        RECT 2387.100 483.070 2387.700 483.210 ;
        RECT 2387.100 189.710 2387.240 483.070 ;
        RECT 2387.040 189.390 2387.300 189.710 ;
        RECT 2774.360 189.390 2774.620 189.710 ;
        RECT 2774.420 62.210 2774.560 189.390 ;
        RECT 2774.360 61.890 2774.620 62.210 ;
        RECT 2779.880 61.890 2780.140 62.210 ;
        RECT 2779.940 2.400 2780.080 61.890 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2403.110 503.440 2403.430 503.500 ;
        RECT 2407.710 503.440 2408.030 503.500 ;
        RECT 2403.110 503.300 2408.030 503.440 ;
        RECT 2403.110 503.240 2403.430 503.300 ;
        RECT 2407.710 503.240 2408.030 503.300 ;
        RECT 2407.710 176.020 2408.030 176.080 ;
        RECT 2794.570 176.020 2794.890 176.080 ;
        RECT 2407.710 175.880 2794.890 176.020 ;
        RECT 2407.710 175.820 2408.030 175.880 ;
        RECT 2794.570 175.820 2794.890 175.880 ;
        RECT 2794.570 62.120 2794.890 62.180 ;
        RECT 2797.790 62.120 2798.110 62.180 ;
        RECT 2794.570 61.980 2798.110 62.120 ;
        RECT 2794.570 61.920 2794.890 61.980 ;
        RECT 2797.790 61.920 2798.110 61.980 ;
      LAYER via ;
        RECT 2403.140 503.240 2403.400 503.500 ;
        RECT 2407.740 503.240 2408.000 503.500 ;
        RECT 2407.740 175.820 2408.000 176.080 ;
        RECT 2794.600 175.820 2794.860 176.080 ;
        RECT 2794.600 61.920 2794.860 62.180 ;
        RECT 2797.820 61.920 2798.080 62.180 ;
      LAYER met2 ;
        RECT 2403.270 510.340 2403.550 514.000 ;
        RECT 2403.200 510.000 2403.550 510.340 ;
        RECT 2403.200 503.530 2403.340 510.000 ;
        RECT 2403.140 503.210 2403.400 503.530 ;
        RECT 2407.740 503.210 2408.000 503.530 ;
        RECT 2407.800 176.110 2407.940 503.210 ;
        RECT 2407.740 175.790 2408.000 176.110 ;
        RECT 2794.600 175.790 2794.860 176.110 ;
        RECT 2794.660 62.210 2794.800 175.790 ;
        RECT 2794.600 61.890 2794.860 62.210 ;
        RECT 2797.820 61.890 2798.080 62.210 ;
        RECT 2797.880 2.400 2798.020 61.890 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2421.510 182.820 2421.830 182.880 ;
        RECT 2815.730 182.820 2816.050 182.880 ;
        RECT 2421.510 182.680 2816.050 182.820 ;
        RECT 2421.510 182.620 2421.830 182.680 ;
        RECT 2815.730 182.620 2816.050 182.680 ;
      LAYER via ;
        RECT 2421.540 182.620 2421.800 182.880 ;
        RECT 2815.760 182.620 2816.020 182.880 ;
      LAYER met2 ;
        RECT 2419.370 510.410 2419.650 514.000 ;
        RECT 2419.370 510.270 2421.740 510.410 ;
        RECT 2419.370 510.000 2419.650 510.270 ;
        RECT 2421.600 182.910 2421.740 510.270 ;
        RECT 2421.540 182.590 2421.800 182.910 ;
        RECT 2815.760 182.590 2816.020 182.910 ;
        RECT 2815.820 2.400 2815.960 182.590 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2435.770 496.980 2436.090 497.040 ;
        RECT 2441.750 496.980 2442.070 497.040 ;
        RECT 2435.770 496.840 2442.070 496.980 ;
        RECT 2435.770 496.780 2436.090 496.840 ;
        RECT 2441.750 496.780 2442.070 496.840 ;
        RECT 2441.750 217.160 2442.070 217.220 ;
        RECT 2829.070 217.160 2829.390 217.220 ;
        RECT 2441.750 217.020 2829.390 217.160 ;
        RECT 2441.750 216.960 2442.070 217.020 ;
        RECT 2829.070 216.960 2829.390 217.020 ;
      LAYER via ;
        RECT 2435.800 496.780 2436.060 497.040 ;
        RECT 2441.780 496.780 2442.040 497.040 ;
        RECT 2441.780 216.960 2442.040 217.220 ;
        RECT 2829.100 216.960 2829.360 217.220 ;
      LAYER met2 ;
        RECT 2435.930 510.340 2436.210 514.000 ;
        RECT 2435.860 510.000 2436.210 510.340 ;
        RECT 2435.860 497.070 2436.000 510.000 ;
        RECT 2435.800 496.750 2436.060 497.070 ;
        RECT 2441.780 496.750 2442.040 497.070 ;
        RECT 2441.840 217.250 2441.980 496.750 ;
        RECT 2441.780 216.930 2442.040 217.250 ;
        RECT 2829.100 216.930 2829.360 217.250 ;
        RECT 2829.160 17.410 2829.300 216.930 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2451.870 496.980 2452.190 497.040 ;
        RECT 2456.010 496.980 2456.330 497.040 ;
        RECT 2451.870 496.840 2456.330 496.980 ;
        RECT 2451.870 496.780 2452.190 496.840 ;
        RECT 2456.010 496.780 2456.330 496.840 ;
        RECT 2456.010 417.420 2456.330 417.480 ;
        RECT 2849.770 417.420 2850.090 417.480 ;
        RECT 2456.010 417.280 2850.090 417.420 ;
        RECT 2456.010 417.220 2456.330 417.280 ;
        RECT 2849.770 417.220 2850.090 417.280 ;
      LAYER via ;
        RECT 2451.900 496.780 2452.160 497.040 ;
        RECT 2456.040 496.780 2456.300 497.040 ;
        RECT 2456.040 417.220 2456.300 417.480 ;
        RECT 2849.800 417.220 2850.060 417.480 ;
      LAYER met2 ;
        RECT 2452.030 510.340 2452.310 514.000 ;
        RECT 2451.960 510.000 2452.310 510.340 ;
        RECT 2451.960 497.070 2452.100 510.000 ;
        RECT 2451.900 496.750 2452.160 497.070 ;
        RECT 2456.040 496.750 2456.300 497.070 ;
        RECT 2456.100 417.510 2456.240 496.750 ;
        RECT 2456.040 417.190 2456.300 417.510 ;
        RECT 2849.800 417.190 2850.060 417.510 ;
        RECT 2849.860 17.410 2850.000 417.190 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2469.810 210.360 2470.130 210.420 ;
        RECT 2863.570 210.360 2863.890 210.420 ;
        RECT 2469.810 210.220 2863.890 210.360 ;
        RECT 2469.810 210.160 2470.130 210.220 ;
        RECT 2863.570 210.160 2863.890 210.220 ;
      LAYER via ;
        RECT 2469.840 210.160 2470.100 210.420 ;
        RECT 2863.600 210.160 2863.860 210.420 ;
      LAYER met2 ;
        RECT 2468.590 510.410 2468.870 514.000 ;
        RECT 2468.590 510.270 2470.040 510.410 ;
        RECT 2468.590 510.000 2468.870 510.270 ;
        RECT 2469.900 210.450 2470.040 510.270 ;
        RECT 2469.840 210.130 2470.100 210.450 ;
        RECT 2863.600 210.130 2863.860 210.450 ;
        RECT 2863.660 17.410 2863.800 210.130 ;
        RECT 2863.660 17.270 2869.320 17.410 ;
        RECT 2869.180 2.400 2869.320 17.270 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2484.530 496.980 2484.850 497.040 ;
        RECT 2490.050 496.980 2490.370 497.040 ;
        RECT 2484.530 496.840 2490.370 496.980 ;
        RECT 2484.530 496.780 2484.850 496.840 ;
        RECT 2490.050 496.780 2490.370 496.840 ;
        RECT 2490.050 444.960 2490.370 445.020 ;
        RECT 2873.690 444.960 2874.010 445.020 ;
        RECT 2490.050 444.820 2874.010 444.960 ;
        RECT 2490.050 444.760 2490.370 444.820 ;
        RECT 2873.690 444.760 2874.010 444.820 ;
        RECT 2873.690 19.960 2874.010 20.020 ;
        RECT 2887.030 19.960 2887.350 20.020 ;
        RECT 2873.690 19.820 2887.350 19.960 ;
        RECT 2873.690 19.760 2874.010 19.820 ;
        RECT 2887.030 19.760 2887.350 19.820 ;
      LAYER via ;
        RECT 2484.560 496.780 2484.820 497.040 ;
        RECT 2490.080 496.780 2490.340 497.040 ;
        RECT 2490.080 444.760 2490.340 445.020 ;
        RECT 2873.720 444.760 2873.980 445.020 ;
        RECT 2873.720 19.760 2873.980 20.020 ;
        RECT 2887.060 19.760 2887.320 20.020 ;
      LAYER met2 ;
        RECT 2484.690 510.340 2484.970 514.000 ;
        RECT 2484.620 510.000 2484.970 510.340 ;
        RECT 2484.620 497.070 2484.760 510.000 ;
        RECT 2484.560 496.750 2484.820 497.070 ;
        RECT 2490.080 496.750 2490.340 497.070 ;
        RECT 2490.140 445.050 2490.280 496.750 ;
        RECT 2490.080 444.730 2490.340 445.050 ;
        RECT 2873.720 444.730 2873.980 445.050 ;
        RECT 2873.780 20.050 2873.920 444.730 ;
        RECT 2873.720 19.730 2873.980 20.050 ;
        RECT 2887.060 19.730 2887.320 20.050 ;
        RECT 2887.120 2.400 2887.260 19.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2504.310 58.720 2504.630 58.780 ;
        RECT 2905.430 58.720 2905.750 58.780 ;
        RECT 2504.310 58.580 2905.750 58.720 ;
        RECT 2504.310 58.520 2504.630 58.580 ;
        RECT 2905.430 58.520 2905.750 58.580 ;
      LAYER via ;
        RECT 2504.340 58.520 2504.600 58.780 ;
        RECT 2905.460 58.520 2905.720 58.780 ;
      LAYER met2 ;
        RECT 2501.250 510.410 2501.530 514.000 ;
        RECT 2501.250 510.270 2504.540 510.410 ;
        RECT 2501.250 510.000 2501.530 510.270 ;
        RECT 2504.400 58.810 2504.540 510.270 ;
        RECT 2504.340 58.490 2504.600 58.810 ;
        RECT 2905.460 58.490 2905.720 58.810 ;
        RECT 2905.520 3.130 2905.660 58.490 ;
        RECT 2905.060 2.990 2905.660 3.130 ;
        RECT 2905.060 2.400 2905.200 2.990 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 128.080 627.830 128.140 ;
        RECT 848.770 128.080 849.090 128.140 ;
        RECT 627.510 127.940 849.090 128.080 ;
        RECT 627.510 127.880 627.830 127.940 ;
        RECT 848.770 127.880 849.090 127.940 ;
      LAYER via ;
        RECT 627.540 127.880 627.800 128.140 ;
        RECT 848.800 127.880 849.060 128.140 ;
      LAYER met2 ;
        RECT 624.450 510.410 624.730 514.000 ;
        RECT 624.450 510.270 627.740 510.410 ;
        RECT 624.450 510.000 624.730 510.270 ;
        RECT 627.600 128.170 627.740 510.270 ;
        RECT 627.540 127.850 627.800 128.170 ;
        RECT 848.800 127.850 849.060 128.170 ;
        RECT 848.860 17.410 849.000 127.850 ;
        RECT 848.860 17.270 853.140 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 134.880 641.630 134.940 ;
        RECT 869.470 134.880 869.790 134.940 ;
        RECT 641.310 134.740 869.790 134.880 ;
        RECT 641.310 134.680 641.630 134.740 ;
        RECT 869.470 134.680 869.790 134.740 ;
      LAYER via ;
        RECT 641.340 134.680 641.600 134.940 ;
        RECT 869.500 134.680 869.760 134.940 ;
      LAYER met2 ;
        RECT 640.550 510.410 640.830 514.000 ;
        RECT 640.550 510.270 641.540 510.410 ;
        RECT 640.550 510.000 640.830 510.270 ;
        RECT 641.400 134.970 641.540 510.270 ;
        RECT 641.340 134.650 641.600 134.970 ;
        RECT 869.500 134.650 869.760 134.970 ;
        RECT 869.560 17.410 869.700 134.650 ;
        RECT 869.560 17.270 871.080 17.410 ;
        RECT 870.940 2.400 871.080 17.270 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 496.980 657.270 497.040 ;
        RECT 662.010 496.980 662.330 497.040 ;
        RECT 656.950 496.840 662.330 496.980 ;
        RECT 656.950 496.780 657.270 496.840 ;
        RECT 662.010 496.780 662.330 496.840 ;
        RECT 662.010 141.340 662.330 141.400 ;
        RECT 883.270 141.340 883.590 141.400 ;
        RECT 662.010 141.200 883.590 141.340 ;
        RECT 662.010 141.140 662.330 141.200 ;
        RECT 883.270 141.140 883.590 141.200 ;
      LAYER via ;
        RECT 656.980 496.780 657.240 497.040 ;
        RECT 662.040 496.780 662.300 497.040 ;
        RECT 662.040 141.140 662.300 141.400 ;
        RECT 883.300 141.140 883.560 141.400 ;
      LAYER met2 ;
        RECT 657.110 510.340 657.390 514.000 ;
        RECT 657.040 510.000 657.390 510.340 ;
        RECT 657.040 497.070 657.180 510.000 ;
        RECT 656.980 496.750 657.240 497.070 ;
        RECT 662.040 496.750 662.300 497.070 ;
        RECT 662.100 141.430 662.240 496.750 ;
        RECT 662.040 141.110 662.300 141.430 ;
        RECT 883.300 141.110 883.560 141.430 ;
        RECT 883.360 17.410 883.500 141.110 ;
        RECT 883.360 17.270 889.020 17.410 ;
        RECT 888.880 2.400 889.020 17.270 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 148.480 676.130 148.540 ;
        RECT 903.970 148.480 904.290 148.540 ;
        RECT 675.810 148.340 904.290 148.480 ;
        RECT 675.810 148.280 676.130 148.340 ;
        RECT 903.970 148.280 904.290 148.340 ;
      LAYER via ;
        RECT 675.840 148.280 676.100 148.540 ;
        RECT 904.000 148.280 904.260 148.540 ;
      LAYER met2 ;
        RECT 673.210 510.410 673.490 514.000 ;
        RECT 673.210 510.270 676.040 510.410 ;
        RECT 673.210 510.000 673.490 510.270 ;
        RECT 675.900 148.570 676.040 510.270 ;
        RECT 675.840 148.250 676.100 148.570 ;
        RECT 904.000 148.250 904.260 148.570 ;
        RECT 904.060 17.410 904.200 148.250 ;
        RECT 904.060 17.270 906.960 17.410 ;
        RECT 906.820 2.400 906.960 17.270 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.610 155.280 689.930 155.340 ;
        RECT 917.770 155.280 918.090 155.340 ;
        RECT 689.610 155.140 918.090 155.280 ;
        RECT 689.610 155.080 689.930 155.140 ;
        RECT 917.770 155.080 918.090 155.140 ;
        RECT 917.770 17.580 918.090 17.640 ;
        RECT 924.210 17.580 924.530 17.640 ;
        RECT 917.770 17.440 924.530 17.580 ;
        RECT 917.770 17.380 918.090 17.440 ;
        RECT 924.210 17.380 924.530 17.440 ;
      LAYER via ;
        RECT 689.640 155.080 689.900 155.340 ;
        RECT 917.800 155.080 918.060 155.340 ;
        RECT 917.800 17.380 918.060 17.640 ;
        RECT 924.240 17.380 924.500 17.640 ;
      LAYER met2 ;
        RECT 689.770 510.340 690.050 514.000 ;
        RECT 689.700 510.000 690.050 510.340 ;
        RECT 689.700 155.370 689.840 510.000 ;
        RECT 689.640 155.050 689.900 155.370 ;
        RECT 917.800 155.050 918.060 155.370 ;
        RECT 917.860 17.670 918.000 155.050 ;
        RECT 917.800 17.350 918.060 17.670 ;
        RECT 924.240 17.350 924.500 17.670 ;
        RECT 924.300 2.400 924.440 17.350 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 705.710 496.980 706.030 497.040 ;
        RECT 710.310 496.980 710.630 497.040 ;
        RECT 705.710 496.840 710.630 496.980 ;
        RECT 705.710 496.780 706.030 496.840 ;
        RECT 710.310 496.780 710.630 496.840 ;
        RECT 710.310 162.420 710.630 162.480 ;
        RECT 938.470 162.420 938.790 162.480 ;
        RECT 710.310 162.280 938.790 162.420 ;
        RECT 710.310 162.220 710.630 162.280 ;
        RECT 938.470 162.220 938.790 162.280 ;
      LAYER via ;
        RECT 705.740 496.780 706.000 497.040 ;
        RECT 710.340 496.780 710.600 497.040 ;
        RECT 710.340 162.220 710.600 162.480 ;
        RECT 938.500 162.220 938.760 162.480 ;
      LAYER met2 ;
        RECT 705.870 510.340 706.150 514.000 ;
        RECT 705.800 510.000 706.150 510.340 ;
        RECT 705.800 497.070 705.940 510.000 ;
        RECT 705.740 496.750 706.000 497.070 ;
        RECT 710.340 496.750 710.600 497.070 ;
        RECT 710.400 162.510 710.540 496.750 ;
        RECT 710.340 162.190 710.600 162.510 ;
        RECT 938.500 162.190 938.760 162.510 ;
        RECT 938.560 17.410 938.700 162.190 ;
        RECT 938.560 17.270 942.380 17.410 ;
        RECT 942.240 2.400 942.380 17.270 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 724.110 169.220 724.430 169.280 ;
        RECT 959.170 169.220 959.490 169.280 ;
        RECT 724.110 169.080 959.490 169.220 ;
        RECT 724.110 169.020 724.430 169.080 ;
        RECT 959.170 169.020 959.490 169.080 ;
      LAYER via ;
        RECT 724.140 169.020 724.400 169.280 ;
        RECT 959.200 169.020 959.460 169.280 ;
      LAYER met2 ;
        RECT 722.430 510.410 722.710 514.000 ;
        RECT 722.430 510.270 724.340 510.410 ;
        RECT 722.430 510.000 722.710 510.270 ;
        RECT 724.200 169.310 724.340 510.270 ;
        RECT 724.140 168.990 724.400 169.310 ;
        RECT 959.200 168.990 959.460 169.310 ;
        RECT 959.260 17.410 959.400 168.990 ;
        RECT 959.260 17.270 960.320 17.410 ;
        RECT 960.180 2.400 960.320 17.270 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 738.370 493.240 738.690 493.300 ;
        RECT 972.970 493.240 973.290 493.300 ;
        RECT 738.370 493.100 973.290 493.240 ;
        RECT 738.370 493.040 738.690 493.100 ;
        RECT 972.970 493.040 973.290 493.100 ;
      LAYER via ;
        RECT 738.400 493.040 738.660 493.300 ;
        RECT 973.000 493.040 973.260 493.300 ;
      LAYER met2 ;
        RECT 738.530 510.340 738.810 514.000 ;
        RECT 738.460 510.000 738.810 510.340 ;
        RECT 738.460 493.330 738.600 510.000 ;
        RECT 738.400 493.010 738.660 493.330 ;
        RECT 973.000 493.010 973.260 493.330 ;
        RECT 973.060 17.410 973.200 493.010 ;
        RECT 973.060 17.270 978.260 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 444.430 503.440 444.750 503.500 ;
        RECT 448.110 503.440 448.430 503.500 ;
        RECT 444.430 503.300 448.430 503.440 ;
        RECT 444.430 503.240 444.750 503.300 ;
        RECT 448.110 503.240 448.430 503.300 ;
        RECT 448.110 141.340 448.430 141.400 ;
        RECT 655.570 141.340 655.890 141.400 ;
        RECT 448.110 141.200 655.890 141.340 ;
        RECT 448.110 141.140 448.430 141.200 ;
        RECT 655.570 141.140 655.890 141.200 ;
        RECT 655.570 2.960 655.890 3.020 ;
        RECT 656.950 2.960 657.270 3.020 ;
        RECT 655.570 2.820 657.270 2.960 ;
        RECT 655.570 2.760 655.890 2.820 ;
        RECT 656.950 2.760 657.270 2.820 ;
      LAYER via ;
        RECT 444.460 503.240 444.720 503.500 ;
        RECT 448.140 503.240 448.400 503.500 ;
        RECT 448.140 141.140 448.400 141.400 ;
        RECT 655.600 141.140 655.860 141.400 ;
        RECT 655.600 2.760 655.860 3.020 ;
        RECT 656.980 2.760 657.240 3.020 ;
      LAYER met2 ;
        RECT 444.590 510.340 444.870 514.000 ;
        RECT 444.520 510.000 444.870 510.340 ;
        RECT 444.520 503.530 444.660 510.000 ;
        RECT 444.460 503.210 444.720 503.530 ;
        RECT 448.140 503.210 448.400 503.530 ;
        RECT 448.200 141.430 448.340 503.210 ;
        RECT 448.140 141.110 448.400 141.430 ;
        RECT 655.600 141.110 655.860 141.430 ;
        RECT 655.660 3.050 655.800 141.110 ;
        RECT 655.600 2.730 655.860 3.050 ;
        RECT 656.980 2.730 657.240 3.050 ;
        RECT 657.040 2.400 657.180 2.730 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 758.610 176.020 758.930 176.080 ;
        RECT 993.670 176.020 993.990 176.080 ;
        RECT 758.610 175.880 993.990 176.020 ;
        RECT 758.610 175.820 758.930 175.880 ;
        RECT 993.670 175.820 993.990 175.880 ;
      LAYER via ;
        RECT 758.640 175.820 758.900 176.080 ;
        RECT 993.700 175.820 993.960 176.080 ;
      LAYER met2 ;
        RECT 755.090 510.410 755.370 514.000 ;
        RECT 755.090 510.270 758.840 510.410 ;
        RECT 755.090 510.000 755.370 510.270 ;
        RECT 758.700 176.110 758.840 510.270 ;
        RECT 758.640 175.790 758.900 176.110 ;
        RECT 993.700 175.790 993.960 176.110 ;
        RECT 993.760 17.410 993.900 175.790 ;
        RECT 993.760 17.270 996.200 17.410 ;
        RECT 996.060 2.400 996.200 17.270 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 772.410 183.160 772.730 183.220 ;
        RECT 1007.470 183.160 1007.790 183.220 ;
        RECT 772.410 183.020 1007.790 183.160 ;
        RECT 772.410 182.960 772.730 183.020 ;
        RECT 1007.470 182.960 1007.790 183.020 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 1013.450 17.920 1013.770 17.980 ;
        RECT 1007.470 17.780 1013.770 17.920 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
        RECT 1013.450 17.720 1013.770 17.780 ;
      LAYER via ;
        RECT 772.440 182.960 772.700 183.220 ;
        RECT 1007.500 182.960 1007.760 183.220 ;
        RECT 1007.500 17.720 1007.760 17.980 ;
        RECT 1013.480 17.720 1013.740 17.980 ;
      LAYER met2 ;
        RECT 771.190 510.410 771.470 514.000 ;
        RECT 771.190 510.270 772.640 510.410 ;
        RECT 771.190 510.000 771.470 510.270 ;
        RECT 772.500 183.250 772.640 510.270 ;
        RECT 772.440 182.930 772.700 183.250 ;
        RECT 1007.500 182.930 1007.760 183.250 ;
        RECT 1007.560 18.010 1007.700 182.930 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 1013.480 17.690 1013.740 18.010 ;
        RECT 1013.540 2.400 1013.680 17.690 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 787.590 496.980 787.910 497.040 ;
        RECT 793.110 496.980 793.430 497.040 ;
        RECT 787.590 496.840 793.430 496.980 ;
        RECT 787.590 496.780 787.910 496.840 ;
        RECT 793.110 496.780 793.430 496.840 ;
        RECT 793.110 189.620 793.430 189.680 ;
        RECT 1028.170 189.620 1028.490 189.680 ;
        RECT 793.110 189.480 1028.490 189.620 ;
        RECT 793.110 189.420 793.430 189.480 ;
        RECT 1028.170 189.420 1028.490 189.480 ;
      LAYER via ;
        RECT 787.620 496.780 787.880 497.040 ;
        RECT 793.140 496.780 793.400 497.040 ;
        RECT 793.140 189.420 793.400 189.680 ;
        RECT 1028.200 189.420 1028.460 189.680 ;
      LAYER met2 ;
        RECT 787.750 510.340 788.030 514.000 ;
        RECT 787.680 510.000 788.030 510.340 ;
        RECT 787.680 497.070 787.820 510.000 ;
        RECT 787.620 496.750 787.880 497.070 ;
        RECT 793.140 496.750 793.400 497.070 ;
        RECT 793.200 189.710 793.340 496.750 ;
        RECT 793.140 189.390 793.400 189.710 ;
        RECT 1028.200 189.390 1028.460 189.710 ;
        RECT 1028.260 17.410 1028.400 189.390 ;
        RECT 1028.260 17.270 1031.620 17.410 ;
        RECT 1031.480 2.400 1031.620 17.270 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 806.910 114.140 807.230 114.200 ;
        RECT 1049.330 114.140 1049.650 114.200 ;
        RECT 806.910 114.000 1049.650 114.140 ;
        RECT 806.910 113.940 807.230 114.000 ;
        RECT 1049.330 113.940 1049.650 114.000 ;
      LAYER via ;
        RECT 806.940 113.940 807.200 114.200 ;
        RECT 1049.360 113.940 1049.620 114.200 ;
      LAYER met2 ;
        RECT 803.850 510.410 804.130 514.000 ;
        RECT 803.850 510.270 807.140 510.410 ;
        RECT 803.850 510.000 804.130 510.270 ;
        RECT 807.000 114.230 807.140 510.270 ;
        RECT 806.940 113.910 807.200 114.230 ;
        RECT 1049.360 113.910 1049.620 114.230 ;
        RECT 1049.420 2.400 1049.560 113.910 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 820.710 237.900 821.030 237.960 ;
        RECT 1062.670 237.900 1062.990 237.960 ;
        RECT 820.710 237.760 1062.990 237.900 ;
        RECT 820.710 237.700 821.030 237.760 ;
        RECT 1062.670 237.700 1062.990 237.760 ;
      LAYER via ;
        RECT 820.740 237.700 821.000 237.960 ;
        RECT 1062.700 237.700 1062.960 237.960 ;
      LAYER met2 ;
        RECT 819.950 510.410 820.230 514.000 ;
        RECT 819.950 510.270 820.940 510.410 ;
        RECT 819.950 510.000 820.230 510.270 ;
        RECT 820.800 237.990 820.940 510.270 ;
        RECT 820.740 237.670 821.000 237.990 ;
        RECT 1062.700 237.670 1062.960 237.990 ;
        RECT 1062.760 17.410 1062.900 237.670 ;
        RECT 1062.760 17.270 1067.500 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 836.350 496.980 836.670 497.040 ;
        RECT 841.410 496.980 841.730 497.040 ;
        RECT 836.350 496.840 841.730 496.980 ;
        RECT 836.350 496.780 836.670 496.840 ;
        RECT 841.410 496.780 841.730 496.840 ;
        RECT 841.410 127.740 841.730 127.800 ;
        RECT 1083.370 127.740 1083.690 127.800 ;
        RECT 841.410 127.600 1083.690 127.740 ;
        RECT 841.410 127.540 841.730 127.600 ;
        RECT 1083.370 127.540 1083.690 127.600 ;
      LAYER via ;
        RECT 836.380 496.780 836.640 497.040 ;
        RECT 841.440 496.780 841.700 497.040 ;
        RECT 841.440 127.540 841.700 127.800 ;
        RECT 1083.400 127.540 1083.660 127.800 ;
      LAYER met2 ;
        RECT 836.510 510.340 836.790 514.000 ;
        RECT 836.440 510.000 836.790 510.340 ;
        RECT 836.440 497.070 836.580 510.000 ;
        RECT 836.380 496.750 836.640 497.070 ;
        RECT 841.440 496.750 841.700 497.070 ;
        RECT 841.500 127.830 841.640 496.750 ;
        RECT 841.440 127.510 841.700 127.830 ;
        RECT 1083.400 127.510 1083.660 127.830 ;
        RECT 1083.460 17.410 1083.600 127.510 ;
        RECT 1083.460 17.270 1085.440 17.410 ;
        RECT 1085.300 2.400 1085.440 17.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 134.540 855.530 134.600 ;
        RECT 1097.170 134.540 1097.490 134.600 ;
        RECT 855.210 134.400 1097.490 134.540 ;
        RECT 855.210 134.340 855.530 134.400 ;
        RECT 1097.170 134.340 1097.490 134.400 ;
      LAYER via ;
        RECT 855.240 134.340 855.500 134.600 ;
        RECT 1097.200 134.340 1097.460 134.600 ;
      LAYER met2 ;
        RECT 852.610 510.410 852.890 514.000 ;
        RECT 852.610 510.270 855.440 510.410 ;
        RECT 852.610 510.000 852.890 510.270 ;
        RECT 855.300 134.630 855.440 510.270 ;
        RECT 855.240 134.310 855.500 134.630 ;
        RECT 1097.200 134.310 1097.460 134.630 ;
        RECT 1097.260 17.410 1097.400 134.310 ;
        RECT 1097.260 17.270 1102.920 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 868.550 203.560 868.870 203.620 ;
        RECT 1117.870 203.560 1118.190 203.620 ;
        RECT 868.550 203.420 1118.190 203.560 ;
        RECT 868.550 203.360 868.870 203.420 ;
        RECT 1117.870 203.360 1118.190 203.420 ;
      LAYER via ;
        RECT 868.580 203.360 868.840 203.620 ;
        RECT 1117.900 203.360 1118.160 203.620 ;
      LAYER met2 ;
        RECT 869.170 510.410 869.450 514.000 ;
        RECT 868.640 510.270 869.450 510.410 ;
        RECT 868.640 203.650 868.780 510.270 ;
        RECT 869.170 510.000 869.450 510.270 ;
        RECT 868.580 203.330 868.840 203.650 ;
        RECT 1117.900 203.330 1118.160 203.650 ;
        RECT 1117.960 17.410 1118.100 203.330 ;
        RECT 1117.960 17.270 1120.860 17.410 ;
        RECT 1120.720 2.400 1120.860 17.270 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 885.110 496.980 885.430 497.040 ;
        RECT 889.710 496.980 890.030 497.040 ;
        RECT 885.110 496.840 890.030 496.980 ;
        RECT 885.110 496.780 885.430 496.840 ;
        RECT 889.710 496.780 890.030 496.840 ;
        RECT 889.710 141.340 890.030 141.400 ;
        RECT 1139.030 141.340 1139.350 141.400 ;
        RECT 889.710 141.200 1139.350 141.340 ;
        RECT 889.710 141.140 890.030 141.200 ;
        RECT 1139.030 141.140 1139.350 141.200 ;
      LAYER via ;
        RECT 885.140 496.780 885.400 497.040 ;
        RECT 889.740 496.780 890.000 497.040 ;
        RECT 889.740 141.140 890.000 141.400 ;
        RECT 1139.060 141.140 1139.320 141.400 ;
      LAYER met2 ;
        RECT 885.270 510.340 885.550 514.000 ;
        RECT 885.200 510.000 885.550 510.340 ;
        RECT 885.200 497.070 885.340 510.000 ;
        RECT 885.140 496.750 885.400 497.070 ;
        RECT 889.740 496.750 890.000 497.070 ;
        RECT 889.800 141.430 889.940 496.750 ;
        RECT 889.740 141.110 890.000 141.430 ;
        RECT 1139.060 141.110 1139.320 141.430 ;
        RECT 1139.120 17.410 1139.260 141.110 ;
        RECT 1138.660 17.270 1139.260 17.410 ;
        RECT 1138.660 2.400 1138.800 17.270 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 903.510 148.140 903.830 148.200 ;
        RECT 1152.370 148.140 1152.690 148.200 ;
        RECT 903.510 148.000 1152.690 148.140 ;
        RECT 903.510 147.940 903.830 148.000 ;
        RECT 1152.370 147.940 1152.690 148.000 ;
      LAYER via ;
        RECT 903.540 147.940 903.800 148.200 ;
        RECT 1152.400 147.940 1152.660 148.200 ;
      LAYER met2 ;
        RECT 901.830 510.410 902.110 514.000 ;
        RECT 901.830 510.270 903.740 510.410 ;
        RECT 901.830 510.000 902.110 510.270 ;
        RECT 903.600 148.230 903.740 510.270 ;
        RECT 903.540 147.910 903.800 148.230 ;
        RECT 1152.400 147.910 1152.660 148.230 ;
        RECT 1152.460 18.090 1152.600 147.910 ;
        RECT 1152.460 17.950 1156.740 18.090 ;
        RECT 1156.600 2.400 1156.740 17.950 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 461.450 148.140 461.770 148.200 ;
        RECT 669.370 148.140 669.690 148.200 ;
        RECT 461.450 148.000 669.690 148.140 ;
        RECT 461.450 147.940 461.770 148.000 ;
        RECT 669.370 147.940 669.690 148.000 ;
      LAYER via ;
        RECT 461.480 147.940 461.740 148.200 ;
        RECT 669.400 147.940 669.660 148.200 ;
      LAYER met2 ;
        RECT 461.150 511.090 461.430 514.000 ;
        RECT 461.150 510.950 462.140 511.090 ;
        RECT 461.150 510.000 461.430 510.950 ;
        RECT 462.000 503.610 462.140 510.950 ;
        RECT 461.540 503.470 462.140 503.610 ;
        RECT 461.540 148.230 461.680 503.470 ;
        RECT 461.480 147.910 461.740 148.230 ;
        RECT 669.400 147.910 669.660 148.230 ;
        RECT 669.460 17.410 669.600 147.910 ;
        RECT 669.460 17.270 674.660 17.410 ;
        RECT 674.520 2.400 674.660 17.270 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 917.770 496.980 918.090 497.040 ;
        RECT 927.890 496.980 928.210 497.040 ;
        RECT 917.770 496.840 928.210 496.980 ;
        RECT 917.770 496.780 918.090 496.840 ;
        RECT 927.890 496.780 928.210 496.840 ;
        RECT 927.890 155.280 928.210 155.340 ;
        RECT 1173.070 155.280 1173.390 155.340 ;
        RECT 927.890 155.140 1173.390 155.280 ;
        RECT 927.890 155.080 928.210 155.140 ;
        RECT 1173.070 155.080 1173.390 155.140 ;
      LAYER via ;
        RECT 917.800 496.780 918.060 497.040 ;
        RECT 927.920 496.780 928.180 497.040 ;
        RECT 927.920 155.080 928.180 155.340 ;
        RECT 1173.100 155.080 1173.360 155.340 ;
      LAYER met2 ;
        RECT 917.930 510.340 918.210 514.000 ;
        RECT 917.860 510.000 918.210 510.340 ;
        RECT 917.860 497.070 918.000 510.000 ;
        RECT 917.800 496.750 918.060 497.070 ;
        RECT 927.920 496.750 928.180 497.070 ;
        RECT 927.980 155.370 928.120 496.750 ;
        RECT 927.920 155.050 928.180 155.370 ;
        RECT 1173.100 155.050 1173.360 155.370 ;
        RECT 1173.160 17.410 1173.300 155.050 ;
        RECT 1173.160 17.270 1174.220 17.410 ;
        RECT 1174.080 2.400 1174.220 17.270 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 938.010 162.080 938.330 162.140 ;
        RECT 1186.870 162.080 1187.190 162.140 ;
        RECT 938.010 161.940 1187.190 162.080 ;
        RECT 938.010 161.880 938.330 161.940 ;
        RECT 1186.870 161.880 1187.190 161.940 ;
      LAYER via ;
        RECT 938.040 161.880 938.300 162.140 ;
        RECT 1186.900 161.880 1187.160 162.140 ;
      LAYER met2 ;
        RECT 934.490 510.410 934.770 514.000 ;
        RECT 934.490 510.270 938.240 510.410 ;
        RECT 934.490 510.000 934.770 510.270 ;
        RECT 938.100 162.170 938.240 510.270 ;
        RECT 938.040 161.850 938.300 162.170 ;
        RECT 1186.900 161.850 1187.160 162.170 ;
        RECT 1186.960 17.410 1187.100 161.850 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 951.810 168.880 952.130 168.940 ;
        RECT 1207.570 168.880 1207.890 168.940 ;
        RECT 951.810 168.740 1207.890 168.880 ;
        RECT 951.810 168.680 952.130 168.740 ;
        RECT 1207.570 168.680 1207.890 168.740 ;
      LAYER via ;
        RECT 951.840 168.680 952.100 168.940 ;
        RECT 1207.600 168.680 1207.860 168.940 ;
      LAYER met2 ;
        RECT 950.590 510.410 950.870 514.000 ;
        RECT 950.590 510.270 952.040 510.410 ;
        RECT 950.590 510.000 950.870 510.270 ;
        RECT 951.900 168.970 952.040 510.270 ;
        RECT 951.840 168.650 952.100 168.970 ;
        RECT 1207.600 168.650 1207.860 168.970 ;
        RECT 1207.660 17.410 1207.800 168.650 ;
        RECT 1207.660 17.270 1210.100 17.410 ;
        RECT 1209.960 2.400 1210.100 17.270 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 966.990 496.980 967.310 497.040 ;
        RECT 972.510 496.980 972.830 497.040 ;
        RECT 966.990 496.840 972.830 496.980 ;
        RECT 966.990 496.780 967.310 496.840 ;
        RECT 972.510 496.780 972.830 496.840 ;
        RECT 972.510 217.160 972.830 217.220 ;
        RECT 1221.370 217.160 1221.690 217.220 ;
        RECT 972.510 217.020 1221.690 217.160 ;
        RECT 972.510 216.960 972.830 217.020 ;
        RECT 1221.370 216.960 1221.690 217.020 ;
        RECT 1221.370 17.580 1221.690 17.640 ;
        RECT 1227.810 17.580 1228.130 17.640 ;
        RECT 1221.370 17.440 1228.130 17.580 ;
        RECT 1221.370 17.380 1221.690 17.440 ;
        RECT 1227.810 17.380 1228.130 17.440 ;
      LAYER via ;
        RECT 967.020 496.780 967.280 497.040 ;
        RECT 972.540 496.780 972.800 497.040 ;
        RECT 972.540 216.960 972.800 217.220 ;
        RECT 1221.400 216.960 1221.660 217.220 ;
        RECT 1221.400 17.380 1221.660 17.640 ;
        RECT 1227.840 17.380 1228.100 17.640 ;
      LAYER met2 ;
        RECT 967.150 510.340 967.430 514.000 ;
        RECT 967.080 510.000 967.430 510.340 ;
        RECT 967.080 497.070 967.220 510.000 ;
        RECT 967.020 496.750 967.280 497.070 ;
        RECT 972.540 496.750 972.800 497.070 ;
        RECT 972.600 217.250 972.740 496.750 ;
        RECT 972.540 216.930 972.800 217.250 ;
        RECT 1221.400 216.930 1221.660 217.250 ;
        RECT 1221.460 17.670 1221.600 216.930 ;
        RECT 1221.400 17.350 1221.660 17.670 ;
        RECT 1227.840 17.350 1228.100 17.670 ;
        RECT 1227.900 2.400 1228.040 17.350 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 986.310 231.100 986.630 231.160 ;
        RECT 1242.070 231.100 1242.390 231.160 ;
        RECT 986.310 230.960 1242.390 231.100 ;
        RECT 986.310 230.900 986.630 230.960 ;
        RECT 1242.070 230.900 1242.390 230.960 ;
      LAYER via ;
        RECT 986.340 230.900 986.600 231.160 ;
        RECT 1242.100 230.900 1242.360 231.160 ;
      LAYER met2 ;
        RECT 983.250 510.410 983.530 514.000 ;
        RECT 983.250 510.270 986.540 510.410 ;
        RECT 983.250 510.000 983.530 510.270 ;
        RECT 986.400 231.190 986.540 510.270 ;
        RECT 986.340 230.870 986.600 231.190 ;
        RECT 1242.100 230.870 1242.360 231.190 ;
        RECT 1242.160 17.410 1242.300 230.870 ;
        RECT 1242.160 17.270 1245.980 17.410 ;
        RECT 1245.840 2.400 1245.980 17.270 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 999.650 176.020 999.970 176.080 ;
        RECT 1263.230 176.020 1263.550 176.080 ;
        RECT 999.650 175.880 1263.550 176.020 ;
        RECT 999.650 175.820 999.970 175.880 ;
        RECT 1263.230 175.820 1263.550 175.880 ;
      LAYER via ;
        RECT 999.680 175.820 999.940 176.080 ;
        RECT 1263.260 175.820 1263.520 176.080 ;
      LAYER met2 ;
        RECT 999.810 510.340 1000.090 514.000 ;
        RECT 999.740 510.000 1000.090 510.340 ;
        RECT 999.740 176.110 999.880 510.000 ;
        RECT 999.680 175.790 999.940 176.110 ;
        RECT 1263.260 175.790 1263.520 176.110 ;
        RECT 1263.320 2.400 1263.460 175.790 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1015.750 496.980 1016.070 497.040 ;
        RECT 1020.810 496.980 1021.130 497.040 ;
        RECT 1015.750 496.840 1021.130 496.980 ;
        RECT 1015.750 496.780 1016.070 496.840 ;
        RECT 1020.810 496.780 1021.130 496.840 ;
        RECT 1020.810 113.800 1021.130 113.860 ;
        RECT 1276.570 113.800 1276.890 113.860 ;
        RECT 1020.810 113.660 1276.890 113.800 ;
        RECT 1020.810 113.600 1021.130 113.660 ;
        RECT 1276.570 113.600 1276.890 113.660 ;
      LAYER via ;
        RECT 1015.780 496.780 1016.040 497.040 ;
        RECT 1020.840 496.780 1021.100 497.040 ;
        RECT 1020.840 113.600 1021.100 113.860 ;
        RECT 1276.600 113.600 1276.860 113.860 ;
      LAYER met2 ;
        RECT 1015.910 510.340 1016.190 514.000 ;
        RECT 1015.840 510.000 1016.190 510.340 ;
        RECT 1015.840 497.070 1015.980 510.000 ;
        RECT 1015.780 496.750 1016.040 497.070 ;
        RECT 1020.840 496.750 1021.100 497.070 ;
        RECT 1020.900 113.890 1021.040 496.750 ;
        RECT 1020.840 113.570 1021.100 113.890 ;
        RECT 1276.600 113.570 1276.860 113.890 ;
        RECT 1276.660 17.410 1276.800 113.570 ;
        RECT 1276.660 17.270 1281.400 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 189.620 1034.930 189.680 ;
        RECT 1297.270 189.620 1297.590 189.680 ;
        RECT 1034.610 189.480 1297.590 189.620 ;
        RECT 1034.610 189.420 1034.930 189.480 ;
        RECT 1297.270 189.420 1297.590 189.480 ;
      LAYER via ;
        RECT 1034.640 189.420 1034.900 189.680 ;
        RECT 1297.300 189.420 1297.560 189.680 ;
      LAYER met2 ;
        RECT 1032.470 510.410 1032.750 514.000 ;
        RECT 1032.470 510.270 1034.840 510.410 ;
        RECT 1032.470 510.000 1032.750 510.270 ;
        RECT 1034.700 189.710 1034.840 510.270 ;
        RECT 1034.640 189.390 1034.900 189.710 ;
        RECT 1297.300 189.390 1297.560 189.710 ;
        RECT 1297.360 17.410 1297.500 189.390 ;
        RECT 1297.360 17.270 1299.340 17.410 ;
        RECT 1299.200 2.400 1299.340 17.270 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1047.950 251.840 1048.270 251.900 ;
        RECT 1311.070 251.840 1311.390 251.900 ;
        RECT 1047.950 251.700 1311.390 251.840 ;
        RECT 1047.950 251.640 1048.270 251.700 ;
        RECT 1311.070 251.640 1311.390 251.700 ;
        RECT 1311.070 17.920 1311.390 17.980 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1311.070 17.780 1317.370 17.920 ;
        RECT 1311.070 17.720 1311.390 17.780 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
      LAYER via ;
        RECT 1047.980 251.640 1048.240 251.900 ;
        RECT 1311.100 251.640 1311.360 251.900 ;
        RECT 1311.100 17.720 1311.360 17.980 ;
        RECT 1317.080 17.720 1317.340 17.980 ;
      LAYER met2 ;
        RECT 1048.570 510.410 1048.850 514.000 ;
        RECT 1048.040 510.270 1048.850 510.410 ;
        RECT 1048.040 251.930 1048.180 510.270 ;
        RECT 1048.570 510.000 1048.850 510.270 ;
        RECT 1047.980 251.610 1048.240 251.930 ;
        RECT 1311.100 251.610 1311.360 251.930 ;
        RECT 1311.160 18.010 1311.300 251.610 ;
        RECT 1311.100 17.690 1311.360 18.010 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1317.140 2.400 1317.280 17.690 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1064.970 496.980 1065.290 497.040 ;
        RECT 1069.110 496.980 1069.430 497.040 ;
        RECT 1064.970 496.840 1069.430 496.980 ;
        RECT 1064.970 496.780 1065.290 496.840 ;
        RECT 1069.110 496.780 1069.430 496.840 ;
        RECT 1069.110 237.900 1069.430 237.960 ;
        RECT 1331.770 237.900 1332.090 237.960 ;
        RECT 1069.110 237.760 1332.090 237.900 ;
        RECT 1069.110 237.700 1069.430 237.760 ;
        RECT 1331.770 237.700 1332.090 237.760 ;
      LAYER via ;
        RECT 1065.000 496.780 1065.260 497.040 ;
        RECT 1069.140 496.780 1069.400 497.040 ;
        RECT 1069.140 237.700 1069.400 237.960 ;
        RECT 1331.800 237.700 1332.060 237.960 ;
      LAYER met2 ;
        RECT 1065.130 510.340 1065.410 514.000 ;
        RECT 1065.060 510.000 1065.410 510.340 ;
        RECT 1065.060 497.070 1065.200 510.000 ;
        RECT 1065.000 496.750 1065.260 497.070 ;
        RECT 1069.140 496.750 1069.400 497.070 ;
        RECT 1069.200 237.990 1069.340 496.750 ;
        RECT 1069.140 237.670 1069.400 237.990 ;
        RECT 1331.800 237.670 1332.060 237.990 ;
        RECT 1331.860 17.410 1332.000 237.670 ;
        RECT 1331.860 17.270 1335.220 17.410 ;
        RECT 1335.080 2.400 1335.220 17.270 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 477.090 503.440 477.410 503.500 ;
        RECT 482.150 503.440 482.470 503.500 ;
        RECT 477.090 503.300 482.470 503.440 ;
        RECT 477.090 503.240 477.410 503.300 ;
        RECT 482.150 503.240 482.470 503.300 ;
        RECT 482.150 162.080 482.470 162.140 ;
        RECT 690.070 162.080 690.390 162.140 ;
        RECT 482.150 161.940 690.390 162.080 ;
        RECT 482.150 161.880 482.470 161.940 ;
        RECT 690.070 161.880 690.390 161.940 ;
      LAYER via ;
        RECT 477.120 503.240 477.380 503.500 ;
        RECT 482.180 503.240 482.440 503.500 ;
        RECT 482.180 161.880 482.440 162.140 ;
        RECT 690.100 161.880 690.360 162.140 ;
      LAYER met2 ;
        RECT 477.250 510.340 477.530 514.000 ;
        RECT 477.180 510.000 477.530 510.340 ;
        RECT 477.180 503.530 477.320 510.000 ;
        RECT 477.120 503.210 477.380 503.530 ;
        RECT 482.180 503.210 482.440 503.530 ;
        RECT 482.240 162.170 482.380 503.210 ;
        RECT 482.180 161.850 482.440 162.170 ;
        RECT 690.100 161.850 690.360 162.170 ;
        RECT 690.160 17.410 690.300 161.850 ;
        RECT 690.160 17.270 692.600 17.410 ;
        RECT 692.460 2.400 692.600 17.270 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1082.910 128.080 1083.230 128.140 ;
        RECT 1352.930 128.080 1353.250 128.140 ;
        RECT 1082.910 127.940 1353.250 128.080 ;
        RECT 1082.910 127.880 1083.230 127.940 ;
        RECT 1352.930 127.880 1353.250 127.940 ;
      LAYER via ;
        RECT 1082.940 127.880 1083.200 128.140 ;
        RECT 1352.960 127.880 1353.220 128.140 ;
      LAYER met2 ;
        RECT 1081.230 510.410 1081.510 514.000 ;
        RECT 1081.230 510.270 1083.140 510.410 ;
        RECT 1081.230 510.000 1081.510 510.270 ;
        RECT 1083.000 128.170 1083.140 510.270 ;
        RECT 1082.940 127.850 1083.200 128.170 ;
        RECT 1352.960 127.850 1353.220 128.170 ;
        RECT 1353.020 17.410 1353.160 127.850 ;
        RECT 1352.560 17.270 1353.160 17.410 ;
        RECT 1352.560 2.400 1352.700 17.270 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1097.630 479.640 1097.950 479.700 ;
        RECT 1366.270 479.640 1366.590 479.700 ;
        RECT 1097.630 479.500 1366.590 479.640 ;
        RECT 1097.630 479.440 1097.950 479.500 ;
        RECT 1366.270 479.440 1366.590 479.500 ;
      LAYER via ;
        RECT 1097.660 479.440 1097.920 479.700 ;
        RECT 1366.300 479.440 1366.560 479.700 ;
      LAYER met2 ;
        RECT 1097.790 510.340 1098.070 514.000 ;
        RECT 1097.720 510.000 1098.070 510.340 ;
        RECT 1097.720 479.730 1097.860 510.000 ;
        RECT 1097.660 479.410 1097.920 479.730 ;
        RECT 1366.300 479.410 1366.560 479.730 ;
        RECT 1366.360 17.410 1366.500 479.410 ;
        RECT 1366.360 17.270 1370.640 17.410 ;
        RECT 1370.500 2.400 1370.640 17.270 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1117.410 134.540 1117.730 134.600 ;
        RECT 1386.970 134.540 1387.290 134.600 ;
        RECT 1117.410 134.400 1387.290 134.540 ;
        RECT 1117.410 134.340 1117.730 134.400 ;
        RECT 1386.970 134.340 1387.290 134.400 ;
      LAYER via ;
        RECT 1117.440 134.340 1117.700 134.600 ;
        RECT 1387.000 134.340 1387.260 134.600 ;
      LAYER met2 ;
        RECT 1113.890 510.410 1114.170 514.000 ;
        RECT 1113.890 510.270 1117.640 510.410 ;
        RECT 1113.890 510.000 1114.170 510.270 ;
        RECT 1117.500 134.630 1117.640 510.270 ;
        RECT 1117.440 134.310 1117.700 134.630 ;
        RECT 1387.000 134.310 1387.260 134.630 ;
        RECT 1387.060 17.410 1387.200 134.310 ;
        RECT 1387.060 17.270 1388.580 17.410 ;
        RECT 1388.440 2.400 1388.580 17.270 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1129.445 338.045 1129.615 386.155 ;
      LAYER mcon ;
        RECT 1129.445 385.985 1129.615 386.155 ;
      LAYER met1 ;
        RECT 1129.830 448.700 1130.150 448.760 ;
        RECT 1130.750 448.700 1131.070 448.760 ;
        RECT 1129.830 448.560 1131.070 448.700 ;
        RECT 1129.830 448.500 1130.150 448.560 ;
        RECT 1130.750 448.500 1131.070 448.560 ;
        RECT 1129.385 386.140 1129.675 386.185 ;
        RECT 1129.830 386.140 1130.150 386.200 ;
        RECT 1129.385 386.000 1130.150 386.140 ;
        RECT 1129.385 385.955 1129.675 386.000 ;
        RECT 1129.830 385.940 1130.150 386.000 ;
        RECT 1129.370 338.200 1129.690 338.260 ;
        RECT 1129.175 338.060 1129.690 338.200 ;
        RECT 1129.370 338.000 1129.690 338.060 ;
        RECT 1129.830 245.040 1130.150 245.100 ;
        RECT 1400.770 245.040 1401.090 245.100 ;
        RECT 1129.830 244.900 1401.090 245.040 ;
        RECT 1129.830 244.840 1130.150 244.900 ;
        RECT 1400.770 244.840 1401.090 244.900 ;
      LAYER via ;
        RECT 1129.860 448.500 1130.120 448.760 ;
        RECT 1130.780 448.500 1131.040 448.760 ;
        RECT 1129.860 385.940 1130.120 386.200 ;
        RECT 1129.400 338.000 1129.660 338.260 ;
        RECT 1129.860 244.840 1130.120 245.100 ;
        RECT 1400.800 244.840 1401.060 245.100 ;
      LAYER met2 ;
        RECT 1130.450 510.410 1130.730 514.000 ;
        RECT 1129.920 510.270 1130.730 510.410 ;
        RECT 1129.920 483.325 1130.060 510.270 ;
        RECT 1130.450 510.000 1130.730 510.270 ;
        RECT 1129.850 482.955 1130.130 483.325 ;
        RECT 1130.770 482.955 1131.050 483.325 ;
        RECT 1130.840 448.790 1130.980 482.955 ;
        RECT 1129.860 448.470 1130.120 448.790 ;
        RECT 1130.780 448.470 1131.040 448.790 ;
        RECT 1129.920 386.230 1130.060 448.470 ;
        RECT 1129.860 385.910 1130.120 386.230 ;
        RECT 1129.400 337.970 1129.660 338.290 ;
        RECT 1129.460 303.690 1129.600 337.970 ;
        RECT 1129.460 303.550 1130.520 303.690 ;
        RECT 1130.380 255.410 1130.520 303.550 ;
        RECT 1129.920 255.270 1130.520 255.410 ;
        RECT 1129.920 245.130 1130.060 255.270 ;
        RECT 1129.860 244.810 1130.120 245.130 ;
        RECT 1400.800 244.810 1401.060 245.130 ;
        RECT 1400.860 17.410 1401.000 244.810 ;
        RECT 1400.860 17.270 1406.520 17.410 ;
        RECT 1406.380 2.400 1406.520 17.270 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
      LAYER via2 ;
        RECT 1129.850 483.000 1130.130 483.280 ;
        RECT 1130.770 483.000 1131.050 483.280 ;
      LAYER met3 ;
        RECT 1129.825 483.290 1130.155 483.305 ;
        RECT 1130.745 483.290 1131.075 483.305 ;
        RECT 1129.825 482.990 1131.075 483.290 ;
        RECT 1129.825 482.975 1130.155 482.990 ;
        RECT 1130.745 482.975 1131.075 482.990 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1146.390 503.440 1146.710 503.500 ;
        RECT 1151.910 503.440 1152.230 503.500 ;
        RECT 1146.390 503.300 1152.230 503.440 ;
        RECT 1146.390 503.240 1146.710 503.300 ;
        RECT 1151.910 503.240 1152.230 503.300 ;
        RECT 1151.910 203.560 1152.230 203.620 ;
        RECT 1421.470 203.560 1421.790 203.620 ;
        RECT 1151.910 203.420 1421.790 203.560 ;
        RECT 1151.910 203.360 1152.230 203.420 ;
        RECT 1421.470 203.360 1421.790 203.420 ;
      LAYER via ;
        RECT 1146.420 503.240 1146.680 503.500 ;
        RECT 1151.940 503.240 1152.200 503.500 ;
        RECT 1151.940 203.360 1152.200 203.620 ;
        RECT 1421.500 203.360 1421.760 203.620 ;
      LAYER met2 ;
        RECT 1146.550 510.340 1146.830 514.000 ;
        RECT 1146.480 510.000 1146.830 510.340 ;
        RECT 1146.480 503.530 1146.620 510.000 ;
        RECT 1146.420 503.210 1146.680 503.530 ;
        RECT 1151.940 503.210 1152.200 503.530 ;
        RECT 1152.000 203.650 1152.140 503.210 ;
        RECT 1151.940 203.330 1152.200 203.650 ;
        RECT 1421.500 203.330 1421.760 203.650 ;
        RECT 1421.560 17.410 1421.700 203.330 ;
        RECT 1421.560 17.270 1424.000 17.410 ;
        RECT 1423.860 2.400 1424.000 17.270 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1165.710 141.340 1166.030 141.400 ;
        RECT 1435.730 141.340 1436.050 141.400 ;
        RECT 1165.710 141.200 1436.050 141.340 ;
        RECT 1165.710 141.140 1166.030 141.200 ;
        RECT 1435.730 141.140 1436.050 141.200 ;
        RECT 1435.730 17.580 1436.050 17.640 ;
        RECT 1441.710 17.580 1442.030 17.640 ;
        RECT 1435.730 17.440 1442.030 17.580 ;
        RECT 1435.730 17.380 1436.050 17.440 ;
        RECT 1441.710 17.380 1442.030 17.440 ;
      LAYER via ;
        RECT 1165.740 141.140 1166.000 141.400 ;
        RECT 1435.760 141.140 1436.020 141.400 ;
        RECT 1435.760 17.380 1436.020 17.640 ;
        RECT 1441.740 17.380 1442.000 17.640 ;
      LAYER met2 ;
        RECT 1163.110 510.410 1163.390 514.000 ;
        RECT 1163.110 510.270 1165.940 510.410 ;
        RECT 1163.110 510.000 1163.390 510.270 ;
        RECT 1165.800 141.430 1165.940 510.270 ;
        RECT 1165.740 141.110 1166.000 141.430 ;
        RECT 1435.760 141.110 1436.020 141.430 ;
        RECT 1435.820 17.670 1435.960 141.110 ;
        RECT 1435.760 17.350 1436.020 17.670 ;
        RECT 1441.740 17.350 1442.000 17.670 ;
        RECT 1441.800 2.400 1441.940 17.350 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1178.205 338.045 1178.375 386.155 ;
        RECT 1179.125 227.885 1179.295 252.195 ;
        RECT 1178.665 147.985 1178.835 207.315 ;
      LAYER mcon ;
        RECT 1178.205 385.985 1178.375 386.155 ;
        RECT 1179.125 252.025 1179.295 252.195 ;
        RECT 1178.665 207.145 1178.835 207.315 ;
      LAYER met1 ;
        RECT 1178.590 448.700 1178.910 448.760 ;
        RECT 1179.510 448.700 1179.830 448.760 ;
        RECT 1178.590 448.560 1179.830 448.700 ;
        RECT 1178.590 448.500 1178.910 448.560 ;
        RECT 1179.510 448.500 1179.830 448.560 ;
        RECT 1178.145 386.140 1178.435 386.185 ;
        RECT 1178.590 386.140 1178.910 386.200 ;
        RECT 1178.145 386.000 1178.910 386.140 ;
        RECT 1178.145 385.955 1178.435 386.000 ;
        RECT 1178.590 385.940 1178.910 386.000 ;
        RECT 1178.130 338.200 1178.450 338.260 ;
        RECT 1177.935 338.060 1178.450 338.200 ;
        RECT 1178.130 338.000 1178.450 338.060 ;
        RECT 1179.050 252.180 1179.370 252.240 ;
        RECT 1178.855 252.040 1179.370 252.180 ;
        RECT 1179.050 251.980 1179.370 252.040 ;
        RECT 1179.065 228.040 1179.355 228.085 ;
        RECT 1179.510 228.040 1179.830 228.100 ;
        RECT 1179.065 227.900 1179.830 228.040 ;
        RECT 1179.065 227.855 1179.355 227.900 ;
        RECT 1179.510 227.840 1179.830 227.900 ;
        RECT 1178.605 207.300 1178.895 207.345 ;
        RECT 1179.050 207.300 1179.370 207.360 ;
        RECT 1178.605 207.160 1179.370 207.300 ;
        RECT 1178.605 207.115 1178.895 207.160 ;
        RECT 1179.050 207.100 1179.370 207.160 ;
        RECT 1178.605 148.140 1178.895 148.185 ;
        RECT 1455.970 148.140 1456.290 148.200 ;
        RECT 1178.605 148.000 1456.290 148.140 ;
        RECT 1178.605 147.955 1178.895 148.000 ;
        RECT 1455.970 147.940 1456.290 148.000 ;
      LAYER via ;
        RECT 1178.620 448.500 1178.880 448.760 ;
        RECT 1179.540 448.500 1179.800 448.760 ;
        RECT 1178.620 385.940 1178.880 386.200 ;
        RECT 1178.160 338.000 1178.420 338.260 ;
        RECT 1179.080 251.980 1179.340 252.240 ;
        RECT 1179.540 227.840 1179.800 228.100 ;
        RECT 1179.080 207.100 1179.340 207.360 ;
        RECT 1456.000 147.940 1456.260 148.200 ;
      LAYER met2 ;
        RECT 1179.210 511.090 1179.490 514.000 ;
        RECT 1179.210 510.950 1180.200 511.090 ;
        RECT 1179.210 510.000 1179.490 510.950 ;
        RECT 1180.060 483.210 1180.200 510.950 ;
        RECT 1179.600 483.070 1180.200 483.210 ;
        RECT 1179.600 448.790 1179.740 483.070 ;
        RECT 1178.620 448.470 1178.880 448.790 ;
        RECT 1179.540 448.470 1179.800 448.790 ;
        RECT 1178.680 386.230 1178.820 448.470 ;
        RECT 1178.620 385.910 1178.880 386.230 ;
        RECT 1178.160 337.970 1178.420 338.290 ;
        RECT 1178.220 303.690 1178.360 337.970 ;
        RECT 1178.220 303.550 1179.280 303.690 ;
        RECT 1179.140 252.270 1179.280 303.550 ;
        RECT 1179.080 251.950 1179.340 252.270 ;
        RECT 1179.540 227.810 1179.800 228.130 ;
        RECT 1179.600 227.530 1179.740 227.810 ;
        RECT 1179.140 227.390 1179.740 227.530 ;
        RECT 1179.140 207.390 1179.280 227.390 ;
        RECT 1179.080 207.070 1179.340 207.390 ;
        RECT 1456.000 147.910 1456.260 148.230 ;
        RECT 1456.060 17.410 1456.200 147.910 ;
        RECT 1456.060 17.270 1459.880 17.410 ;
        RECT 1459.740 2.400 1459.880 17.270 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1195.610 498.680 1195.930 498.740 ;
        RECT 1200.210 498.680 1200.530 498.740 ;
        RECT 1195.610 498.540 1200.530 498.680 ;
        RECT 1195.610 498.480 1195.930 498.540 ;
        RECT 1200.210 498.480 1200.530 498.540 ;
        RECT 1200.210 155.280 1200.530 155.340 ;
        RECT 1476.670 155.280 1476.990 155.340 ;
        RECT 1200.210 155.140 1476.990 155.280 ;
        RECT 1200.210 155.080 1200.530 155.140 ;
        RECT 1476.670 155.080 1476.990 155.140 ;
      LAYER via ;
        RECT 1195.640 498.480 1195.900 498.740 ;
        RECT 1200.240 498.480 1200.500 498.740 ;
        RECT 1200.240 155.080 1200.500 155.340 ;
        RECT 1476.700 155.080 1476.960 155.340 ;
      LAYER met2 ;
        RECT 1195.770 510.340 1196.050 514.000 ;
        RECT 1195.700 510.000 1196.050 510.340 ;
        RECT 1195.700 498.770 1195.840 510.000 ;
        RECT 1195.640 498.450 1195.900 498.770 ;
        RECT 1200.240 498.450 1200.500 498.770 ;
        RECT 1200.300 155.370 1200.440 498.450 ;
        RECT 1200.240 155.050 1200.500 155.370 ;
        RECT 1476.700 155.050 1476.960 155.370 ;
        RECT 1476.760 17.410 1476.900 155.050 ;
        RECT 1476.760 17.270 1477.820 17.410 ;
        RECT 1477.680 2.400 1477.820 17.270 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 258.640 1214.330 258.700 ;
        RECT 1490.470 258.640 1490.790 258.700 ;
        RECT 1214.010 258.500 1490.790 258.640 ;
        RECT 1214.010 258.440 1214.330 258.500 ;
        RECT 1490.470 258.440 1490.790 258.500 ;
      LAYER via ;
        RECT 1214.040 258.440 1214.300 258.700 ;
        RECT 1490.500 258.440 1490.760 258.700 ;
      LAYER met2 ;
        RECT 1211.870 510.410 1212.150 514.000 ;
        RECT 1211.870 510.270 1214.240 510.410 ;
        RECT 1211.870 510.000 1212.150 510.270 ;
        RECT 1214.100 258.730 1214.240 510.270 ;
        RECT 1214.040 258.410 1214.300 258.730 ;
        RECT 1490.500 258.410 1490.760 258.730 ;
        RECT 1490.560 17.410 1490.700 258.410 ;
        RECT 1490.560 17.270 1495.760 17.410 ;
        RECT 1495.620 2.400 1495.760 17.270 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.350 217.160 1227.670 217.220 ;
        RECT 1511.170 217.160 1511.490 217.220 ;
        RECT 1227.350 217.020 1511.490 217.160 ;
        RECT 1227.350 216.960 1227.670 217.020 ;
        RECT 1511.170 216.960 1511.490 217.020 ;
      LAYER via ;
        RECT 1227.380 216.960 1227.640 217.220 ;
        RECT 1511.200 216.960 1511.460 217.220 ;
      LAYER met2 ;
        RECT 1227.970 510.410 1228.250 514.000 ;
        RECT 1227.440 510.270 1228.250 510.410 ;
        RECT 1227.440 217.250 1227.580 510.270 ;
        RECT 1227.970 510.000 1228.250 510.270 ;
        RECT 1227.380 216.930 1227.640 217.250 ;
        RECT 1511.200 216.930 1511.460 217.250 ;
        RECT 1511.260 17.410 1511.400 216.930 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 496.410 168.880 496.730 168.940 ;
        RECT 703.870 168.880 704.190 168.940 ;
        RECT 496.410 168.740 704.190 168.880 ;
        RECT 496.410 168.680 496.730 168.740 ;
        RECT 703.870 168.680 704.190 168.740 ;
        RECT 703.870 15.200 704.190 15.260 ;
        RECT 710.310 15.200 710.630 15.260 ;
        RECT 703.870 15.060 710.630 15.200 ;
        RECT 703.870 15.000 704.190 15.060 ;
        RECT 710.310 15.000 710.630 15.060 ;
      LAYER via ;
        RECT 496.440 168.680 496.700 168.940 ;
        RECT 703.900 168.680 704.160 168.940 ;
        RECT 703.900 15.000 704.160 15.260 ;
        RECT 710.340 15.000 710.600 15.260 ;
      LAYER met2 ;
        RECT 493.810 510.410 494.090 514.000 ;
        RECT 493.810 510.270 496.640 510.410 ;
        RECT 493.810 510.000 494.090 510.270 ;
        RECT 496.500 168.970 496.640 510.270 ;
        RECT 496.440 168.650 496.700 168.970 ;
        RECT 703.900 168.650 704.160 168.970 ;
        RECT 703.960 15.290 704.100 168.650 ;
        RECT 703.900 14.970 704.160 15.290 ;
        RECT 710.340 14.970 710.600 15.290 ;
        RECT 710.400 2.400 710.540 14.970 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1244.370 496.980 1244.690 497.040 ;
        RECT 1248.510 496.980 1248.830 497.040 ;
        RECT 1244.370 496.840 1248.830 496.980 ;
        RECT 1244.370 496.780 1244.690 496.840 ;
        RECT 1248.510 496.780 1248.830 496.840 ;
        RECT 1248.510 162.420 1248.830 162.480 ;
        RECT 1524.970 162.420 1525.290 162.480 ;
        RECT 1248.510 162.280 1525.290 162.420 ;
        RECT 1248.510 162.220 1248.830 162.280 ;
        RECT 1524.970 162.220 1525.290 162.280 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1524.970 17.440 1531.270 17.580 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
      LAYER via ;
        RECT 1244.400 496.780 1244.660 497.040 ;
        RECT 1248.540 496.780 1248.800 497.040 ;
        RECT 1248.540 162.220 1248.800 162.480 ;
        RECT 1525.000 162.220 1525.260 162.480 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
        RECT 1530.980 17.380 1531.240 17.640 ;
      LAYER met2 ;
        RECT 1244.530 510.340 1244.810 514.000 ;
        RECT 1244.460 510.000 1244.810 510.340 ;
        RECT 1244.460 497.070 1244.600 510.000 ;
        RECT 1244.400 496.750 1244.660 497.070 ;
        RECT 1248.540 496.750 1248.800 497.070 ;
        RECT 1248.600 162.510 1248.740 496.750 ;
        RECT 1248.540 162.190 1248.800 162.510 ;
        RECT 1525.000 162.190 1525.260 162.510 ;
        RECT 1525.060 17.670 1525.200 162.190 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1531.040 2.400 1531.180 17.350 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.310 120.600 1262.630 120.660 ;
        RECT 1545.670 120.600 1545.990 120.660 ;
        RECT 1262.310 120.460 1545.990 120.600 ;
        RECT 1262.310 120.400 1262.630 120.460 ;
        RECT 1545.670 120.400 1545.990 120.460 ;
      LAYER via ;
        RECT 1262.340 120.400 1262.600 120.660 ;
        RECT 1545.700 120.400 1545.960 120.660 ;
      LAYER met2 ;
        RECT 1260.630 510.410 1260.910 514.000 ;
        RECT 1260.630 510.270 1262.540 510.410 ;
        RECT 1260.630 510.000 1260.910 510.270 ;
        RECT 1262.400 120.690 1262.540 510.270 ;
        RECT 1262.340 120.370 1262.600 120.690 ;
        RECT 1545.700 120.370 1545.960 120.690 ;
        RECT 1545.760 17.410 1545.900 120.370 ;
        RECT 1545.760 17.270 1549.120 17.410 ;
        RECT 1548.980 2.400 1549.120 17.270 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.030 496.980 1277.350 497.040 ;
        RECT 1283.010 496.980 1283.330 497.040 ;
        RECT 1277.030 496.840 1283.330 496.980 ;
        RECT 1277.030 496.780 1277.350 496.840 ;
        RECT 1283.010 496.780 1283.330 496.840 ;
        RECT 1283.010 113.800 1283.330 113.860 ;
        RECT 1566.830 113.800 1567.150 113.860 ;
        RECT 1283.010 113.660 1567.150 113.800 ;
        RECT 1283.010 113.600 1283.330 113.660 ;
        RECT 1566.830 113.600 1567.150 113.660 ;
      LAYER via ;
        RECT 1277.060 496.780 1277.320 497.040 ;
        RECT 1283.040 496.780 1283.300 497.040 ;
        RECT 1283.040 113.600 1283.300 113.860 ;
        RECT 1566.860 113.600 1567.120 113.860 ;
      LAYER met2 ;
        RECT 1277.190 510.340 1277.470 514.000 ;
        RECT 1277.120 510.000 1277.470 510.340 ;
        RECT 1277.120 497.070 1277.260 510.000 ;
        RECT 1277.060 496.750 1277.320 497.070 ;
        RECT 1283.040 496.750 1283.300 497.070 ;
        RECT 1283.100 113.890 1283.240 496.750 ;
        RECT 1283.040 113.570 1283.300 113.890 ;
        RECT 1566.860 113.570 1567.120 113.890 ;
        RECT 1566.920 2.400 1567.060 113.570 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.810 176.020 1297.130 176.080 ;
        RECT 1580.170 176.020 1580.490 176.080 ;
        RECT 1296.810 175.880 1580.490 176.020 ;
        RECT 1296.810 175.820 1297.130 175.880 ;
        RECT 1580.170 175.820 1580.490 175.880 ;
      LAYER via ;
        RECT 1296.840 175.820 1297.100 176.080 ;
        RECT 1580.200 175.820 1580.460 176.080 ;
      LAYER met2 ;
        RECT 1293.290 510.410 1293.570 514.000 ;
        RECT 1293.290 510.270 1297.040 510.410 ;
        RECT 1293.290 510.000 1293.570 510.270 ;
        RECT 1296.900 176.110 1297.040 510.270 ;
        RECT 1296.840 175.790 1297.100 176.110 ;
        RECT 1580.200 175.790 1580.460 176.110 ;
        RECT 1580.260 16.730 1580.400 175.790 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 189.620 1310.930 189.680 ;
        RECT 1600.870 189.620 1601.190 189.680 ;
        RECT 1310.610 189.480 1601.190 189.620 ;
        RECT 1310.610 189.420 1310.930 189.480 ;
        RECT 1600.870 189.420 1601.190 189.480 ;
      LAYER via ;
        RECT 1310.640 189.420 1310.900 189.680 ;
        RECT 1600.900 189.420 1601.160 189.680 ;
      LAYER met2 ;
        RECT 1309.850 510.410 1310.130 514.000 ;
        RECT 1309.850 510.270 1310.840 510.410 ;
        RECT 1309.850 510.000 1310.130 510.270 ;
        RECT 1310.700 189.710 1310.840 510.270 ;
        RECT 1310.640 189.390 1310.900 189.710 ;
        RECT 1600.900 189.390 1601.160 189.710 ;
        RECT 1600.960 16.730 1601.100 189.390 ;
        RECT 1600.960 16.590 1602.480 16.730 ;
        RECT 1602.340 2.400 1602.480 16.590 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1325.790 496.980 1326.110 497.040 ;
        RECT 1330.850 496.980 1331.170 497.040 ;
        RECT 1325.790 496.840 1331.170 496.980 ;
        RECT 1325.790 496.780 1326.110 496.840 ;
        RECT 1330.850 496.780 1331.170 496.840 ;
        RECT 1330.850 127.740 1331.170 127.800 ;
        RECT 1614.670 127.740 1614.990 127.800 ;
        RECT 1330.850 127.600 1614.990 127.740 ;
        RECT 1330.850 127.540 1331.170 127.600 ;
        RECT 1614.670 127.540 1614.990 127.600 ;
      LAYER via ;
        RECT 1325.820 496.780 1326.080 497.040 ;
        RECT 1330.880 496.780 1331.140 497.040 ;
        RECT 1330.880 127.540 1331.140 127.800 ;
        RECT 1614.700 127.540 1614.960 127.800 ;
      LAYER met2 ;
        RECT 1325.950 510.340 1326.230 514.000 ;
        RECT 1325.880 510.000 1326.230 510.340 ;
        RECT 1325.880 497.070 1326.020 510.000 ;
        RECT 1325.820 496.750 1326.080 497.070 ;
        RECT 1330.880 496.750 1331.140 497.070 ;
        RECT 1330.940 127.830 1331.080 496.750 ;
        RECT 1330.880 127.510 1331.140 127.830 ;
        RECT 1614.700 127.510 1614.960 127.830 ;
        RECT 1614.760 16.730 1614.900 127.510 ;
        RECT 1614.760 16.590 1620.420 16.730 ;
        RECT 1620.280 2.400 1620.420 16.590 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 231.100 1345.430 231.160 ;
        RECT 1635.370 231.100 1635.690 231.160 ;
        RECT 1345.110 230.960 1635.690 231.100 ;
        RECT 1345.110 230.900 1345.430 230.960 ;
        RECT 1635.370 230.900 1635.690 230.960 ;
      LAYER via ;
        RECT 1345.140 230.900 1345.400 231.160 ;
        RECT 1635.400 230.900 1635.660 231.160 ;
      LAYER met2 ;
        RECT 1342.510 510.410 1342.790 514.000 ;
        RECT 1342.510 510.270 1345.340 510.410 ;
        RECT 1342.510 510.000 1342.790 510.270 ;
        RECT 1345.200 231.190 1345.340 510.270 ;
        RECT 1345.140 230.870 1345.400 231.190 ;
        RECT 1635.400 230.870 1635.660 231.190 ;
        RECT 1635.460 17.410 1635.600 230.870 ;
        RECT 1635.460 17.270 1638.360 17.410 ;
        RECT 1638.220 2.400 1638.360 17.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.450 237.900 1358.770 237.960 ;
        RECT 1656.530 237.900 1656.850 237.960 ;
        RECT 1358.450 237.760 1656.850 237.900 ;
        RECT 1358.450 237.700 1358.770 237.760 ;
        RECT 1656.530 237.700 1656.850 237.760 ;
      LAYER via ;
        RECT 1358.480 237.700 1358.740 237.960 ;
        RECT 1656.560 237.700 1656.820 237.960 ;
      LAYER met2 ;
        RECT 1358.610 510.340 1358.890 514.000 ;
        RECT 1358.540 510.000 1358.890 510.340 ;
        RECT 1358.540 237.990 1358.680 510.000 ;
        RECT 1358.480 237.670 1358.740 237.990 ;
        RECT 1656.560 237.670 1656.820 237.990 ;
        RECT 1656.620 17.410 1656.760 237.670 ;
        RECT 1656.160 17.270 1656.760 17.410 ;
        RECT 1656.160 2.400 1656.300 17.270 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.010 496.980 1375.330 497.040 ;
        RECT 1379.610 496.980 1379.930 497.040 ;
        RECT 1375.010 496.840 1379.930 496.980 ;
        RECT 1375.010 496.780 1375.330 496.840 ;
        RECT 1379.610 496.780 1379.930 496.840 ;
        RECT 1379.610 251.840 1379.930 251.900 ;
        RECT 1669.870 251.840 1670.190 251.900 ;
        RECT 1379.610 251.700 1670.190 251.840 ;
        RECT 1379.610 251.640 1379.930 251.700 ;
        RECT 1669.870 251.640 1670.190 251.700 ;
      LAYER via ;
        RECT 1375.040 496.780 1375.300 497.040 ;
        RECT 1379.640 496.780 1379.900 497.040 ;
        RECT 1379.640 251.640 1379.900 251.900 ;
        RECT 1669.900 251.640 1670.160 251.900 ;
      LAYER met2 ;
        RECT 1375.170 510.340 1375.450 514.000 ;
        RECT 1375.100 510.000 1375.450 510.340 ;
        RECT 1375.100 497.070 1375.240 510.000 ;
        RECT 1375.040 496.750 1375.300 497.070 ;
        RECT 1379.640 496.750 1379.900 497.070 ;
        RECT 1379.700 251.930 1379.840 496.750 ;
        RECT 1379.640 251.610 1379.900 251.930 ;
        RECT 1669.900 251.610 1670.160 251.930 ;
        RECT 1669.960 17.410 1670.100 251.610 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.410 134.540 1393.730 134.600 ;
        RECT 1690.570 134.540 1690.890 134.600 ;
        RECT 1393.410 134.400 1690.890 134.540 ;
        RECT 1393.410 134.340 1393.730 134.400 ;
        RECT 1690.570 134.340 1690.890 134.400 ;
      LAYER via ;
        RECT 1393.440 134.340 1393.700 134.600 ;
        RECT 1690.600 134.340 1690.860 134.600 ;
      LAYER met2 ;
        RECT 1391.270 510.410 1391.550 514.000 ;
        RECT 1391.270 510.270 1393.640 510.410 ;
        RECT 1391.270 510.000 1391.550 510.270 ;
        RECT 1393.500 134.630 1393.640 510.270 ;
        RECT 1393.440 134.310 1393.700 134.630 ;
        RECT 1690.600 134.310 1690.860 134.630 ;
        RECT 1690.660 17.410 1690.800 134.310 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.210 176.020 510.530 176.080 ;
        RECT 724.570 176.020 724.890 176.080 ;
        RECT 510.210 175.880 724.890 176.020 ;
        RECT 510.210 175.820 510.530 175.880 ;
        RECT 724.570 175.820 724.890 175.880 ;
      LAYER via ;
        RECT 510.240 175.820 510.500 176.080 ;
        RECT 724.600 175.820 724.860 176.080 ;
      LAYER met2 ;
        RECT 509.910 511.090 510.190 514.000 ;
        RECT 509.910 510.950 510.900 511.090 ;
        RECT 509.910 510.000 510.190 510.950 ;
        RECT 510.760 496.810 510.900 510.950 ;
        RECT 510.300 496.670 510.900 496.810 ;
        RECT 510.300 176.110 510.440 496.670 ;
        RECT 510.240 175.790 510.500 176.110 ;
        RECT 724.600 175.790 724.860 176.110 ;
        RECT 724.660 17.410 724.800 175.790 ;
        RECT 724.660 17.270 728.480 17.410 ;
        RECT 728.340 2.400 728.480 17.270 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.670 479.640 1407.990 479.700 ;
        RECT 1704.370 479.640 1704.690 479.700 ;
        RECT 1407.670 479.500 1704.690 479.640 ;
        RECT 1407.670 479.440 1407.990 479.500 ;
        RECT 1704.370 479.440 1704.690 479.500 ;
      LAYER via ;
        RECT 1407.700 479.440 1407.960 479.700 ;
        RECT 1704.400 479.440 1704.660 479.700 ;
      LAYER met2 ;
        RECT 1407.830 510.340 1408.110 514.000 ;
        RECT 1407.760 510.000 1408.110 510.340 ;
        RECT 1407.760 479.730 1407.900 510.000 ;
        RECT 1407.700 479.410 1407.960 479.730 ;
        RECT 1704.400 479.410 1704.660 479.730 ;
        RECT 1704.460 17.410 1704.600 479.410 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.770 496.980 1424.090 497.040 ;
        RECT 1427.910 496.980 1428.230 497.040 ;
        RECT 1423.770 496.840 1428.230 496.980 ;
        RECT 1423.770 496.780 1424.090 496.840 ;
        RECT 1427.910 496.780 1428.230 496.840 ;
        RECT 1427.910 203.560 1428.230 203.620 ;
        RECT 1725.070 203.560 1725.390 203.620 ;
        RECT 1427.910 203.420 1725.390 203.560 ;
        RECT 1427.910 203.360 1428.230 203.420 ;
        RECT 1725.070 203.360 1725.390 203.420 ;
      LAYER via ;
        RECT 1423.800 496.780 1424.060 497.040 ;
        RECT 1427.940 496.780 1428.200 497.040 ;
        RECT 1427.940 203.360 1428.200 203.620 ;
        RECT 1725.100 203.360 1725.360 203.620 ;
      LAYER met2 ;
        RECT 1423.930 510.340 1424.210 514.000 ;
        RECT 1423.860 510.000 1424.210 510.340 ;
        RECT 1423.860 497.070 1424.000 510.000 ;
        RECT 1423.800 496.750 1424.060 497.070 ;
        RECT 1427.940 496.750 1428.200 497.070 ;
        RECT 1428.000 203.650 1428.140 496.750 ;
        RECT 1427.940 203.330 1428.200 203.650 ;
        RECT 1725.100 203.330 1725.360 203.650 ;
        RECT 1725.160 17.410 1725.300 203.330 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 141.340 1442.030 141.400 ;
        RECT 1738.870 141.340 1739.190 141.400 ;
        RECT 1441.710 141.200 1739.190 141.340 ;
        RECT 1441.710 141.140 1442.030 141.200 ;
        RECT 1738.870 141.140 1739.190 141.200 ;
        RECT 1738.870 17.580 1739.190 17.640 ;
        RECT 1745.310 17.580 1745.630 17.640 ;
        RECT 1738.870 17.440 1745.630 17.580 ;
        RECT 1738.870 17.380 1739.190 17.440 ;
        RECT 1745.310 17.380 1745.630 17.440 ;
      LAYER via ;
        RECT 1441.740 141.140 1442.000 141.400 ;
        RECT 1738.900 141.140 1739.160 141.400 ;
        RECT 1738.900 17.380 1739.160 17.640 ;
        RECT 1745.340 17.380 1745.600 17.640 ;
      LAYER met2 ;
        RECT 1440.490 510.410 1440.770 514.000 ;
        RECT 1440.490 510.270 1441.940 510.410 ;
        RECT 1440.490 510.000 1440.770 510.270 ;
        RECT 1441.800 141.430 1441.940 510.270 ;
        RECT 1441.740 141.110 1442.000 141.430 ;
        RECT 1738.900 141.110 1739.160 141.430 ;
        RECT 1738.960 17.670 1739.100 141.110 ;
        RECT 1738.900 17.350 1739.160 17.670 ;
        RECT 1745.340 17.350 1745.600 17.670 ;
        RECT 1745.400 2.400 1745.540 17.350 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1456.430 496.980 1456.750 497.040 ;
        RECT 1462.410 496.980 1462.730 497.040 ;
        RECT 1456.430 496.840 1462.730 496.980 ;
        RECT 1456.430 496.780 1456.750 496.840 ;
        RECT 1462.410 496.780 1462.730 496.840 ;
        RECT 1462.410 245.040 1462.730 245.100 ;
        RECT 1759.570 245.040 1759.890 245.100 ;
        RECT 1462.410 244.900 1759.890 245.040 ;
        RECT 1462.410 244.840 1462.730 244.900 ;
        RECT 1759.570 244.840 1759.890 244.900 ;
        RECT 1759.570 62.120 1759.890 62.180 ;
        RECT 1762.790 62.120 1763.110 62.180 ;
        RECT 1759.570 61.980 1763.110 62.120 ;
        RECT 1759.570 61.920 1759.890 61.980 ;
        RECT 1762.790 61.920 1763.110 61.980 ;
      LAYER via ;
        RECT 1456.460 496.780 1456.720 497.040 ;
        RECT 1462.440 496.780 1462.700 497.040 ;
        RECT 1462.440 244.840 1462.700 245.100 ;
        RECT 1759.600 244.840 1759.860 245.100 ;
        RECT 1759.600 61.920 1759.860 62.180 ;
        RECT 1762.820 61.920 1763.080 62.180 ;
      LAYER met2 ;
        RECT 1456.590 510.340 1456.870 514.000 ;
        RECT 1456.520 510.000 1456.870 510.340 ;
        RECT 1456.520 497.070 1456.660 510.000 ;
        RECT 1456.460 496.750 1456.720 497.070 ;
        RECT 1462.440 496.750 1462.700 497.070 ;
        RECT 1462.500 245.130 1462.640 496.750 ;
        RECT 1462.440 244.810 1462.700 245.130 ;
        RECT 1759.600 244.810 1759.860 245.130 ;
        RECT 1759.660 62.210 1759.800 244.810 ;
        RECT 1759.600 61.890 1759.860 62.210 ;
        RECT 1762.820 61.890 1763.080 62.210 ;
        RECT 1762.880 2.400 1763.020 61.890 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1476.210 210.360 1476.530 210.420 ;
        RECT 1780.730 210.360 1781.050 210.420 ;
        RECT 1476.210 210.220 1781.050 210.360 ;
        RECT 1476.210 210.160 1476.530 210.220 ;
        RECT 1780.730 210.160 1781.050 210.220 ;
      LAYER via ;
        RECT 1476.240 210.160 1476.500 210.420 ;
        RECT 1780.760 210.160 1781.020 210.420 ;
      LAYER met2 ;
        RECT 1473.150 510.410 1473.430 514.000 ;
        RECT 1473.150 510.270 1476.440 510.410 ;
        RECT 1473.150 510.000 1473.430 510.270 ;
        RECT 1476.300 210.450 1476.440 510.270 ;
        RECT 1476.240 210.130 1476.500 210.450 ;
        RECT 1780.760 210.130 1781.020 210.450 ;
        RECT 1780.820 2.400 1780.960 210.130 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1488.705 338.045 1488.875 386.155 ;
      LAYER mcon ;
        RECT 1488.705 385.985 1488.875 386.155 ;
      LAYER met1 ;
        RECT 1488.630 448.700 1488.950 448.760 ;
        RECT 1489.550 448.700 1489.870 448.760 ;
        RECT 1488.630 448.560 1489.870 448.700 ;
        RECT 1488.630 448.500 1488.950 448.560 ;
        RECT 1489.550 448.500 1489.870 448.560 ;
        RECT 1488.630 386.140 1488.950 386.200 ;
        RECT 1488.435 386.000 1488.950 386.140 ;
        RECT 1488.630 385.940 1488.950 386.000 ;
        RECT 1488.645 338.200 1488.935 338.245 ;
        RECT 1489.090 338.200 1489.410 338.260 ;
        RECT 1488.645 338.060 1489.410 338.200 ;
        RECT 1488.645 338.015 1488.935 338.060 ;
        RECT 1489.090 338.000 1489.410 338.060 ;
        RECT 1489.090 304.200 1489.410 304.260 ;
        RECT 1488.720 304.060 1489.410 304.200 ;
        RECT 1488.720 303.580 1488.860 304.060 ;
        RECT 1489.090 304.000 1489.410 304.060 ;
        RECT 1488.630 303.320 1488.950 303.580 ;
        RECT 1488.630 265.440 1488.950 265.500 ;
        RECT 1794.070 265.440 1794.390 265.500 ;
        RECT 1488.630 265.300 1794.390 265.440 ;
        RECT 1488.630 265.240 1488.950 265.300 ;
        RECT 1794.070 265.240 1794.390 265.300 ;
        RECT 1794.070 62.120 1794.390 62.180 ;
        RECT 1798.670 62.120 1798.990 62.180 ;
        RECT 1794.070 61.980 1798.990 62.120 ;
        RECT 1794.070 61.920 1794.390 61.980 ;
        RECT 1798.670 61.920 1798.990 61.980 ;
      LAYER via ;
        RECT 1488.660 448.500 1488.920 448.760 ;
        RECT 1489.580 448.500 1489.840 448.760 ;
        RECT 1488.660 385.940 1488.920 386.200 ;
        RECT 1489.120 338.000 1489.380 338.260 ;
        RECT 1489.120 304.000 1489.380 304.260 ;
        RECT 1488.660 303.320 1488.920 303.580 ;
        RECT 1488.660 265.240 1488.920 265.500 ;
        RECT 1794.100 265.240 1794.360 265.500 ;
        RECT 1794.100 61.920 1794.360 62.180 ;
        RECT 1798.700 61.920 1798.960 62.180 ;
      LAYER met2 ;
        RECT 1489.250 510.410 1489.530 514.000 ;
        RECT 1488.720 510.270 1489.530 510.410 ;
        RECT 1488.720 483.325 1488.860 510.270 ;
        RECT 1489.250 510.000 1489.530 510.270 ;
        RECT 1488.650 482.955 1488.930 483.325 ;
        RECT 1489.570 482.955 1489.850 483.325 ;
        RECT 1489.640 448.790 1489.780 482.955 ;
        RECT 1488.660 448.470 1488.920 448.790 ;
        RECT 1489.580 448.470 1489.840 448.790 ;
        RECT 1488.720 386.230 1488.860 448.470 ;
        RECT 1488.660 385.910 1488.920 386.230 ;
        RECT 1489.120 337.970 1489.380 338.290 ;
        RECT 1489.180 304.290 1489.320 337.970 ;
        RECT 1489.120 303.970 1489.380 304.290 ;
        RECT 1488.660 303.290 1488.920 303.610 ;
        RECT 1488.720 265.530 1488.860 303.290 ;
        RECT 1488.660 265.210 1488.920 265.530 ;
        RECT 1794.100 265.210 1794.360 265.530 ;
        RECT 1794.160 62.210 1794.300 265.210 ;
        RECT 1794.100 61.890 1794.360 62.210 ;
        RECT 1798.700 61.890 1798.960 62.210 ;
        RECT 1798.760 2.400 1798.900 61.890 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 1488.650 483.000 1488.930 483.280 ;
        RECT 1489.570 483.000 1489.850 483.280 ;
      LAYER met3 ;
        RECT 1488.625 483.290 1488.955 483.305 ;
        RECT 1489.545 483.290 1489.875 483.305 ;
        RECT 1488.625 482.990 1489.875 483.290 ;
        RECT 1488.625 482.975 1488.955 482.990 ;
        RECT 1489.545 482.975 1489.875 482.990 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1505.650 501.060 1505.970 501.120 ;
        RECT 1510.710 501.060 1511.030 501.120 ;
        RECT 1505.650 500.920 1511.030 501.060 ;
        RECT 1505.650 500.860 1505.970 500.920 ;
        RECT 1510.710 500.860 1511.030 500.920 ;
        RECT 1510.710 162.080 1511.030 162.140 ;
        RECT 1814.770 162.080 1815.090 162.140 ;
        RECT 1510.710 161.940 1815.090 162.080 ;
        RECT 1510.710 161.880 1511.030 161.940 ;
        RECT 1814.770 161.880 1815.090 161.940 ;
      LAYER via ;
        RECT 1505.680 500.860 1505.940 501.120 ;
        RECT 1510.740 500.860 1511.000 501.120 ;
        RECT 1510.740 161.880 1511.000 162.140 ;
        RECT 1814.800 161.880 1815.060 162.140 ;
      LAYER met2 ;
        RECT 1505.810 510.340 1506.090 514.000 ;
        RECT 1505.740 510.000 1506.090 510.340 ;
        RECT 1505.740 501.150 1505.880 510.000 ;
        RECT 1505.680 500.830 1505.940 501.150 ;
        RECT 1510.740 500.830 1511.000 501.150 ;
        RECT 1510.800 162.170 1510.940 500.830 ;
        RECT 1510.740 161.850 1511.000 162.170 ;
        RECT 1814.800 161.850 1815.060 162.170 ;
        RECT 1814.860 17.410 1815.000 161.850 ;
        RECT 1814.860 17.270 1816.840 17.410 ;
        RECT 1816.700 2.400 1816.840 17.270 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.510 217.160 1524.830 217.220 ;
        RECT 1828.570 217.160 1828.890 217.220 ;
        RECT 1524.510 217.020 1828.890 217.160 ;
        RECT 1524.510 216.960 1524.830 217.020 ;
        RECT 1828.570 216.960 1828.890 217.020 ;
        RECT 1828.570 17.920 1828.890 17.980 ;
        RECT 1834.550 17.920 1834.870 17.980 ;
        RECT 1828.570 17.780 1834.870 17.920 ;
        RECT 1828.570 17.720 1828.890 17.780 ;
        RECT 1834.550 17.720 1834.870 17.780 ;
      LAYER via ;
        RECT 1524.540 216.960 1524.800 217.220 ;
        RECT 1828.600 216.960 1828.860 217.220 ;
        RECT 1828.600 17.720 1828.860 17.980 ;
        RECT 1834.580 17.720 1834.840 17.980 ;
      LAYER met2 ;
        RECT 1521.910 510.410 1522.190 514.000 ;
        RECT 1521.910 510.270 1524.740 510.410 ;
        RECT 1521.910 510.000 1522.190 510.270 ;
        RECT 1524.600 217.250 1524.740 510.270 ;
        RECT 1524.540 216.930 1524.800 217.250 ;
        RECT 1828.600 216.930 1828.860 217.250 ;
        RECT 1828.660 18.010 1828.800 216.930 ;
        RECT 1828.600 17.690 1828.860 18.010 ;
        RECT 1834.580 17.690 1834.840 18.010 ;
        RECT 1834.640 2.400 1834.780 17.690 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1849.345 48.365 1849.515 96.475 ;
      LAYER mcon ;
        RECT 1849.345 96.305 1849.515 96.475 ;
      LAYER met1 ;
        RECT 1538.310 279.380 1538.630 279.440 ;
        RECT 1849.270 279.380 1849.590 279.440 ;
        RECT 1538.310 279.240 1849.590 279.380 ;
        RECT 1538.310 279.180 1538.630 279.240 ;
        RECT 1849.270 279.180 1849.590 279.240 ;
        RECT 1849.270 96.460 1849.590 96.520 ;
        RECT 1849.075 96.320 1849.590 96.460 ;
        RECT 1849.270 96.260 1849.590 96.320 ;
        RECT 1849.285 48.520 1849.575 48.565 ;
        RECT 1852.030 48.520 1852.350 48.580 ;
        RECT 1849.285 48.380 1852.350 48.520 ;
        RECT 1849.285 48.335 1849.575 48.380 ;
        RECT 1852.030 48.320 1852.350 48.380 ;
      LAYER via ;
        RECT 1538.340 279.180 1538.600 279.440 ;
        RECT 1849.300 279.180 1849.560 279.440 ;
        RECT 1849.300 96.260 1849.560 96.520 ;
        RECT 1852.060 48.320 1852.320 48.580 ;
      LAYER met2 ;
        RECT 1538.470 510.340 1538.750 514.000 ;
        RECT 1538.400 510.000 1538.750 510.340 ;
        RECT 1538.400 279.470 1538.540 510.000 ;
        RECT 1538.340 279.150 1538.600 279.470 ;
        RECT 1849.300 279.150 1849.560 279.470 ;
        RECT 1849.360 96.550 1849.500 279.150 ;
        RECT 1849.300 96.230 1849.560 96.550 ;
        RECT 1852.060 48.290 1852.320 48.610 ;
        RECT 1852.120 2.400 1852.260 48.290 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1554.410 496.980 1554.730 497.040 ;
        RECT 1559.010 496.980 1559.330 497.040 ;
        RECT 1554.410 496.840 1559.330 496.980 ;
        RECT 1554.410 496.780 1554.730 496.840 ;
        RECT 1559.010 496.780 1559.330 496.840 ;
        RECT 1559.010 182.820 1559.330 182.880 ;
        RECT 1870.430 182.820 1870.750 182.880 ;
        RECT 1559.010 182.680 1870.750 182.820 ;
        RECT 1559.010 182.620 1559.330 182.680 ;
        RECT 1870.430 182.620 1870.750 182.680 ;
      LAYER via ;
        RECT 1554.440 496.780 1554.700 497.040 ;
        RECT 1559.040 496.780 1559.300 497.040 ;
        RECT 1559.040 182.620 1559.300 182.880 ;
        RECT 1870.460 182.620 1870.720 182.880 ;
      LAYER met2 ;
        RECT 1554.570 510.340 1554.850 514.000 ;
        RECT 1554.500 510.000 1554.850 510.340 ;
        RECT 1554.500 497.070 1554.640 510.000 ;
        RECT 1554.440 496.750 1554.700 497.070 ;
        RECT 1559.040 496.750 1559.300 497.070 ;
        RECT 1559.100 182.910 1559.240 496.750 ;
        RECT 1559.040 182.590 1559.300 182.910 ;
        RECT 1870.460 182.590 1870.720 182.910 ;
        RECT 1870.520 7.210 1870.660 182.590 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 526.310 503.440 526.630 503.500 ;
        RECT 530.910 503.440 531.230 503.500 ;
        RECT 526.310 503.300 531.230 503.440 ;
        RECT 526.310 503.240 526.630 503.300 ;
        RECT 530.910 503.240 531.230 503.300 ;
        RECT 530.910 182.820 531.230 182.880 ;
        RECT 745.270 182.820 745.590 182.880 ;
        RECT 530.910 182.680 745.590 182.820 ;
        RECT 530.910 182.620 531.230 182.680 ;
        RECT 745.270 182.620 745.590 182.680 ;
      LAYER via ;
        RECT 526.340 503.240 526.600 503.500 ;
        RECT 530.940 503.240 531.200 503.500 ;
        RECT 530.940 182.620 531.200 182.880 ;
        RECT 745.300 182.620 745.560 182.880 ;
      LAYER met2 ;
        RECT 526.470 510.340 526.750 514.000 ;
        RECT 526.400 510.000 526.750 510.340 ;
        RECT 526.400 503.530 526.540 510.000 ;
        RECT 526.340 503.210 526.600 503.530 ;
        RECT 530.940 503.210 531.200 503.530 ;
        RECT 531.000 182.910 531.140 503.210 ;
        RECT 530.940 182.590 531.200 182.910 ;
        RECT 745.300 182.590 745.560 182.910 ;
        RECT 745.360 17.410 745.500 182.590 ;
        RECT 745.360 17.270 746.420 17.410 ;
        RECT 746.280 2.400 746.420 17.270 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.810 293.320 1573.130 293.380 ;
        RECT 1883.770 293.320 1884.090 293.380 ;
        RECT 1572.810 293.180 1884.090 293.320 ;
        RECT 1572.810 293.120 1573.130 293.180 ;
        RECT 1883.770 293.120 1884.090 293.180 ;
        RECT 1883.770 62.120 1884.090 62.180 ;
        RECT 1887.910 62.120 1888.230 62.180 ;
        RECT 1883.770 61.980 1888.230 62.120 ;
        RECT 1883.770 61.920 1884.090 61.980 ;
        RECT 1887.910 61.920 1888.230 61.980 ;
      LAYER via ;
        RECT 1572.840 293.120 1573.100 293.380 ;
        RECT 1883.800 293.120 1884.060 293.380 ;
        RECT 1883.800 61.920 1884.060 62.180 ;
        RECT 1887.940 61.920 1888.200 62.180 ;
      LAYER met2 ;
        RECT 1571.130 510.410 1571.410 514.000 ;
        RECT 1571.130 510.270 1573.040 510.410 ;
        RECT 1571.130 510.000 1571.410 510.270 ;
        RECT 1572.900 293.410 1573.040 510.270 ;
        RECT 1572.840 293.090 1573.100 293.410 ;
        RECT 1883.800 293.090 1884.060 293.410 ;
        RECT 1883.860 62.210 1884.000 293.090 ;
        RECT 1883.800 61.890 1884.060 62.210 ;
        RECT 1887.940 61.890 1888.200 62.210 ;
        RECT 1888.000 2.400 1888.140 61.890 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1587.070 486.440 1587.390 486.500 ;
        RECT 1904.470 486.440 1904.790 486.500 ;
        RECT 1587.070 486.300 1904.790 486.440 ;
        RECT 1587.070 486.240 1587.390 486.300 ;
        RECT 1904.470 486.240 1904.790 486.300 ;
      LAYER via ;
        RECT 1587.100 486.240 1587.360 486.500 ;
        RECT 1904.500 486.240 1904.760 486.500 ;
      LAYER met2 ;
        RECT 1587.230 510.340 1587.510 514.000 ;
        RECT 1587.160 510.000 1587.510 510.340 ;
        RECT 1587.160 486.530 1587.300 510.000 ;
        RECT 1587.100 486.210 1587.360 486.530 ;
        RECT 1904.500 486.210 1904.760 486.530 ;
        RECT 1904.560 16.730 1904.700 486.210 ;
        RECT 1904.560 16.590 1906.080 16.730 ;
        RECT 1905.940 2.400 1906.080 16.590 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1603.170 496.980 1603.490 497.040 ;
        RECT 1607.310 496.980 1607.630 497.040 ;
        RECT 1603.170 496.840 1607.630 496.980 ;
        RECT 1603.170 496.780 1603.490 496.840 ;
        RECT 1607.310 496.780 1607.630 496.840 ;
        RECT 1607.310 176.020 1607.630 176.080 ;
        RECT 1918.270 176.020 1918.590 176.080 ;
        RECT 1607.310 175.880 1918.590 176.020 ;
        RECT 1607.310 175.820 1607.630 175.880 ;
        RECT 1918.270 175.820 1918.590 175.880 ;
      LAYER via ;
        RECT 1603.200 496.780 1603.460 497.040 ;
        RECT 1607.340 496.780 1607.600 497.040 ;
        RECT 1607.340 175.820 1607.600 176.080 ;
        RECT 1918.300 175.820 1918.560 176.080 ;
      LAYER met2 ;
        RECT 1603.330 510.340 1603.610 514.000 ;
        RECT 1603.260 510.000 1603.610 510.340 ;
        RECT 1603.260 497.070 1603.400 510.000 ;
        RECT 1603.200 496.750 1603.460 497.070 ;
        RECT 1607.340 496.750 1607.600 497.070 ;
        RECT 1607.400 176.110 1607.540 496.750 ;
        RECT 1607.340 175.790 1607.600 176.110 ;
        RECT 1918.300 175.790 1918.560 176.110 ;
        RECT 1918.360 16.730 1918.500 175.790 ;
        RECT 1918.360 16.590 1923.560 16.730 ;
        RECT 1923.420 2.400 1923.560 16.590 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1621.110 224.300 1621.430 224.360 ;
        RECT 1938.970 224.300 1939.290 224.360 ;
        RECT 1621.110 224.160 1939.290 224.300 ;
        RECT 1621.110 224.100 1621.430 224.160 ;
        RECT 1938.970 224.100 1939.290 224.160 ;
      LAYER via ;
        RECT 1621.140 224.100 1621.400 224.360 ;
        RECT 1939.000 224.100 1939.260 224.360 ;
      LAYER met2 ;
        RECT 1619.890 510.410 1620.170 514.000 ;
        RECT 1619.890 510.270 1621.340 510.410 ;
        RECT 1619.890 510.000 1620.170 510.270 ;
        RECT 1621.200 224.390 1621.340 510.270 ;
        RECT 1621.140 224.070 1621.400 224.390 ;
        RECT 1939.000 224.070 1939.260 224.390 ;
        RECT 1939.060 16.730 1939.200 224.070 ;
        RECT 1939.060 16.590 1941.500 16.730 ;
        RECT 1941.360 2.400 1941.500 16.590 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1635.830 503.440 1636.150 503.500 ;
        RECT 1645.490 503.440 1645.810 503.500 ;
        RECT 1635.830 503.300 1645.810 503.440 ;
        RECT 1635.830 503.240 1636.150 503.300 ;
        RECT 1645.490 503.240 1645.810 503.300 ;
        RECT 1645.490 231.100 1645.810 231.160 ;
        RECT 1952.770 231.100 1953.090 231.160 ;
        RECT 1645.490 230.960 1953.090 231.100 ;
        RECT 1645.490 230.900 1645.810 230.960 ;
        RECT 1952.770 230.900 1953.090 230.960 ;
        RECT 1952.770 37.980 1953.090 38.040 ;
        RECT 1959.210 37.980 1959.530 38.040 ;
        RECT 1952.770 37.840 1959.530 37.980 ;
        RECT 1952.770 37.780 1953.090 37.840 ;
        RECT 1959.210 37.780 1959.530 37.840 ;
      LAYER via ;
        RECT 1635.860 503.240 1636.120 503.500 ;
        RECT 1645.520 503.240 1645.780 503.500 ;
        RECT 1645.520 230.900 1645.780 231.160 ;
        RECT 1952.800 230.900 1953.060 231.160 ;
        RECT 1952.800 37.780 1953.060 38.040 ;
        RECT 1959.240 37.780 1959.500 38.040 ;
      LAYER met2 ;
        RECT 1635.990 510.340 1636.270 514.000 ;
        RECT 1635.920 510.000 1636.270 510.340 ;
        RECT 1635.920 503.530 1636.060 510.000 ;
        RECT 1635.860 503.210 1636.120 503.530 ;
        RECT 1645.520 503.210 1645.780 503.530 ;
        RECT 1645.580 231.190 1645.720 503.210 ;
        RECT 1645.520 230.870 1645.780 231.190 ;
        RECT 1952.800 230.870 1953.060 231.190 ;
        RECT 1952.860 38.070 1953.000 230.870 ;
        RECT 1952.800 37.750 1953.060 38.070 ;
        RECT 1959.240 37.750 1959.500 38.070 ;
        RECT 1959.300 2.400 1959.440 37.750 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 189.620 1655.930 189.680 ;
        RECT 1973.470 189.620 1973.790 189.680 ;
        RECT 1655.610 189.480 1973.790 189.620 ;
        RECT 1655.610 189.420 1655.930 189.480 ;
        RECT 1973.470 189.420 1973.790 189.480 ;
        RECT 1973.470 62.260 1973.790 62.520 ;
        RECT 1973.560 61.780 1973.700 62.260 ;
        RECT 1977.150 61.780 1977.470 61.840 ;
        RECT 1973.560 61.640 1977.470 61.780 ;
        RECT 1977.150 61.580 1977.470 61.640 ;
        RECT 1977.150 47.980 1977.470 48.240 ;
        RECT 1977.240 47.560 1977.380 47.980 ;
        RECT 1977.150 47.300 1977.470 47.560 ;
      LAYER via ;
        RECT 1655.640 189.420 1655.900 189.680 ;
        RECT 1973.500 189.420 1973.760 189.680 ;
        RECT 1973.500 62.260 1973.760 62.520 ;
        RECT 1977.180 61.580 1977.440 61.840 ;
        RECT 1977.180 47.980 1977.440 48.240 ;
        RECT 1977.180 47.300 1977.440 47.560 ;
      LAYER met2 ;
        RECT 1652.550 510.410 1652.830 514.000 ;
        RECT 1652.550 510.270 1655.840 510.410 ;
        RECT 1652.550 510.000 1652.830 510.270 ;
        RECT 1655.700 189.710 1655.840 510.270 ;
        RECT 1655.640 189.390 1655.900 189.710 ;
        RECT 1973.500 189.390 1973.760 189.710 ;
        RECT 1973.560 62.550 1973.700 189.390 ;
        RECT 1973.500 62.230 1973.760 62.550 ;
        RECT 1977.180 61.550 1977.440 61.870 ;
        RECT 1977.240 48.270 1977.380 61.550 ;
        RECT 1977.180 47.950 1977.440 48.270 ;
        RECT 1977.180 47.270 1977.440 47.590 ;
        RECT 1977.240 2.400 1977.380 47.270 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1669.025 237.745 1669.195 240.975 ;
      LAYER mcon ;
        RECT 1669.025 240.805 1669.195 240.975 ;
      LAYER met1 ;
        RECT 1668.490 289.920 1668.810 289.980 ;
        RECT 1668.950 289.920 1669.270 289.980 ;
        RECT 1668.490 289.780 1669.270 289.920 ;
        RECT 1668.490 289.720 1668.810 289.780 ;
        RECT 1668.950 289.720 1669.270 289.780 ;
        RECT 1668.950 240.960 1669.270 241.020 ;
        RECT 1668.755 240.820 1669.270 240.960 ;
        RECT 1668.950 240.760 1669.270 240.820 ;
        RECT 1668.965 237.900 1669.255 237.945 ;
        RECT 1994.170 237.900 1994.490 237.960 ;
        RECT 1668.965 237.760 1994.490 237.900 ;
        RECT 1668.965 237.715 1669.255 237.760 ;
        RECT 1994.170 237.700 1994.490 237.760 ;
      LAYER via ;
        RECT 1668.520 289.720 1668.780 289.980 ;
        RECT 1668.980 289.720 1669.240 289.980 ;
        RECT 1668.980 240.760 1669.240 241.020 ;
        RECT 1994.200 237.700 1994.460 237.960 ;
      LAYER met2 ;
        RECT 1668.650 510.410 1668.930 514.000 ;
        RECT 1668.120 510.270 1668.930 510.410 ;
        RECT 1668.120 483.325 1668.260 510.270 ;
        RECT 1668.650 510.000 1668.930 510.270 ;
        RECT 1668.050 482.955 1668.330 483.325 ;
        RECT 1668.970 482.955 1669.250 483.325 ;
        RECT 1669.040 337.690 1669.180 482.955 ;
        RECT 1668.580 337.550 1669.180 337.690 ;
        RECT 1668.580 290.010 1668.720 337.550 ;
        RECT 1668.520 289.690 1668.780 290.010 ;
        RECT 1668.980 289.690 1669.240 290.010 ;
        RECT 1669.040 241.050 1669.180 289.690 ;
        RECT 1668.980 240.730 1669.240 241.050 ;
        RECT 1994.200 237.670 1994.460 237.990 ;
        RECT 1994.260 16.730 1994.400 237.670 ;
        RECT 1994.260 16.590 1995.320 16.730 ;
        RECT 1995.180 2.400 1995.320 16.590 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
      LAYER via2 ;
        RECT 1668.050 483.000 1668.330 483.280 ;
        RECT 1668.970 483.000 1669.250 483.280 ;
      LAYER met3 ;
        RECT 1668.025 483.290 1668.355 483.305 ;
        RECT 1668.945 483.290 1669.275 483.305 ;
        RECT 1668.025 482.990 1669.275 483.290 ;
        RECT 1668.025 482.975 1668.355 482.990 ;
        RECT 1668.945 482.975 1669.275 482.990 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1685.050 503.440 1685.370 503.500 ;
        RECT 1690.110 503.440 1690.430 503.500 ;
        RECT 1685.050 503.300 1690.430 503.440 ;
        RECT 1685.050 503.240 1685.370 503.300 ;
        RECT 1690.110 503.240 1690.430 503.300 ;
        RECT 1690.110 251.840 1690.430 251.900 ;
        RECT 2007.970 251.840 2008.290 251.900 ;
        RECT 1690.110 251.700 2008.290 251.840 ;
        RECT 1690.110 251.640 1690.430 251.700 ;
        RECT 2007.970 251.640 2008.290 251.700 ;
      LAYER via ;
        RECT 1685.080 503.240 1685.340 503.500 ;
        RECT 1690.140 503.240 1690.400 503.500 ;
        RECT 1690.140 251.640 1690.400 251.900 ;
        RECT 2008.000 251.640 2008.260 251.900 ;
      LAYER met2 ;
        RECT 1685.210 510.340 1685.490 514.000 ;
        RECT 1685.140 510.000 1685.490 510.340 ;
        RECT 1685.140 503.530 1685.280 510.000 ;
        RECT 1685.080 503.210 1685.340 503.530 ;
        RECT 1690.140 503.210 1690.400 503.530 ;
        RECT 1690.200 251.930 1690.340 503.210 ;
        RECT 1690.140 251.610 1690.400 251.930 ;
        RECT 2008.000 251.610 2008.260 251.930 ;
        RECT 2008.060 16.730 2008.200 251.610 ;
        RECT 2008.060 16.590 2012.800 16.730 ;
        RECT 2012.660 2.400 2012.800 16.590 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.910 258.640 1704.230 258.700 ;
        RECT 2028.670 258.640 2028.990 258.700 ;
        RECT 1703.910 258.500 2028.990 258.640 ;
        RECT 1703.910 258.440 1704.230 258.500 ;
        RECT 2028.670 258.440 2028.990 258.500 ;
      LAYER via ;
        RECT 1703.940 258.440 1704.200 258.700 ;
        RECT 2028.700 258.440 2028.960 258.700 ;
      LAYER met2 ;
        RECT 1701.310 510.410 1701.590 514.000 ;
        RECT 1701.310 510.270 1704.140 510.410 ;
        RECT 1701.310 510.000 1701.590 510.270 ;
        RECT 1704.000 258.730 1704.140 510.270 ;
        RECT 1703.940 258.410 1704.200 258.730 ;
        RECT 2028.700 258.410 2028.960 258.730 ;
        RECT 2028.760 17.410 2028.900 258.410 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.710 496.980 1718.030 497.040 ;
        RECT 1728.290 496.980 1728.610 497.040 ;
        RECT 1717.710 496.840 1728.610 496.980 ;
        RECT 1717.710 496.780 1718.030 496.840 ;
        RECT 1728.290 496.780 1728.610 496.840 ;
        RECT 1728.290 203.900 1728.610 203.960 ;
        RECT 2042.930 203.900 2043.250 203.960 ;
        RECT 1728.290 203.760 2043.250 203.900 ;
        RECT 1728.290 203.700 1728.610 203.760 ;
        RECT 2042.930 203.700 2043.250 203.760 ;
        RECT 2042.930 96.460 2043.250 96.520 ;
        RECT 2048.450 96.460 2048.770 96.520 ;
        RECT 2042.930 96.320 2048.770 96.460 ;
        RECT 2042.930 96.260 2043.250 96.320 ;
        RECT 2048.450 96.260 2048.770 96.320 ;
      LAYER via ;
        RECT 1717.740 496.780 1718.000 497.040 ;
        RECT 1728.320 496.780 1728.580 497.040 ;
        RECT 1728.320 203.700 1728.580 203.960 ;
        RECT 2042.960 203.700 2043.220 203.960 ;
        RECT 2042.960 96.260 2043.220 96.520 ;
        RECT 2048.480 96.260 2048.740 96.520 ;
      LAYER met2 ;
        RECT 1717.870 510.340 1718.150 514.000 ;
        RECT 1717.800 510.000 1718.150 510.340 ;
        RECT 1717.800 497.070 1717.940 510.000 ;
        RECT 1717.740 496.750 1718.000 497.070 ;
        RECT 1728.320 496.750 1728.580 497.070 ;
        RECT 1728.380 203.990 1728.520 496.750 ;
        RECT 1728.320 203.670 1728.580 203.990 ;
        RECT 2042.960 203.670 2043.220 203.990 ;
        RECT 2043.020 96.550 2043.160 203.670 ;
        RECT 2042.960 96.230 2043.220 96.550 ;
        RECT 2048.480 96.230 2048.740 96.550 ;
        RECT 2048.540 2.400 2048.680 96.230 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 544.710 189.620 545.030 189.680 ;
        RECT 759.070 189.620 759.390 189.680 ;
        RECT 544.710 189.480 759.390 189.620 ;
        RECT 544.710 189.420 545.030 189.480 ;
        RECT 759.070 189.420 759.390 189.480 ;
      LAYER via ;
        RECT 544.740 189.420 545.000 189.680 ;
        RECT 759.100 189.420 759.360 189.680 ;
      LAYER met2 ;
        RECT 542.570 510.410 542.850 514.000 ;
        RECT 542.570 510.270 544.940 510.410 ;
        RECT 542.570 510.000 542.850 510.270 ;
        RECT 544.800 189.710 544.940 510.270 ;
        RECT 544.740 189.390 545.000 189.710 ;
        RECT 759.100 189.390 759.360 189.710 ;
        RECT 759.160 16.730 759.300 189.390 ;
        RECT 759.160 16.590 763.900 16.730 ;
        RECT 763.760 2.400 763.900 16.590 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1733.810 496.980 1734.130 497.040 ;
        RECT 1738.410 496.980 1738.730 497.040 ;
        RECT 1733.810 496.840 1738.730 496.980 ;
        RECT 1733.810 496.780 1734.130 496.840 ;
        RECT 1738.410 496.780 1738.730 496.840 ;
        RECT 1738.410 306.920 1738.730 306.980 ;
        RECT 2063.170 306.920 2063.490 306.980 ;
        RECT 1738.410 306.780 2063.490 306.920 ;
        RECT 1738.410 306.720 1738.730 306.780 ;
        RECT 2063.170 306.720 2063.490 306.780 ;
        RECT 2063.170 62.120 2063.490 62.180 ;
        RECT 2066.390 62.120 2066.710 62.180 ;
        RECT 2063.170 61.980 2066.710 62.120 ;
        RECT 2063.170 61.920 2063.490 61.980 ;
        RECT 2066.390 61.920 2066.710 61.980 ;
      LAYER via ;
        RECT 1733.840 496.780 1734.100 497.040 ;
        RECT 1738.440 496.780 1738.700 497.040 ;
        RECT 1738.440 306.720 1738.700 306.980 ;
        RECT 2063.200 306.720 2063.460 306.980 ;
        RECT 2063.200 61.920 2063.460 62.180 ;
        RECT 2066.420 61.920 2066.680 62.180 ;
      LAYER met2 ;
        RECT 1733.970 510.340 1734.250 514.000 ;
        RECT 1733.900 510.000 1734.250 510.340 ;
        RECT 1733.900 497.070 1734.040 510.000 ;
        RECT 1733.840 496.750 1734.100 497.070 ;
        RECT 1738.440 496.750 1738.700 497.070 ;
        RECT 1738.500 307.010 1738.640 496.750 ;
        RECT 1738.440 306.690 1738.700 307.010 ;
        RECT 2063.200 306.690 2063.460 307.010 ;
        RECT 2063.260 62.210 2063.400 306.690 ;
        RECT 2063.200 61.890 2063.460 62.210 ;
        RECT 2066.420 61.890 2066.680 62.210 ;
        RECT 2066.480 2.400 2066.620 61.890 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1752.210 272.920 1752.530 272.980 ;
        RECT 2084.330 272.920 2084.650 272.980 ;
        RECT 1752.210 272.780 2084.650 272.920 ;
        RECT 1752.210 272.720 1752.530 272.780 ;
        RECT 2084.330 272.720 2084.650 272.780 ;
      LAYER via ;
        RECT 1752.240 272.720 1752.500 272.980 ;
        RECT 2084.360 272.720 2084.620 272.980 ;
      LAYER met2 ;
        RECT 1750.530 510.410 1750.810 514.000 ;
        RECT 1750.530 510.270 1752.440 510.410 ;
        RECT 1750.530 510.000 1750.810 510.270 ;
        RECT 1752.300 273.010 1752.440 510.270 ;
        RECT 1752.240 272.690 1752.500 273.010 ;
        RECT 2084.360 272.690 2084.620 273.010 ;
        RECT 2084.420 2.400 2084.560 272.690 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.470 500.380 1766.790 500.440 ;
        RECT 1811.090 500.380 1811.410 500.440 ;
        RECT 1766.470 500.240 1811.410 500.380 ;
        RECT 1766.470 500.180 1766.790 500.240 ;
        RECT 1811.090 500.180 1811.410 500.240 ;
        RECT 1811.090 58.720 1811.410 58.780 ;
        RECT 2097.670 58.720 2097.990 58.780 ;
        RECT 1811.090 58.580 2097.990 58.720 ;
        RECT 1811.090 58.520 1811.410 58.580 ;
        RECT 2097.670 58.520 2097.990 58.580 ;
      LAYER via ;
        RECT 1766.500 500.180 1766.760 500.440 ;
        RECT 1811.120 500.180 1811.380 500.440 ;
        RECT 1811.120 58.520 1811.380 58.780 ;
        RECT 2097.700 58.520 2097.960 58.780 ;
      LAYER met2 ;
        RECT 1766.630 510.340 1766.910 514.000 ;
        RECT 1766.560 510.000 1766.910 510.340 ;
        RECT 1766.560 500.470 1766.700 510.000 ;
        RECT 1766.500 500.150 1766.760 500.470 ;
        RECT 1811.120 500.150 1811.380 500.470 ;
        RECT 1811.180 58.810 1811.320 500.150 ;
        RECT 1811.120 58.490 1811.380 58.810 ;
        RECT 2097.700 58.490 2097.960 58.810 ;
        RECT 2097.760 17.410 2097.900 58.490 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1783.030 496.980 1783.350 497.040 ;
        RECT 1786.710 496.980 1787.030 497.040 ;
        RECT 1783.030 496.840 1787.030 496.980 ;
        RECT 1783.030 496.780 1783.350 496.840 ;
        RECT 1786.710 496.780 1787.030 496.840 ;
        RECT 1786.710 245.040 1787.030 245.100 ;
        RECT 2118.370 245.040 2118.690 245.100 ;
        RECT 1786.710 244.900 2118.690 245.040 ;
        RECT 1786.710 244.840 1787.030 244.900 ;
        RECT 2118.370 244.840 2118.690 244.900 ;
      LAYER via ;
        RECT 1783.060 496.780 1783.320 497.040 ;
        RECT 1786.740 496.780 1787.000 497.040 ;
        RECT 1786.740 244.840 1787.000 245.100 ;
        RECT 2118.400 244.840 2118.660 245.100 ;
      LAYER met2 ;
        RECT 1783.190 510.340 1783.470 514.000 ;
        RECT 1783.120 510.000 1783.470 510.340 ;
        RECT 1783.120 497.070 1783.260 510.000 ;
        RECT 1783.060 496.750 1783.320 497.070 ;
        RECT 1786.740 496.750 1787.000 497.070 ;
        RECT 1786.800 245.130 1786.940 496.750 ;
        RECT 1786.740 244.810 1787.000 245.130 ;
        RECT 2118.400 244.810 2118.660 245.130 ;
        RECT 2118.460 17.410 2118.600 244.810 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 265.440 1800.830 265.500 ;
        RECT 2132.170 265.440 2132.490 265.500 ;
        RECT 1800.510 265.300 2132.490 265.440 ;
        RECT 1800.510 265.240 1800.830 265.300 ;
        RECT 2132.170 265.240 2132.490 265.300 ;
      LAYER via ;
        RECT 1800.540 265.240 1800.800 265.500 ;
        RECT 2132.200 265.240 2132.460 265.500 ;
      LAYER met2 ;
        RECT 1799.290 510.410 1799.570 514.000 ;
        RECT 1799.290 510.270 1800.740 510.410 ;
        RECT 1799.290 510.000 1799.570 510.270 ;
        RECT 1800.600 265.530 1800.740 510.270 ;
        RECT 1800.540 265.210 1800.800 265.530 ;
        RECT 2132.200 265.210 2132.460 265.530 ;
        RECT 2132.260 17.410 2132.400 265.210 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1815.690 496.980 1816.010 497.040 ;
        RECT 1820.750 496.980 1821.070 497.040 ;
        RECT 1815.690 496.840 1821.070 496.980 ;
        RECT 1815.690 496.780 1816.010 496.840 ;
        RECT 1820.750 496.780 1821.070 496.840 ;
        RECT 1820.750 451.760 1821.070 451.820 ;
        RECT 2152.870 451.760 2153.190 451.820 ;
        RECT 1820.750 451.620 2153.190 451.760 ;
        RECT 1820.750 451.560 1821.070 451.620 ;
        RECT 2152.870 451.560 2153.190 451.620 ;
      LAYER via ;
        RECT 1815.720 496.780 1815.980 497.040 ;
        RECT 1820.780 496.780 1821.040 497.040 ;
        RECT 1820.780 451.560 1821.040 451.820 ;
        RECT 2152.900 451.560 2153.160 451.820 ;
      LAYER met2 ;
        RECT 1815.850 510.340 1816.130 514.000 ;
        RECT 1815.780 510.000 1816.130 510.340 ;
        RECT 1815.780 497.070 1815.920 510.000 ;
        RECT 1815.720 496.750 1815.980 497.070 ;
        RECT 1820.780 496.750 1821.040 497.070 ;
        RECT 1820.840 451.850 1820.980 496.750 ;
        RECT 1820.780 451.530 1821.040 451.850 ;
        RECT 2152.900 451.530 2153.160 451.850 ;
        RECT 2152.960 17.410 2153.100 451.530 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 286.180 1835.330 286.240 ;
        RECT 2166.670 286.180 2166.990 286.240 ;
        RECT 1835.010 286.040 2166.990 286.180 ;
        RECT 1835.010 285.980 1835.330 286.040 ;
        RECT 2166.670 285.980 2166.990 286.040 ;
        RECT 2166.670 16.900 2166.990 16.960 ;
        RECT 2173.110 16.900 2173.430 16.960 ;
        RECT 2166.670 16.760 2173.430 16.900 ;
        RECT 2166.670 16.700 2166.990 16.760 ;
        RECT 2173.110 16.700 2173.430 16.760 ;
      LAYER via ;
        RECT 1835.040 285.980 1835.300 286.240 ;
        RECT 2166.700 285.980 2166.960 286.240 ;
        RECT 2166.700 16.700 2166.960 16.960 ;
        RECT 2173.140 16.700 2173.400 16.960 ;
      LAYER met2 ;
        RECT 1831.950 510.410 1832.230 514.000 ;
        RECT 1831.950 510.270 1835.240 510.410 ;
        RECT 1831.950 510.000 1832.230 510.270 ;
        RECT 1835.100 286.270 1835.240 510.270 ;
        RECT 1835.040 285.950 1835.300 286.270 ;
        RECT 2166.700 285.950 2166.960 286.270 ;
        RECT 2166.760 16.990 2166.900 285.950 ;
        RECT 2166.700 16.670 2166.960 16.990 ;
        RECT 2173.140 16.670 2173.400 16.990 ;
        RECT 2173.200 2.400 2173.340 16.670 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.350 300.120 1848.670 300.180 ;
        RECT 2187.370 300.120 2187.690 300.180 ;
        RECT 1848.350 299.980 2187.690 300.120 ;
        RECT 1848.350 299.920 1848.670 299.980 ;
        RECT 2187.370 299.920 2187.690 299.980 ;
      LAYER via ;
        RECT 1848.380 299.920 1848.640 300.180 ;
        RECT 2187.400 299.920 2187.660 300.180 ;
      LAYER met2 ;
        RECT 1848.510 510.340 1848.790 514.000 ;
        RECT 1848.440 510.000 1848.790 510.340 ;
        RECT 1848.440 300.210 1848.580 510.000 ;
        RECT 1848.380 299.890 1848.640 300.210 ;
        RECT 2187.400 299.890 2187.660 300.210 ;
        RECT 2187.460 17.410 2187.600 299.890 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1864.450 496.980 1864.770 497.040 ;
        RECT 1869.510 496.980 1869.830 497.040 ;
        RECT 1864.450 496.840 1869.830 496.980 ;
        RECT 1864.450 496.780 1864.770 496.840 ;
        RECT 1869.510 496.780 1869.830 496.840 ;
        RECT 1869.510 279.380 1869.830 279.440 ;
        RECT 2208.070 279.380 2208.390 279.440 ;
        RECT 1869.510 279.240 2208.390 279.380 ;
        RECT 1869.510 279.180 1869.830 279.240 ;
        RECT 2208.070 279.180 2208.390 279.240 ;
      LAYER via ;
        RECT 1864.480 496.780 1864.740 497.040 ;
        RECT 1869.540 496.780 1869.800 497.040 ;
        RECT 1869.540 279.180 1869.800 279.440 ;
        RECT 2208.100 279.180 2208.360 279.440 ;
      LAYER met2 ;
        RECT 1864.610 510.340 1864.890 514.000 ;
        RECT 1864.540 510.000 1864.890 510.340 ;
        RECT 1864.540 497.070 1864.680 510.000 ;
        RECT 1864.480 496.750 1864.740 497.070 ;
        RECT 1869.540 496.750 1869.800 497.070 ;
        RECT 1869.600 279.470 1869.740 496.750 ;
        RECT 1869.540 279.150 1869.800 279.470 ;
        RECT 2208.100 279.150 2208.360 279.470 ;
        RECT 2208.160 17.410 2208.300 279.150 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1883.310 314.060 1883.630 314.120 ;
        RECT 2221.870 314.060 2222.190 314.120 ;
        RECT 1883.310 313.920 2222.190 314.060 ;
        RECT 1883.310 313.860 1883.630 313.920 ;
        RECT 2221.870 313.860 2222.190 313.920 ;
      LAYER via ;
        RECT 1883.340 313.860 1883.600 314.120 ;
        RECT 2221.900 313.860 2222.160 314.120 ;
      LAYER met2 ;
        RECT 1881.170 510.410 1881.450 514.000 ;
        RECT 1881.170 510.270 1883.540 510.410 ;
        RECT 1881.170 510.000 1881.450 510.270 ;
        RECT 1883.400 314.150 1883.540 510.270 ;
        RECT 1883.340 313.830 1883.600 314.150 ;
        RECT 2221.900 313.830 2222.160 314.150 ;
        RECT 2221.960 17.410 2222.100 313.830 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.970 486.440 559.290 486.500 ;
        RECT 779.770 486.440 780.090 486.500 ;
        RECT 558.970 486.300 780.090 486.440 ;
        RECT 558.970 486.240 559.290 486.300 ;
        RECT 779.770 486.240 780.090 486.300 ;
      LAYER via ;
        RECT 559.000 486.240 559.260 486.500 ;
        RECT 779.800 486.240 780.060 486.500 ;
      LAYER met2 ;
        RECT 559.130 510.340 559.410 514.000 ;
        RECT 559.060 510.000 559.410 510.340 ;
        RECT 559.060 486.530 559.200 510.000 ;
        RECT 559.000 486.210 559.260 486.530 ;
        RECT 779.800 486.210 780.060 486.530 ;
        RECT 779.860 16.730 780.000 486.210 ;
        RECT 779.860 16.590 781.840 16.730 ;
        RECT 781.700 2.400 781.840 16.590 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1897.110 293.320 1897.430 293.380 ;
        RECT 2242.570 293.320 2242.890 293.380 ;
        RECT 1897.110 293.180 2242.890 293.320 ;
        RECT 1897.110 293.120 1897.430 293.180 ;
        RECT 2242.570 293.120 2242.890 293.180 ;
      LAYER via ;
        RECT 1897.140 293.120 1897.400 293.380 ;
        RECT 2242.600 293.120 2242.860 293.380 ;
      LAYER met2 ;
        RECT 1897.270 510.340 1897.550 514.000 ;
        RECT 1897.200 510.000 1897.550 510.340 ;
        RECT 1897.200 293.410 1897.340 510.000 ;
        RECT 1897.140 293.090 1897.400 293.410 ;
        RECT 2242.600 293.090 2242.860 293.410 ;
        RECT 2242.660 17.410 2242.800 293.090 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1913.670 496.980 1913.990 497.040 ;
        RECT 1917.810 496.980 1918.130 497.040 ;
        RECT 1913.670 496.840 1918.130 496.980 ;
        RECT 1913.670 496.780 1913.990 496.840 ;
        RECT 1917.810 496.780 1918.130 496.840 ;
        RECT 1917.810 320.860 1918.130 320.920 ;
        RECT 2256.370 320.860 2256.690 320.920 ;
        RECT 1917.810 320.720 2256.690 320.860 ;
        RECT 1917.810 320.660 1918.130 320.720 ;
        RECT 2256.370 320.660 2256.690 320.720 ;
        RECT 2256.370 16.900 2256.690 16.960 ;
        RECT 2262.350 16.900 2262.670 16.960 ;
        RECT 2256.370 16.760 2262.670 16.900 ;
        RECT 2256.370 16.700 2256.690 16.760 ;
        RECT 2262.350 16.700 2262.670 16.760 ;
      LAYER via ;
        RECT 1913.700 496.780 1913.960 497.040 ;
        RECT 1917.840 496.780 1918.100 497.040 ;
        RECT 1917.840 320.660 1918.100 320.920 ;
        RECT 2256.400 320.660 2256.660 320.920 ;
        RECT 2256.400 16.700 2256.660 16.960 ;
        RECT 2262.380 16.700 2262.640 16.960 ;
      LAYER met2 ;
        RECT 1913.830 510.340 1914.110 514.000 ;
        RECT 1913.760 510.000 1914.110 510.340 ;
        RECT 1913.760 497.070 1913.900 510.000 ;
        RECT 1913.700 496.750 1913.960 497.070 ;
        RECT 1917.840 496.750 1918.100 497.070 ;
        RECT 1917.900 320.950 1918.040 496.750 ;
        RECT 1917.840 320.630 1918.100 320.950 ;
        RECT 2256.400 320.630 2256.660 320.950 ;
        RECT 2256.460 16.990 2256.600 320.630 ;
        RECT 2256.400 16.670 2256.660 16.990 ;
        RECT 2262.380 16.670 2262.640 16.990 ;
        RECT 2262.440 2.400 2262.580 16.670 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1929.770 500.380 1930.090 500.440 ;
        RECT 2059.490 500.380 2059.810 500.440 ;
        RECT 1929.770 500.240 2059.810 500.380 ;
        RECT 1929.770 500.180 1930.090 500.240 ;
        RECT 2059.490 500.180 2059.810 500.240 ;
        RECT 2059.490 93.060 2059.810 93.120 ;
        RECT 2277.070 93.060 2277.390 93.120 ;
        RECT 2059.490 92.920 2277.390 93.060 ;
        RECT 2059.490 92.860 2059.810 92.920 ;
        RECT 2277.070 92.860 2277.390 92.920 ;
      LAYER via ;
        RECT 1929.800 500.180 1930.060 500.440 ;
        RECT 2059.520 500.180 2059.780 500.440 ;
        RECT 2059.520 92.860 2059.780 93.120 ;
        RECT 2277.100 92.860 2277.360 93.120 ;
      LAYER met2 ;
        RECT 1929.930 510.340 1930.210 514.000 ;
        RECT 1929.860 510.000 1930.210 510.340 ;
        RECT 1929.860 500.470 1930.000 510.000 ;
        RECT 1929.800 500.150 1930.060 500.470 ;
        RECT 2059.520 500.150 2059.780 500.470 ;
        RECT 2059.580 93.150 2059.720 500.150 ;
        RECT 2059.520 92.830 2059.780 93.150 ;
        RECT 2277.100 92.830 2277.360 93.150 ;
        RECT 2277.160 17.410 2277.300 92.830 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1946.330 472.500 1946.650 472.560 ;
        RECT 2298.230 472.500 2298.550 472.560 ;
        RECT 1946.330 472.360 2298.550 472.500 ;
        RECT 1946.330 472.300 1946.650 472.360 ;
        RECT 2298.230 472.300 2298.550 472.360 ;
      LAYER via ;
        RECT 1946.360 472.300 1946.620 472.560 ;
        RECT 2298.260 472.300 2298.520 472.560 ;
      LAYER met2 ;
        RECT 1946.490 510.340 1946.770 514.000 ;
        RECT 1946.420 510.000 1946.770 510.340 ;
        RECT 1946.420 472.590 1946.560 510.000 ;
        RECT 1946.360 472.270 1946.620 472.590 ;
        RECT 2298.260 472.270 2298.520 472.590 ;
        RECT 2298.320 2.400 2298.460 472.270 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1962.430 503.440 1962.750 503.500 ;
        RECT 1966.110 503.440 1966.430 503.500 ;
        RECT 1962.430 503.300 1966.430 503.440 ;
        RECT 1962.430 503.240 1962.750 503.300 ;
        RECT 1966.110 503.240 1966.430 503.300 ;
        RECT 1966.110 328.000 1966.430 328.060 ;
        RECT 2311.570 328.000 2311.890 328.060 ;
        RECT 1966.110 327.860 2311.890 328.000 ;
        RECT 1966.110 327.800 1966.430 327.860 ;
        RECT 2311.570 327.800 2311.890 327.860 ;
      LAYER via ;
        RECT 1962.460 503.240 1962.720 503.500 ;
        RECT 1966.140 503.240 1966.400 503.500 ;
        RECT 1966.140 327.800 1966.400 328.060 ;
        RECT 2311.600 327.800 2311.860 328.060 ;
      LAYER met2 ;
        RECT 1962.590 510.340 1962.870 514.000 ;
        RECT 1962.520 510.000 1962.870 510.340 ;
        RECT 1962.520 503.530 1962.660 510.000 ;
        RECT 1962.460 503.210 1962.720 503.530 ;
        RECT 1966.140 503.210 1966.400 503.530 ;
        RECT 1966.200 328.090 1966.340 503.210 ;
        RECT 1966.140 327.770 1966.400 328.090 ;
        RECT 2311.600 327.770 2311.860 328.090 ;
        RECT 2311.660 17.410 2311.800 327.770 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1979.065 434.945 1979.235 483.055 ;
      LAYER mcon ;
        RECT 1979.065 482.885 1979.235 483.055 ;
      LAYER met1 ;
        RECT 1979.005 483.040 1979.295 483.085 ;
        RECT 1979.450 483.040 1979.770 483.100 ;
        RECT 1979.005 482.900 1979.770 483.040 ;
        RECT 1979.005 482.855 1979.295 482.900 ;
        RECT 1979.450 482.840 1979.770 482.900 ;
        RECT 1978.990 435.100 1979.310 435.160 ;
        RECT 1978.795 434.960 1979.310 435.100 ;
        RECT 1978.990 434.900 1979.310 434.960 ;
        RECT 1978.990 400.560 1979.310 400.820 ;
        RECT 1979.080 400.140 1979.220 400.560 ;
        RECT 1978.990 399.880 1979.310 400.140 ;
        RECT 1978.990 334.800 1979.310 334.860 ;
        RECT 2332.270 334.800 2332.590 334.860 ;
        RECT 1978.990 334.660 2332.590 334.800 ;
        RECT 1978.990 334.600 1979.310 334.660 ;
        RECT 2332.270 334.600 2332.590 334.660 ;
      LAYER via ;
        RECT 1979.480 482.840 1979.740 483.100 ;
        RECT 1979.020 434.900 1979.280 435.160 ;
        RECT 1979.020 400.560 1979.280 400.820 ;
        RECT 1979.020 399.880 1979.280 400.140 ;
        RECT 1979.020 334.600 1979.280 334.860 ;
        RECT 2332.300 334.600 2332.560 334.860 ;
      LAYER met2 ;
        RECT 1979.150 511.090 1979.430 514.000 ;
        RECT 1979.150 510.950 1980.140 511.090 ;
        RECT 1979.150 510.000 1979.430 510.950 ;
        RECT 1980.000 498.680 1980.140 510.950 ;
        RECT 1979.540 498.540 1980.140 498.680 ;
        RECT 1979.540 483.130 1979.680 498.540 ;
        RECT 1979.480 482.810 1979.740 483.130 ;
        RECT 1979.020 434.870 1979.280 435.190 ;
        RECT 1979.080 400.850 1979.220 434.870 ;
        RECT 1979.020 400.530 1979.280 400.850 ;
        RECT 1979.020 399.850 1979.280 400.170 ;
        RECT 1979.080 334.890 1979.220 399.850 ;
        RECT 1979.020 334.570 1979.280 334.890 ;
        RECT 2332.300 334.570 2332.560 334.890 ;
        RECT 2332.360 17.410 2332.500 334.570 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 496.980 1995.410 497.040 ;
        RECT 2000.150 496.980 2000.470 497.040 ;
        RECT 1995.090 496.840 2000.470 496.980 ;
        RECT 1995.090 496.780 1995.410 496.840 ;
        RECT 2000.150 496.780 2000.470 496.840 ;
        RECT 2000.150 237.900 2000.470 237.960 ;
        RECT 2346.070 237.900 2346.390 237.960 ;
        RECT 2000.150 237.760 2346.390 237.900 ;
        RECT 2000.150 237.700 2000.470 237.760 ;
        RECT 2346.070 237.700 2346.390 237.760 ;
      LAYER via ;
        RECT 1995.120 496.780 1995.380 497.040 ;
        RECT 2000.180 496.780 2000.440 497.040 ;
        RECT 2000.180 237.700 2000.440 237.960 ;
        RECT 2346.100 237.700 2346.360 237.960 ;
      LAYER met2 ;
        RECT 1995.250 510.340 1995.530 514.000 ;
        RECT 1995.180 510.000 1995.530 510.340 ;
        RECT 1995.180 497.070 1995.320 510.000 ;
        RECT 1995.120 496.750 1995.380 497.070 ;
        RECT 2000.180 496.750 2000.440 497.070 ;
        RECT 2000.240 237.990 2000.380 496.750 ;
        RECT 2000.180 237.670 2000.440 237.990 ;
        RECT 2346.100 237.670 2346.360 237.990 ;
        RECT 2346.160 17.410 2346.300 237.670 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 341.600 2014.730 341.660 ;
        RECT 2366.770 341.600 2367.090 341.660 ;
        RECT 2014.410 341.460 2367.090 341.600 ;
        RECT 2014.410 341.400 2014.730 341.460 ;
        RECT 2366.770 341.400 2367.090 341.460 ;
      LAYER via ;
        RECT 2014.440 341.400 2014.700 341.660 ;
        RECT 2366.800 341.400 2367.060 341.660 ;
      LAYER met2 ;
        RECT 2011.350 510.410 2011.630 514.000 ;
        RECT 2011.350 510.270 2014.640 510.410 ;
        RECT 2011.350 510.000 2011.630 510.270 ;
        RECT 2014.500 341.690 2014.640 510.270 ;
        RECT 2014.440 341.370 2014.700 341.690 ;
        RECT 2366.800 341.370 2367.060 341.690 ;
        RECT 2366.860 16.730 2367.000 341.370 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2027.750 348.400 2028.070 348.460 ;
        RECT 2387.930 348.400 2388.250 348.460 ;
        RECT 2027.750 348.260 2388.250 348.400 ;
        RECT 2027.750 348.200 2028.070 348.260 ;
        RECT 2387.930 348.200 2388.250 348.260 ;
      LAYER via ;
        RECT 2027.780 348.200 2028.040 348.460 ;
        RECT 2387.960 348.200 2388.220 348.460 ;
      LAYER met2 ;
        RECT 2027.910 510.340 2028.190 514.000 ;
        RECT 2027.840 510.000 2028.190 510.340 ;
        RECT 2027.840 348.490 2027.980 510.000 ;
        RECT 2027.780 348.170 2028.040 348.490 ;
        RECT 2387.960 348.170 2388.220 348.490 ;
        RECT 2388.020 17.410 2388.160 348.170 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2043.850 503.440 2044.170 503.500 ;
        RECT 2048.910 503.440 2049.230 503.500 ;
        RECT 2043.850 503.300 2049.230 503.440 ;
        RECT 2043.850 503.240 2044.170 503.300 ;
        RECT 2048.910 503.240 2049.230 503.300 ;
        RECT 2048.910 355.200 2049.230 355.260 ;
        RECT 2401.270 355.200 2401.590 355.260 ;
        RECT 2048.910 355.060 2401.590 355.200 ;
        RECT 2048.910 355.000 2049.230 355.060 ;
        RECT 2401.270 355.000 2401.590 355.060 ;
      LAYER via ;
        RECT 2043.880 503.240 2044.140 503.500 ;
        RECT 2048.940 503.240 2049.200 503.500 ;
        RECT 2048.940 355.000 2049.200 355.260 ;
        RECT 2401.300 355.000 2401.560 355.260 ;
      LAYER met2 ;
        RECT 2044.010 510.340 2044.290 514.000 ;
        RECT 2043.940 510.000 2044.290 510.340 ;
        RECT 2043.940 503.530 2044.080 510.000 ;
        RECT 2043.880 503.210 2044.140 503.530 ;
        RECT 2048.940 503.210 2049.200 503.530 ;
        RECT 2049.000 355.290 2049.140 503.210 ;
        RECT 2048.940 354.970 2049.200 355.290 ;
        RECT 2401.300 354.970 2401.560 355.290 ;
        RECT 2401.360 17.410 2401.500 354.970 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 575.070 496.980 575.390 497.040 ;
        RECT 579.210 496.980 579.530 497.040 ;
        RECT 575.070 496.840 579.530 496.980 ;
        RECT 575.070 496.780 575.390 496.840 ;
        RECT 579.210 496.780 579.530 496.840 ;
        RECT 579.210 196.760 579.530 196.820 ;
        RECT 793.570 196.760 793.890 196.820 ;
        RECT 579.210 196.620 793.890 196.760 ;
        RECT 579.210 196.560 579.530 196.620 ;
        RECT 793.570 196.560 793.890 196.620 ;
        RECT 793.570 17.580 793.890 17.640 ;
        RECT 799.550 17.580 799.870 17.640 ;
        RECT 793.570 17.440 799.870 17.580 ;
        RECT 793.570 17.380 793.890 17.440 ;
        RECT 799.550 17.380 799.870 17.440 ;
      LAYER via ;
        RECT 575.100 496.780 575.360 497.040 ;
        RECT 579.240 496.780 579.500 497.040 ;
        RECT 579.240 196.560 579.500 196.820 ;
        RECT 793.600 196.560 793.860 196.820 ;
        RECT 793.600 17.380 793.860 17.640 ;
        RECT 799.580 17.380 799.840 17.640 ;
      LAYER met2 ;
        RECT 575.230 510.340 575.510 514.000 ;
        RECT 575.160 510.000 575.510 510.340 ;
        RECT 575.160 497.070 575.300 510.000 ;
        RECT 575.100 496.750 575.360 497.070 ;
        RECT 579.240 496.750 579.500 497.070 ;
        RECT 579.300 196.850 579.440 496.750 ;
        RECT 579.240 196.530 579.500 196.850 ;
        RECT 793.600 196.530 793.860 196.850 ;
        RECT 793.660 17.670 793.800 196.530 ;
        RECT 793.600 17.350 793.860 17.670 ;
        RECT 799.580 17.350 799.840 17.670 ;
        RECT 799.640 2.400 799.780 17.350 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 434.310 38.320 434.630 38.380 ;
        RECT 644.530 38.320 644.850 38.380 ;
        RECT 434.310 38.180 644.850 38.320 ;
        RECT 434.310 38.120 434.630 38.180 ;
        RECT 644.530 38.120 644.850 38.180 ;
      LAYER via ;
        RECT 434.340 38.120 434.600 38.380 ;
        RECT 644.560 38.120 644.820 38.380 ;
      LAYER met2 ;
        RECT 434.010 510.410 434.290 514.000 ;
        RECT 433.480 510.270 434.290 510.410 ;
        RECT 433.480 483.325 433.620 510.270 ;
        RECT 434.010 510.000 434.290 510.270 ;
        RECT 433.410 482.955 433.690 483.325 ;
        RECT 434.330 482.955 434.610 483.325 ;
        RECT 434.400 38.410 434.540 482.955 ;
        RECT 434.340 38.090 434.600 38.410 ;
        RECT 644.560 38.090 644.820 38.410 ;
        RECT 644.620 17.410 644.760 38.090 ;
        RECT 644.620 17.270 645.220 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 433.410 483.000 433.690 483.280 ;
        RECT 434.330 483.000 434.610 483.280 ;
      LAYER met3 ;
        RECT 433.385 483.290 433.715 483.305 ;
        RECT 434.305 483.290 434.635 483.305 ;
        RECT 433.385 482.990 434.635 483.290 ;
        RECT 433.385 482.975 433.715 482.990 ;
        RECT 434.305 482.975 434.635 482.990 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.610 306.920 2069.930 306.980 ;
        RECT 2428.870 306.920 2429.190 306.980 ;
        RECT 2069.610 306.780 2429.190 306.920 ;
        RECT 2069.610 306.720 2069.930 306.780 ;
        RECT 2428.870 306.720 2429.190 306.780 ;
      LAYER via ;
        RECT 2069.640 306.720 2069.900 306.980 ;
        RECT 2428.900 306.720 2429.160 306.980 ;
      LAYER met2 ;
        RECT 2066.090 510.410 2066.370 514.000 ;
        RECT 2066.090 510.270 2069.840 510.410 ;
        RECT 2066.090 510.000 2066.370 510.270 ;
        RECT 2069.700 307.010 2069.840 510.270 ;
        RECT 2069.640 306.690 2069.900 307.010 ;
        RECT 2428.900 306.690 2429.160 307.010 ;
        RECT 2428.960 2.400 2429.100 306.690 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 272.580 2083.730 272.640 ;
        RECT 2442.670 272.580 2442.990 272.640 ;
        RECT 2083.410 272.440 2442.990 272.580 ;
        RECT 2083.410 272.380 2083.730 272.440 ;
        RECT 2442.670 272.380 2442.990 272.440 ;
      LAYER via ;
        RECT 2083.440 272.380 2083.700 272.640 ;
        RECT 2442.700 272.380 2442.960 272.640 ;
      LAYER met2 ;
        RECT 2082.190 510.410 2082.470 514.000 ;
        RECT 2082.190 510.270 2083.640 510.410 ;
        RECT 2082.190 510.000 2082.470 510.270 ;
        RECT 2083.500 272.670 2083.640 510.270 ;
        RECT 2083.440 272.350 2083.700 272.670 ;
        RECT 2442.700 272.350 2442.960 272.670 ;
        RECT 2442.760 17.410 2442.900 272.350 ;
        RECT 2442.760 17.270 2447.040 17.410 ;
        RECT 2446.900 2.400 2447.040 17.270 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2098.590 499.020 2098.910 499.080 ;
        RECT 2103.650 499.020 2103.970 499.080 ;
        RECT 2098.590 498.880 2103.970 499.020 ;
        RECT 2098.590 498.820 2098.910 498.880 ;
        RECT 2103.650 498.820 2103.970 498.880 ;
        RECT 2103.650 362.340 2103.970 362.400 ;
        RECT 2463.370 362.340 2463.690 362.400 ;
        RECT 2103.650 362.200 2463.690 362.340 ;
        RECT 2103.650 362.140 2103.970 362.200 ;
        RECT 2463.370 362.140 2463.690 362.200 ;
      LAYER via ;
        RECT 2098.620 498.820 2098.880 499.080 ;
        RECT 2103.680 498.820 2103.940 499.080 ;
        RECT 2103.680 362.140 2103.940 362.400 ;
        RECT 2463.400 362.140 2463.660 362.400 ;
      LAYER met2 ;
        RECT 2098.750 510.340 2099.030 514.000 ;
        RECT 2098.680 510.000 2099.030 510.340 ;
        RECT 2098.680 499.110 2098.820 510.000 ;
        RECT 2098.620 498.790 2098.880 499.110 ;
        RECT 2103.680 498.790 2103.940 499.110 ;
        RECT 2103.740 362.430 2103.880 498.790 ;
        RECT 2103.680 362.110 2103.940 362.430 ;
        RECT 2463.400 362.110 2463.660 362.430 ;
        RECT 2463.460 18.090 2463.600 362.110 ;
        RECT 2463.460 17.950 2464.980 18.090 ;
        RECT 2464.840 2.400 2464.980 17.950 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2477.245 241.485 2477.415 289.595 ;
        RECT 2477.245 144.925 2477.415 193.035 ;
        RECT 2482.765 2.805 2482.935 48.195 ;
      LAYER mcon ;
        RECT 2477.245 289.425 2477.415 289.595 ;
        RECT 2477.245 192.865 2477.415 193.035 ;
        RECT 2482.765 48.025 2482.935 48.195 ;
      LAYER met1 ;
        RECT 2117.910 369.140 2118.230 369.200 ;
        RECT 2477.170 369.140 2477.490 369.200 ;
        RECT 2117.910 369.000 2477.490 369.140 ;
        RECT 2117.910 368.940 2118.230 369.000 ;
        RECT 2477.170 368.940 2477.490 369.000 ;
        RECT 2477.170 289.580 2477.490 289.640 ;
        RECT 2476.975 289.440 2477.490 289.580 ;
        RECT 2477.170 289.380 2477.490 289.440 ;
        RECT 2477.170 241.640 2477.490 241.700 ;
        RECT 2476.975 241.500 2477.490 241.640 ;
        RECT 2477.170 241.440 2477.490 241.500 ;
        RECT 2477.170 193.020 2477.490 193.080 ;
        RECT 2476.975 192.880 2477.490 193.020 ;
        RECT 2477.170 192.820 2477.490 192.880 ;
        RECT 2477.170 145.080 2477.490 145.140 ;
        RECT 2476.975 144.940 2477.490 145.080 ;
        RECT 2477.170 144.880 2477.490 144.940 ;
        RECT 2477.170 96.460 2477.490 96.520 ;
        RECT 2478.090 96.460 2478.410 96.520 ;
        RECT 2477.170 96.320 2478.410 96.460 ;
        RECT 2477.170 96.260 2477.490 96.320 ;
        RECT 2478.090 96.260 2478.410 96.320 ;
        RECT 2477.170 48.180 2477.490 48.240 ;
        RECT 2482.705 48.180 2482.995 48.225 ;
        RECT 2477.170 48.040 2482.995 48.180 ;
        RECT 2477.170 47.980 2477.490 48.040 ;
        RECT 2482.705 47.995 2482.995 48.040 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2482.495 2.820 2483.010 2.960 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 2117.940 368.940 2118.200 369.200 ;
        RECT 2477.200 368.940 2477.460 369.200 ;
        RECT 2477.200 289.380 2477.460 289.640 ;
        RECT 2477.200 241.440 2477.460 241.700 ;
        RECT 2477.200 192.820 2477.460 193.080 ;
        RECT 2477.200 144.880 2477.460 145.140 ;
        RECT 2477.200 96.260 2477.460 96.520 ;
        RECT 2478.120 96.260 2478.380 96.520 ;
        RECT 2477.200 47.980 2477.460 48.240 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 2114.850 510.410 2115.130 514.000 ;
        RECT 2114.850 510.270 2118.140 510.410 ;
        RECT 2114.850 510.000 2115.130 510.270 ;
        RECT 2118.000 369.230 2118.140 510.270 ;
        RECT 2117.940 368.910 2118.200 369.230 ;
        RECT 2477.200 368.910 2477.460 369.230 ;
        RECT 2477.260 290.885 2477.400 368.910 ;
        RECT 2477.190 290.515 2477.470 290.885 ;
        RECT 2477.190 289.835 2477.470 290.205 ;
        RECT 2477.260 289.670 2477.400 289.835 ;
        RECT 2477.200 289.350 2477.460 289.670 ;
        RECT 2477.200 241.410 2477.460 241.730 ;
        RECT 2477.260 193.110 2477.400 241.410 ;
        RECT 2477.200 192.790 2477.460 193.110 ;
        RECT 2477.200 144.850 2477.460 145.170 ;
        RECT 2477.260 96.550 2477.400 144.850 ;
        RECT 2477.200 96.230 2477.460 96.550 ;
        RECT 2478.120 96.230 2478.380 96.550 ;
        RECT 2478.180 48.805 2478.320 96.230 ;
        RECT 2477.190 48.435 2477.470 48.805 ;
        RECT 2478.110 48.435 2478.390 48.805 ;
        RECT 2477.260 48.270 2477.400 48.435 ;
        RECT 2477.200 47.950 2477.460 48.270 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
      LAYER via2 ;
        RECT 2477.190 290.560 2477.470 290.840 ;
        RECT 2477.190 289.880 2477.470 290.160 ;
        RECT 2477.190 48.480 2477.470 48.760 ;
        RECT 2478.110 48.480 2478.390 48.760 ;
      LAYER met3 ;
        RECT 2477.165 290.850 2477.495 290.865 ;
        RECT 2477.165 290.550 2478.170 290.850 ;
        RECT 2477.165 290.535 2477.495 290.550 ;
        RECT 2477.165 290.170 2477.495 290.185 ;
        RECT 2477.870 290.170 2478.170 290.550 ;
        RECT 2477.165 289.870 2478.170 290.170 ;
        RECT 2477.165 289.855 2477.495 289.870 ;
        RECT 2477.165 48.770 2477.495 48.785 ;
        RECT 2478.085 48.770 2478.415 48.785 ;
        RECT 2477.165 48.470 2478.415 48.770 ;
        RECT 2477.165 48.455 2477.495 48.470 ;
        RECT 2478.085 48.455 2478.415 48.470 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2497.945 289.765 2498.115 337.875 ;
      LAYER mcon ;
        RECT 2497.945 337.705 2498.115 337.875 ;
      LAYER met1 ;
        RECT 2131.710 375.940 2132.030 376.000 ;
        RECT 2497.870 375.940 2498.190 376.000 ;
        RECT 2131.710 375.800 2498.190 375.940 ;
        RECT 2131.710 375.740 2132.030 375.800 ;
        RECT 2497.870 375.740 2498.190 375.800 ;
        RECT 2497.870 337.860 2498.190 337.920 ;
        RECT 2497.675 337.720 2498.190 337.860 ;
        RECT 2497.870 337.660 2498.190 337.720 ;
        RECT 2497.870 289.920 2498.190 289.980 ;
        RECT 2497.675 289.780 2498.190 289.920 ;
        RECT 2497.870 289.720 2498.190 289.780 ;
        RECT 2497.870 14.180 2498.190 14.240 ;
        RECT 2497.870 14.040 2500.860 14.180 ;
        RECT 2497.870 13.980 2498.190 14.040 ;
        RECT 2500.720 13.900 2500.860 14.040 ;
        RECT 2500.630 13.640 2500.950 13.900 ;
      LAYER via ;
        RECT 2131.740 375.740 2132.000 376.000 ;
        RECT 2497.900 375.740 2498.160 376.000 ;
        RECT 2497.900 337.660 2498.160 337.920 ;
        RECT 2497.900 289.720 2498.160 289.980 ;
        RECT 2497.900 13.980 2498.160 14.240 ;
        RECT 2500.660 13.640 2500.920 13.900 ;
      LAYER met2 ;
        RECT 2131.410 511.770 2131.690 514.000 ;
        RECT 2131.410 511.630 2132.400 511.770 ;
        RECT 2131.410 510.000 2131.690 511.630 ;
        RECT 2132.260 494.770 2132.400 511.630 ;
        RECT 2131.800 494.630 2132.400 494.770 ;
        RECT 2131.800 376.030 2131.940 494.630 ;
        RECT 2131.740 375.710 2132.000 376.030 ;
        RECT 2497.900 375.710 2498.160 376.030 ;
        RECT 2497.960 337.950 2498.100 375.710 ;
        RECT 2497.900 337.630 2498.160 337.950 ;
        RECT 2497.900 289.690 2498.160 290.010 ;
        RECT 2497.960 14.270 2498.100 289.690 ;
        RECT 2497.900 13.950 2498.160 14.270 ;
        RECT 2500.660 13.610 2500.920 13.930 ;
        RECT 2500.720 2.400 2500.860 13.610 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2147.350 496.980 2147.670 497.040 ;
        RECT 2152.410 496.980 2152.730 497.040 ;
        RECT 2147.350 496.840 2152.730 496.980 ;
        RECT 2147.350 496.780 2147.670 496.840 ;
        RECT 2152.410 496.780 2152.730 496.840 ;
        RECT 2152.410 382.740 2152.730 382.800 ;
        RECT 2511.670 382.740 2511.990 382.800 ;
        RECT 2152.410 382.600 2511.990 382.740 ;
        RECT 2152.410 382.540 2152.730 382.600 ;
        RECT 2511.670 382.540 2511.990 382.600 ;
        RECT 2511.670 10.440 2511.990 10.500 ;
        RECT 2518.110 10.440 2518.430 10.500 ;
        RECT 2511.670 10.300 2518.430 10.440 ;
        RECT 2511.670 10.240 2511.990 10.300 ;
        RECT 2518.110 10.240 2518.430 10.300 ;
      LAYER via ;
        RECT 2147.380 496.780 2147.640 497.040 ;
        RECT 2152.440 496.780 2152.700 497.040 ;
        RECT 2152.440 382.540 2152.700 382.800 ;
        RECT 2511.700 382.540 2511.960 382.800 ;
        RECT 2511.700 10.240 2511.960 10.500 ;
        RECT 2518.140 10.240 2518.400 10.500 ;
      LAYER met2 ;
        RECT 2147.510 510.340 2147.790 514.000 ;
        RECT 2147.440 510.000 2147.790 510.340 ;
        RECT 2147.440 497.070 2147.580 510.000 ;
        RECT 2147.380 496.750 2147.640 497.070 ;
        RECT 2152.440 496.750 2152.700 497.070 ;
        RECT 2152.500 382.830 2152.640 496.750 ;
        RECT 2152.440 382.510 2152.700 382.830 ;
        RECT 2511.700 382.510 2511.960 382.830 ;
        RECT 2511.760 10.530 2511.900 382.510 ;
        RECT 2511.700 10.210 2511.960 10.530 ;
        RECT 2518.140 10.210 2518.400 10.530 ;
        RECT 2518.200 2.400 2518.340 10.210 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 410.620 2166.530 410.680 ;
        RECT 2532.370 410.620 2532.690 410.680 ;
        RECT 2166.210 410.480 2532.690 410.620 ;
        RECT 2166.210 410.420 2166.530 410.480 ;
        RECT 2532.370 410.420 2532.690 410.480 ;
      LAYER via ;
        RECT 2166.240 410.420 2166.500 410.680 ;
        RECT 2532.400 410.420 2532.660 410.680 ;
      LAYER met2 ;
        RECT 2164.070 510.410 2164.350 514.000 ;
        RECT 2164.070 510.270 2166.440 510.410 ;
        RECT 2164.070 510.000 2164.350 510.270 ;
        RECT 2166.300 410.710 2166.440 510.270 ;
        RECT 2166.240 410.390 2166.500 410.710 ;
        RECT 2532.400 410.390 2532.660 410.710 ;
        RECT 2532.460 17.410 2532.600 410.390 ;
        RECT 2532.460 17.270 2536.280 17.410 ;
        RECT 2536.140 2.400 2536.280 17.270 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 286.180 2180.330 286.240 ;
        RECT 2553.070 286.180 2553.390 286.240 ;
        RECT 2180.010 286.040 2553.390 286.180 ;
        RECT 2180.010 285.980 2180.330 286.040 ;
        RECT 2553.070 285.980 2553.390 286.040 ;
      LAYER via ;
        RECT 2180.040 285.980 2180.300 286.240 ;
        RECT 2553.100 285.980 2553.360 286.240 ;
      LAYER met2 ;
        RECT 2180.170 510.340 2180.450 514.000 ;
        RECT 2180.100 510.000 2180.450 510.340 ;
        RECT 2180.100 286.270 2180.240 510.000 ;
        RECT 2180.040 285.950 2180.300 286.270 ;
        RECT 2553.100 285.950 2553.360 286.270 ;
        RECT 2553.160 17.410 2553.300 285.950 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2196.570 496.980 2196.890 497.040 ;
        RECT 2200.710 496.980 2201.030 497.040 ;
        RECT 2196.570 496.840 2201.030 496.980 ;
        RECT 2196.570 496.780 2196.890 496.840 ;
        RECT 2200.710 496.780 2201.030 496.840 ;
        RECT 2200.710 300.120 2201.030 300.180 ;
        RECT 2566.870 300.120 2567.190 300.180 ;
        RECT 2200.710 299.980 2567.190 300.120 ;
        RECT 2200.710 299.920 2201.030 299.980 ;
        RECT 2566.870 299.920 2567.190 299.980 ;
      LAYER via ;
        RECT 2196.600 496.780 2196.860 497.040 ;
        RECT 2200.740 496.780 2201.000 497.040 ;
        RECT 2200.740 299.920 2201.000 300.180 ;
        RECT 2566.900 299.920 2567.160 300.180 ;
      LAYER met2 ;
        RECT 2196.730 510.340 2197.010 514.000 ;
        RECT 2196.660 510.000 2197.010 510.340 ;
        RECT 2196.660 497.070 2196.800 510.000 ;
        RECT 2196.600 496.750 2196.860 497.070 ;
        RECT 2200.740 496.750 2201.000 497.070 ;
        RECT 2200.800 300.210 2200.940 496.750 ;
        RECT 2200.740 299.890 2201.000 300.210 ;
        RECT 2566.900 299.890 2567.160 300.210 ;
        RECT 2566.960 17.410 2567.100 299.890 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.400 2572.160 17.270 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 279.380 2214.830 279.440 ;
        RECT 2587.570 279.380 2587.890 279.440 ;
        RECT 2214.510 279.240 2587.890 279.380 ;
        RECT 2214.510 279.180 2214.830 279.240 ;
        RECT 2587.570 279.180 2587.890 279.240 ;
      LAYER via ;
        RECT 2214.540 279.180 2214.800 279.440 ;
        RECT 2587.600 279.180 2587.860 279.440 ;
      LAYER met2 ;
        RECT 2212.830 510.410 2213.110 514.000 ;
        RECT 2212.830 510.270 2214.740 510.410 ;
        RECT 2212.830 510.000 2213.110 510.270 ;
        RECT 2214.600 279.470 2214.740 510.270 ;
        RECT 2214.540 279.150 2214.800 279.470 ;
        RECT 2587.600 279.150 2587.860 279.470 ;
        RECT 2587.660 17.410 2587.800 279.150 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 203.560 600.230 203.620 ;
        RECT 821.170 203.560 821.490 203.620 ;
        RECT 599.910 203.420 821.490 203.560 ;
        RECT 599.910 203.360 600.230 203.420 ;
        RECT 821.170 203.360 821.490 203.420 ;
      LAYER via ;
        RECT 599.940 203.360 600.200 203.620 ;
        RECT 821.200 203.360 821.460 203.620 ;
      LAYER met2 ;
        RECT 597.310 510.410 597.590 514.000 ;
        RECT 597.310 510.270 600.140 510.410 ;
        RECT 597.310 510.000 597.590 510.270 ;
        RECT 600.000 203.650 600.140 510.270 ;
        RECT 599.940 203.330 600.200 203.650 ;
        RECT 821.200 203.330 821.460 203.650 ;
        RECT 821.260 17.410 821.400 203.330 ;
        RECT 821.260 17.270 823.700 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2229.230 496.980 2229.550 497.040 ;
        RECT 2235.210 496.980 2235.530 497.040 ;
        RECT 2229.230 496.840 2235.530 496.980 ;
        RECT 2229.230 496.780 2229.550 496.840 ;
        RECT 2235.210 496.780 2235.530 496.840 ;
        RECT 2235.210 314.060 2235.530 314.120 ;
        RECT 2601.370 314.060 2601.690 314.120 ;
        RECT 2235.210 313.920 2601.690 314.060 ;
        RECT 2235.210 313.860 2235.530 313.920 ;
        RECT 2601.370 313.860 2601.690 313.920 ;
        RECT 2601.370 20.980 2601.690 21.040 ;
        RECT 2607.350 20.980 2607.670 21.040 ;
        RECT 2601.370 20.840 2607.670 20.980 ;
        RECT 2601.370 20.780 2601.690 20.840 ;
        RECT 2607.350 20.780 2607.670 20.840 ;
      LAYER via ;
        RECT 2229.260 496.780 2229.520 497.040 ;
        RECT 2235.240 496.780 2235.500 497.040 ;
        RECT 2235.240 313.860 2235.500 314.120 ;
        RECT 2601.400 313.860 2601.660 314.120 ;
        RECT 2601.400 20.780 2601.660 21.040 ;
        RECT 2607.380 20.780 2607.640 21.040 ;
      LAYER met2 ;
        RECT 2229.390 510.340 2229.670 514.000 ;
        RECT 2229.320 510.000 2229.670 510.340 ;
        RECT 2229.320 497.070 2229.460 510.000 ;
        RECT 2229.260 496.750 2229.520 497.070 ;
        RECT 2235.240 496.750 2235.500 497.070 ;
        RECT 2235.300 314.150 2235.440 496.750 ;
        RECT 2235.240 313.830 2235.500 314.150 ;
        RECT 2601.400 313.830 2601.660 314.150 ;
        RECT 2601.460 21.070 2601.600 313.830 ;
        RECT 2601.400 20.750 2601.660 21.070 ;
        RECT 2607.380 20.750 2607.640 21.070 ;
        RECT 2607.440 2.400 2607.580 20.750 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2249.010 293.320 2249.330 293.380 ;
        RECT 2622.070 293.320 2622.390 293.380 ;
        RECT 2249.010 293.180 2622.390 293.320 ;
        RECT 2249.010 293.120 2249.330 293.180 ;
        RECT 2622.070 293.120 2622.390 293.180 ;
      LAYER via ;
        RECT 2249.040 293.120 2249.300 293.380 ;
        RECT 2622.100 293.120 2622.360 293.380 ;
      LAYER met2 ;
        RECT 2245.490 510.410 2245.770 514.000 ;
        RECT 2245.490 510.270 2249.240 510.410 ;
        RECT 2245.490 510.000 2245.770 510.270 ;
        RECT 2249.100 293.410 2249.240 510.270 ;
        RECT 2249.040 293.090 2249.300 293.410 ;
        RECT 2622.100 293.090 2622.360 293.410 ;
        RECT 2622.160 17.410 2622.300 293.090 ;
        RECT 2622.160 17.270 2625.520 17.410 ;
        RECT 2625.380 2.400 2625.520 17.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2262.350 403.480 2262.670 403.540 ;
        RECT 2642.770 403.480 2643.090 403.540 ;
        RECT 2262.350 403.340 2643.090 403.480 ;
        RECT 2262.350 403.280 2262.670 403.340 ;
        RECT 2642.770 403.280 2643.090 403.340 ;
      LAYER via ;
        RECT 2262.380 403.280 2262.640 403.540 ;
        RECT 2642.800 403.280 2643.060 403.540 ;
      LAYER met2 ;
        RECT 2261.590 510.410 2261.870 514.000 ;
        RECT 2261.590 510.270 2262.580 510.410 ;
        RECT 2261.590 510.000 2261.870 510.270 ;
        RECT 2262.440 403.570 2262.580 510.270 ;
        RECT 2262.380 403.250 2262.640 403.570 ;
        RECT 2642.800 403.250 2643.060 403.570 ;
        RECT 2642.860 17.410 2643.000 403.250 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2277.990 496.980 2278.310 497.040 ;
        RECT 2283.050 496.980 2283.370 497.040 ;
        RECT 2277.990 496.840 2283.370 496.980 ;
        RECT 2277.990 496.780 2278.310 496.840 ;
        RECT 2283.050 496.780 2283.370 496.840 ;
        RECT 2283.050 396.680 2283.370 396.740 ;
        RECT 2656.570 396.680 2656.890 396.740 ;
        RECT 2283.050 396.540 2656.890 396.680 ;
        RECT 2283.050 396.480 2283.370 396.540 ;
        RECT 2656.570 396.480 2656.890 396.540 ;
      LAYER via ;
        RECT 2278.020 496.780 2278.280 497.040 ;
        RECT 2283.080 496.780 2283.340 497.040 ;
        RECT 2283.080 396.480 2283.340 396.740 ;
        RECT 2656.600 396.480 2656.860 396.740 ;
      LAYER met2 ;
        RECT 2278.150 510.340 2278.430 514.000 ;
        RECT 2278.080 510.000 2278.430 510.340 ;
        RECT 2278.080 497.070 2278.220 510.000 ;
        RECT 2278.020 496.750 2278.280 497.070 ;
        RECT 2283.080 496.750 2283.340 497.070 ;
        RECT 2283.140 396.770 2283.280 496.750 ;
        RECT 2283.080 396.450 2283.340 396.770 ;
        RECT 2656.600 396.450 2656.860 396.770 ;
        RECT 2656.660 17.410 2656.800 396.450 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2297.310 389.880 2297.630 389.940 ;
        RECT 2677.270 389.880 2677.590 389.940 ;
        RECT 2297.310 389.740 2677.590 389.880 ;
        RECT 2297.310 389.680 2297.630 389.740 ;
        RECT 2677.270 389.680 2677.590 389.740 ;
      LAYER via ;
        RECT 2297.340 389.680 2297.600 389.940 ;
        RECT 2677.300 389.680 2677.560 389.940 ;
      LAYER met2 ;
        RECT 2294.250 510.410 2294.530 514.000 ;
        RECT 2294.250 510.270 2297.540 510.410 ;
        RECT 2294.250 510.000 2294.530 510.270 ;
        RECT 2297.400 389.970 2297.540 510.270 ;
        RECT 2297.340 389.650 2297.600 389.970 ;
        RECT 2677.300 389.650 2677.560 389.970 ;
        RECT 2677.360 17.410 2677.500 389.650 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2310.190 448.700 2310.510 448.760 ;
        RECT 2311.110 448.700 2311.430 448.760 ;
        RECT 2310.190 448.560 2311.430 448.700 ;
        RECT 2310.190 448.500 2310.510 448.560 ;
        RECT 2311.110 448.500 2311.430 448.560 ;
        RECT 2310.650 400.560 2310.970 400.820 ;
        RECT 2310.740 400.140 2310.880 400.560 ;
        RECT 2310.650 399.880 2310.970 400.140 ;
        RECT 2310.190 327.660 2310.510 327.720 ;
        RECT 2691.070 327.660 2691.390 327.720 ;
        RECT 2310.190 327.520 2691.390 327.660 ;
        RECT 2310.190 327.460 2310.510 327.520 ;
        RECT 2691.070 327.460 2691.390 327.520 ;
      LAYER via ;
        RECT 2310.220 448.500 2310.480 448.760 ;
        RECT 2311.140 448.500 2311.400 448.760 ;
        RECT 2310.680 400.560 2310.940 400.820 ;
        RECT 2310.680 399.880 2310.940 400.140 ;
        RECT 2310.220 327.460 2310.480 327.720 ;
        RECT 2691.100 327.460 2691.360 327.720 ;
      LAYER met2 ;
        RECT 2310.810 510.410 2311.090 514.000 ;
        RECT 2310.280 510.270 2311.090 510.410 ;
        RECT 2310.280 483.325 2310.420 510.270 ;
        RECT 2310.810 510.000 2311.090 510.270 ;
        RECT 2310.210 482.955 2310.490 483.325 ;
        RECT 2311.130 482.955 2311.410 483.325 ;
        RECT 2311.200 448.790 2311.340 482.955 ;
        RECT 2310.220 448.530 2310.480 448.790 ;
        RECT 2310.220 448.470 2310.880 448.530 ;
        RECT 2311.140 448.470 2311.400 448.790 ;
        RECT 2310.280 448.390 2310.880 448.470 ;
        RECT 2310.740 400.850 2310.880 448.390 ;
        RECT 2310.680 400.530 2310.940 400.850 ;
        RECT 2310.680 399.850 2310.940 400.170 ;
        RECT 2310.740 351.970 2310.880 399.850 ;
        RECT 2310.280 351.830 2310.880 351.970 ;
        RECT 2310.280 327.750 2310.420 351.830 ;
        RECT 2310.220 327.430 2310.480 327.750 ;
        RECT 2691.100 327.430 2691.360 327.750 ;
        RECT 2691.160 17.410 2691.300 327.430 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 2310.210 483.000 2310.490 483.280 ;
        RECT 2311.130 483.000 2311.410 483.280 ;
      LAYER met3 ;
        RECT 2310.185 483.290 2310.515 483.305 ;
        RECT 2311.105 483.290 2311.435 483.305 ;
        RECT 2310.185 482.990 2311.435 483.290 ;
        RECT 2310.185 482.975 2310.515 482.990 ;
        RECT 2311.105 482.975 2311.435 482.990 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2326.750 498.680 2327.070 498.740 ;
        RECT 2331.810 498.680 2332.130 498.740 ;
        RECT 2326.750 498.540 2332.130 498.680 ;
        RECT 2326.750 498.480 2327.070 498.540 ;
        RECT 2331.810 498.480 2332.130 498.540 ;
        RECT 2331.810 334.460 2332.130 334.520 ;
        RECT 2711.770 334.460 2712.090 334.520 ;
        RECT 2331.810 334.320 2712.090 334.460 ;
        RECT 2331.810 334.260 2332.130 334.320 ;
        RECT 2711.770 334.260 2712.090 334.320 ;
      LAYER via ;
        RECT 2326.780 498.480 2327.040 498.740 ;
        RECT 2331.840 498.480 2332.100 498.740 ;
        RECT 2331.840 334.260 2332.100 334.520 ;
        RECT 2711.800 334.260 2712.060 334.520 ;
      LAYER met2 ;
        RECT 2326.910 510.340 2327.190 514.000 ;
        RECT 2326.840 510.000 2327.190 510.340 ;
        RECT 2326.840 498.770 2326.980 510.000 ;
        RECT 2326.780 498.450 2327.040 498.770 ;
        RECT 2331.840 498.450 2332.100 498.770 ;
        RECT 2331.900 334.550 2332.040 498.450 ;
        RECT 2331.840 334.230 2332.100 334.550 ;
        RECT 2711.800 334.230 2712.060 334.550 ;
        RECT 2711.860 17.410 2712.000 334.230 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 18.940 2345.930 19.000 ;
        RECT 2732.470 18.940 2732.790 19.000 ;
        RECT 2345.610 18.800 2732.790 18.940 ;
        RECT 2345.610 18.740 2345.930 18.800 ;
        RECT 2732.470 18.740 2732.790 18.800 ;
      LAYER via ;
        RECT 2345.640 18.740 2345.900 19.000 ;
        RECT 2732.500 18.740 2732.760 19.000 ;
      LAYER met2 ;
        RECT 2343.470 510.410 2343.750 514.000 ;
        RECT 2343.470 510.270 2345.840 510.410 ;
        RECT 2343.470 510.000 2343.750 510.270 ;
        RECT 2345.700 19.030 2345.840 510.270 ;
        RECT 2345.640 18.710 2345.900 19.030 ;
        RECT 2732.500 18.710 2732.760 19.030 ;
        RECT 2732.560 2.400 2732.700 18.710 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2359.410 20.640 2359.730 20.700 ;
        RECT 2750.410 20.640 2750.730 20.700 ;
        RECT 2359.410 20.500 2750.730 20.640 ;
        RECT 2359.410 20.440 2359.730 20.500 ;
        RECT 2750.410 20.440 2750.730 20.500 ;
      LAYER via ;
        RECT 2359.440 20.440 2359.700 20.700 ;
        RECT 2750.440 20.440 2750.700 20.700 ;
      LAYER met2 ;
        RECT 2359.570 510.340 2359.850 514.000 ;
        RECT 2359.500 510.000 2359.850 510.340 ;
        RECT 2359.500 20.730 2359.640 510.000 ;
        RECT 2359.440 20.410 2359.700 20.730 ;
        RECT 2750.440 20.410 2750.700 20.730 ;
        RECT 2750.500 2.400 2750.640 20.410 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2375.970 496.980 2376.290 497.040 ;
        RECT 2380.110 496.980 2380.430 497.040 ;
        RECT 2375.970 496.840 2380.430 496.980 ;
        RECT 2375.970 496.780 2376.290 496.840 ;
        RECT 2380.110 496.780 2380.430 496.840 ;
        RECT 2380.110 20.300 2380.430 20.360 ;
        RECT 2767.890 20.300 2768.210 20.360 ;
        RECT 2380.110 20.160 2768.210 20.300 ;
        RECT 2380.110 20.100 2380.430 20.160 ;
        RECT 2767.890 20.100 2768.210 20.160 ;
      LAYER via ;
        RECT 2376.000 496.780 2376.260 497.040 ;
        RECT 2380.140 496.780 2380.400 497.040 ;
        RECT 2380.140 20.100 2380.400 20.360 ;
        RECT 2767.920 20.100 2768.180 20.360 ;
      LAYER met2 ;
        RECT 2376.130 510.340 2376.410 514.000 ;
        RECT 2376.060 510.000 2376.410 510.340 ;
        RECT 2376.060 497.070 2376.200 510.000 ;
        RECT 2376.000 496.750 2376.260 497.070 ;
        RECT 2380.140 496.750 2380.400 497.070 ;
        RECT 2380.200 20.390 2380.340 496.750 ;
        RECT 2380.140 20.070 2380.400 20.390 ;
        RECT 2767.920 20.070 2768.180 20.390 ;
        RECT 2767.980 2.400 2768.120 20.070 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.250 210.700 613.570 210.760 ;
        RECT 834.970 210.700 835.290 210.760 ;
        RECT 613.250 210.560 835.290 210.700 ;
        RECT 613.250 210.500 613.570 210.560 ;
        RECT 834.970 210.500 835.290 210.560 ;
        RECT 834.970 17.580 835.290 17.640 ;
        RECT 840.950 17.580 841.270 17.640 ;
        RECT 834.970 17.440 841.270 17.580 ;
        RECT 834.970 17.380 835.290 17.440 ;
        RECT 840.950 17.380 841.270 17.440 ;
      LAYER via ;
        RECT 613.280 210.500 613.540 210.760 ;
        RECT 835.000 210.500 835.260 210.760 ;
        RECT 835.000 17.380 835.260 17.640 ;
        RECT 840.980 17.380 841.240 17.640 ;
      LAYER met2 ;
        RECT 613.410 510.340 613.690 514.000 ;
        RECT 613.340 510.000 613.690 510.340 ;
        RECT 613.340 210.790 613.480 510.000 ;
        RECT 613.280 210.470 613.540 210.790 ;
        RECT 835.000 210.470 835.260 210.790 ;
        RECT 835.060 17.670 835.200 210.470 ;
        RECT 835.000 17.350 835.260 17.670 ;
        RECT 840.980 17.350 841.240 17.670 ;
        RECT 841.040 2.400 841.180 17.350 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2393.910 19.960 2394.230 20.020 ;
        RECT 2785.830 19.960 2786.150 20.020 ;
        RECT 2393.910 19.820 2786.150 19.960 ;
        RECT 2393.910 19.760 2394.230 19.820 ;
        RECT 2785.830 19.760 2786.150 19.820 ;
      LAYER via ;
        RECT 2393.940 19.760 2394.200 20.020 ;
        RECT 2785.860 19.760 2786.120 20.020 ;
      LAYER met2 ;
        RECT 2392.230 510.410 2392.510 514.000 ;
        RECT 2392.230 510.270 2394.140 510.410 ;
        RECT 2392.230 510.000 2392.510 510.270 ;
        RECT 2394.000 20.050 2394.140 510.270 ;
        RECT 2393.940 19.730 2394.200 20.050 ;
        RECT 2785.860 19.730 2786.120 20.050 ;
        RECT 2785.920 2.400 2786.060 19.730 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2408.630 503.440 2408.950 503.500 ;
        RECT 2414.610 503.440 2414.930 503.500 ;
        RECT 2408.630 503.300 2414.930 503.440 ;
        RECT 2408.630 503.240 2408.950 503.300 ;
        RECT 2414.610 503.240 2414.930 503.300 ;
        RECT 2414.610 19.620 2414.930 19.680 ;
        RECT 2803.770 19.620 2804.090 19.680 ;
        RECT 2414.610 19.480 2804.090 19.620 ;
        RECT 2414.610 19.420 2414.930 19.480 ;
        RECT 2803.770 19.420 2804.090 19.480 ;
      LAYER via ;
        RECT 2408.660 503.240 2408.920 503.500 ;
        RECT 2414.640 503.240 2414.900 503.500 ;
        RECT 2414.640 19.420 2414.900 19.680 ;
        RECT 2803.800 19.420 2804.060 19.680 ;
      LAYER met2 ;
        RECT 2408.790 510.340 2409.070 514.000 ;
        RECT 2408.720 510.000 2409.070 510.340 ;
        RECT 2408.720 503.530 2408.860 510.000 ;
        RECT 2408.660 503.210 2408.920 503.530 ;
        RECT 2414.640 503.210 2414.900 503.530 ;
        RECT 2414.700 19.710 2414.840 503.210 ;
        RECT 2414.640 19.390 2414.900 19.710 ;
        RECT 2803.800 19.390 2804.060 19.710 ;
        RECT 2803.860 2.400 2804.000 19.390 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2428.410 19.280 2428.730 19.340 ;
        RECT 2821.710 19.280 2822.030 19.340 ;
        RECT 2428.410 19.140 2822.030 19.280 ;
        RECT 2428.410 19.080 2428.730 19.140 ;
        RECT 2821.710 19.080 2822.030 19.140 ;
      LAYER via ;
        RECT 2428.440 19.080 2428.700 19.340 ;
        RECT 2821.740 19.080 2822.000 19.340 ;
      LAYER met2 ;
        RECT 2424.890 510.410 2425.170 514.000 ;
        RECT 2424.890 510.270 2428.640 510.410 ;
        RECT 2424.890 510.000 2425.170 510.270 ;
        RECT 2428.500 19.370 2428.640 510.270 ;
        RECT 2428.440 19.050 2428.700 19.370 ;
        RECT 2821.740 19.050 2822.000 19.370 ;
        RECT 2821.800 2.400 2821.940 19.050 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2500.245 18.105 2501.795 18.275 ;
        RECT 2739.445 18.105 2739.615 18.955 ;
        RECT 2790.965 18.105 2791.135 18.955 ;
      LAYER mcon ;
        RECT 2739.445 18.785 2739.615 18.955 ;
        RECT 2501.625 18.105 2501.795 18.275 ;
        RECT 2790.965 18.785 2791.135 18.955 ;
      LAYER met1 ;
        RECT 2739.385 18.940 2739.675 18.985 ;
        RECT 2790.905 18.940 2791.195 18.985 ;
        RECT 2739.385 18.800 2791.195 18.940 ;
        RECT 2739.385 18.755 2739.675 18.800 ;
        RECT 2790.905 18.755 2791.195 18.800 ;
        RECT 2442.210 18.260 2442.530 18.320 ;
        RECT 2500.185 18.260 2500.475 18.305 ;
        RECT 2442.210 18.120 2500.475 18.260 ;
        RECT 2442.210 18.060 2442.530 18.120 ;
        RECT 2500.185 18.075 2500.475 18.120 ;
        RECT 2501.565 18.260 2501.855 18.305 ;
        RECT 2739.385 18.260 2739.675 18.305 ;
        RECT 2501.565 18.120 2739.675 18.260 ;
        RECT 2501.565 18.075 2501.855 18.120 ;
        RECT 2739.385 18.075 2739.675 18.120 ;
        RECT 2790.905 18.260 2791.195 18.305 ;
        RECT 2835.970 18.260 2836.290 18.320 ;
        RECT 2790.905 18.120 2836.290 18.260 ;
        RECT 2790.905 18.075 2791.195 18.120 ;
        RECT 2835.970 18.060 2836.290 18.120 ;
        RECT 2835.970 16.900 2836.290 16.960 ;
        RECT 2839.190 16.900 2839.510 16.960 ;
        RECT 2835.970 16.760 2839.510 16.900 ;
        RECT 2835.970 16.700 2836.290 16.760 ;
        RECT 2839.190 16.700 2839.510 16.760 ;
      LAYER via ;
        RECT 2442.240 18.060 2442.500 18.320 ;
        RECT 2836.000 18.060 2836.260 18.320 ;
        RECT 2836.000 16.700 2836.260 16.960 ;
        RECT 2839.220 16.700 2839.480 16.960 ;
      LAYER met2 ;
        RECT 2441.450 510.410 2441.730 514.000 ;
        RECT 2441.450 510.270 2442.440 510.410 ;
        RECT 2441.450 510.000 2441.730 510.270 ;
        RECT 2442.300 18.350 2442.440 510.270 ;
        RECT 2442.240 18.030 2442.500 18.350 ;
        RECT 2836.000 18.030 2836.260 18.350 ;
        RECT 2836.060 16.990 2836.200 18.030 ;
        RECT 2836.000 16.670 2836.260 16.990 ;
        RECT 2839.220 16.670 2839.480 16.990 ;
        RECT 2839.280 2.400 2839.420 16.670 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2457.390 496.980 2457.710 497.040 ;
        RECT 2462.910 496.980 2463.230 497.040 ;
        RECT 2457.390 496.840 2463.230 496.980 ;
        RECT 2457.390 496.780 2457.710 496.840 ;
        RECT 2462.910 496.780 2463.230 496.840 ;
        RECT 2462.910 18.600 2463.230 18.660 ;
        RECT 2462.910 18.460 2501.320 18.600 ;
        RECT 2462.910 18.400 2463.230 18.460 ;
        RECT 2501.180 17.920 2501.320 18.460 ;
        RECT 2857.130 17.920 2857.450 17.980 ;
        RECT 2501.180 17.780 2857.450 17.920 ;
        RECT 2857.130 17.720 2857.450 17.780 ;
      LAYER via ;
        RECT 2457.420 496.780 2457.680 497.040 ;
        RECT 2462.940 496.780 2463.200 497.040 ;
        RECT 2462.940 18.400 2463.200 18.660 ;
        RECT 2857.160 17.720 2857.420 17.980 ;
      LAYER met2 ;
        RECT 2457.550 510.340 2457.830 514.000 ;
        RECT 2457.480 510.000 2457.830 510.340 ;
        RECT 2457.480 497.070 2457.620 510.000 ;
        RECT 2457.420 496.750 2457.680 497.070 ;
        RECT 2462.940 496.750 2463.200 497.070 ;
        RECT 2463.000 18.690 2463.140 496.750 ;
        RECT 2462.940 18.370 2463.200 18.690 ;
        RECT 2857.160 17.690 2857.420 18.010 ;
        RECT 2857.220 2.400 2857.360 17.690 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2476.250 17.920 2476.570 17.980 ;
        RECT 2476.250 17.780 2478.320 17.920 ;
        RECT 2476.250 17.720 2476.570 17.780 ;
        RECT 2478.180 17.580 2478.320 17.780 ;
        RECT 2875.070 17.580 2875.390 17.640 ;
        RECT 2478.180 17.440 2875.390 17.580 ;
        RECT 2875.070 17.380 2875.390 17.440 ;
      LAYER via ;
        RECT 2476.280 17.720 2476.540 17.980 ;
        RECT 2875.100 17.380 2875.360 17.640 ;
      LAYER met2 ;
        RECT 2474.110 510.410 2474.390 514.000 ;
        RECT 2474.110 510.270 2476.940 510.410 ;
        RECT 2474.110 510.000 2474.390 510.270 ;
        RECT 2476.800 26.250 2476.940 510.270 ;
        RECT 2476.340 26.110 2476.940 26.250 ;
        RECT 2476.340 18.010 2476.480 26.110 ;
        RECT 2476.280 17.690 2476.540 18.010 ;
        RECT 2875.100 17.350 2875.360 17.670 ;
        RECT 2875.160 2.400 2875.300 17.350 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 17.240 2490.830 17.300 ;
        RECT 2893.010 17.240 2893.330 17.300 ;
        RECT 2490.510 17.100 2893.330 17.240 ;
        RECT 2490.510 17.040 2490.830 17.100 ;
        RECT 2893.010 17.040 2893.330 17.100 ;
      LAYER via ;
        RECT 2490.540 17.040 2490.800 17.300 ;
        RECT 2893.040 17.040 2893.300 17.300 ;
      LAYER met2 ;
        RECT 2490.210 510.340 2490.490 514.000 ;
        RECT 2490.140 510.000 2490.490 510.340 ;
        RECT 2490.140 497.490 2490.280 510.000 ;
        RECT 2490.140 497.350 2490.740 497.490 ;
        RECT 2490.600 17.330 2490.740 497.350 ;
        RECT 2490.540 17.010 2490.800 17.330 ;
        RECT 2893.040 17.010 2893.300 17.330 ;
        RECT 2893.100 2.400 2893.240 17.010 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2506.610 496.980 2506.930 497.040 ;
        RECT 2511.210 496.980 2511.530 497.040 ;
        RECT 2506.610 496.840 2511.530 496.980 ;
        RECT 2506.610 496.780 2506.930 496.840 ;
        RECT 2511.210 496.780 2511.530 496.840 ;
        RECT 2511.210 18.600 2511.530 18.660 ;
        RECT 2910.950 18.600 2911.270 18.660 ;
        RECT 2511.210 18.460 2911.270 18.600 ;
        RECT 2511.210 18.400 2511.530 18.460 ;
        RECT 2910.950 18.400 2911.270 18.460 ;
      LAYER via ;
        RECT 2506.640 496.780 2506.900 497.040 ;
        RECT 2511.240 496.780 2511.500 497.040 ;
        RECT 2511.240 18.400 2511.500 18.660 ;
        RECT 2910.980 18.400 2911.240 18.660 ;
      LAYER met2 ;
        RECT 2506.770 510.340 2507.050 514.000 ;
        RECT 2506.700 510.000 2507.050 510.340 ;
        RECT 2506.700 497.070 2506.840 510.000 ;
        RECT 2506.640 496.750 2506.900 497.070 ;
        RECT 2511.240 496.750 2511.500 497.070 ;
        RECT 2511.300 18.690 2511.440 496.750 ;
        RECT 2511.240 18.370 2511.500 18.690 ;
        RECT 2910.980 18.370 2911.240 18.690 ;
        RECT 2911.040 2.400 2911.180 18.370 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 629.810 496.980 630.130 497.040 ;
        RECT 634.410 496.980 634.730 497.040 ;
        RECT 629.810 496.840 634.730 496.980 ;
        RECT 629.810 496.780 630.130 496.840 ;
        RECT 634.410 496.780 634.730 496.840 ;
        RECT 634.410 217.160 634.730 217.220 ;
        RECT 855.670 217.160 855.990 217.220 ;
        RECT 634.410 217.020 855.990 217.160 ;
        RECT 634.410 216.960 634.730 217.020 ;
        RECT 855.670 216.960 855.990 217.020 ;
      LAYER via ;
        RECT 629.840 496.780 630.100 497.040 ;
        RECT 634.440 496.780 634.700 497.040 ;
        RECT 634.440 216.960 634.700 217.220 ;
        RECT 855.700 216.960 855.960 217.220 ;
      LAYER met2 ;
        RECT 629.970 510.340 630.250 514.000 ;
        RECT 629.900 510.000 630.250 510.340 ;
        RECT 629.900 497.070 630.040 510.000 ;
        RECT 629.840 496.750 630.100 497.070 ;
        RECT 634.440 496.750 634.700 497.070 ;
        RECT 634.500 217.250 634.640 496.750 ;
        RECT 634.440 216.930 634.700 217.250 ;
        RECT 855.700 216.930 855.960 217.250 ;
        RECT 855.760 17.410 855.900 216.930 ;
        RECT 855.760 17.270 859.120 17.410 ;
        RECT 858.980 2.400 859.120 17.270 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 231.100 648.530 231.160 ;
        RECT 876.370 231.100 876.690 231.160 ;
        RECT 648.210 230.960 876.690 231.100 ;
        RECT 648.210 230.900 648.530 230.960 ;
        RECT 876.370 230.900 876.690 230.960 ;
      LAYER via ;
        RECT 648.240 230.900 648.500 231.160 ;
        RECT 876.400 230.900 876.660 231.160 ;
      LAYER met2 ;
        RECT 646.070 510.410 646.350 514.000 ;
        RECT 646.070 510.270 648.440 510.410 ;
        RECT 646.070 510.000 646.350 510.270 ;
        RECT 648.300 231.190 648.440 510.270 ;
        RECT 648.240 230.870 648.500 231.190 ;
        RECT 876.400 230.870 876.660 231.190 ;
        RECT 876.460 17.410 876.600 230.870 ;
        RECT 876.460 17.270 877.060 17.410 ;
        RECT 876.920 2.400 877.060 17.270 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.470 496.980 662.790 497.040 ;
        RECT 668.450 496.980 668.770 497.040 ;
        RECT 662.470 496.840 668.770 496.980 ;
        RECT 662.470 496.780 662.790 496.840 ;
        RECT 668.450 496.780 668.770 496.840 ;
        RECT 668.450 245.380 668.770 245.440 ;
        RECT 890.170 245.380 890.490 245.440 ;
        RECT 668.450 245.240 890.490 245.380 ;
        RECT 668.450 245.180 668.770 245.240 ;
        RECT 890.170 245.180 890.490 245.240 ;
      LAYER via ;
        RECT 662.500 496.780 662.760 497.040 ;
        RECT 668.480 496.780 668.740 497.040 ;
        RECT 668.480 245.180 668.740 245.440 ;
        RECT 890.200 245.180 890.460 245.440 ;
      LAYER met2 ;
        RECT 662.630 510.340 662.910 514.000 ;
        RECT 662.560 510.000 662.910 510.340 ;
        RECT 662.560 497.070 662.700 510.000 ;
        RECT 662.500 496.750 662.760 497.070 ;
        RECT 668.480 496.750 668.740 497.070 ;
        RECT 668.540 245.470 668.680 496.750 ;
        RECT 668.480 245.150 668.740 245.470 ;
        RECT 890.200 245.150 890.460 245.470 ;
        RECT 890.260 17.410 890.400 245.150 ;
        RECT 890.260 17.270 895.000 17.410 ;
        RECT 894.860 2.400 895.000 17.270 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 678.570 496.980 678.890 497.040 ;
        RECT 682.710 496.980 683.030 497.040 ;
        RECT 678.570 496.840 683.030 496.980 ;
        RECT 678.570 496.780 678.890 496.840 ;
        RECT 682.710 496.780 683.030 496.840 ;
        RECT 682.710 251.840 683.030 251.900 ;
        RECT 910.870 251.840 911.190 251.900 ;
        RECT 682.710 251.700 911.190 251.840 ;
        RECT 682.710 251.640 683.030 251.700 ;
        RECT 910.870 251.640 911.190 251.700 ;
      LAYER via ;
        RECT 678.600 496.780 678.860 497.040 ;
        RECT 682.740 496.780 683.000 497.040 ;
        RECT 682.740 251.640 683.000 251.900 ;
        RECT 910.900 251.640 911.160 251.900 ;
      LAYER met2 ;
        RECT 678.730 510.340 679.010 514.000 ;
        RECT 678.660 510.000 679.010 510.340 ;
        RECT 678.660 497.070 678.800 510.000 ;
        RECT 678.600 496.750 678.860 497.070 ;
        RECT 682.740 496.750 683.000 497.070 ;
        RECT 682.800 251.930 682.940 496.750 ;
        RECT 682.740 251.610 683.000 251.930 ;
        RECT 910.900 251.610 911.160 251.930 ;
        RECT 910.960 17.410 911.100 251.610 ;
        RECT 910.960 17.270 912.940 17.410 ;
        RECT 912.800 2.400 912.940 17.270 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.510 258.640 696.830 258.700 ;
        RECT 924.670 258.640 924.990 258.700 ;
        RECT 696.510 258.500 924.990 258.640 ;
        RECT 696.510 258.440 696.830 258.500 ;
        RECT 924.670 258.440 924.990 258.500 ;
      LAYER via ;
        RECT 696.540 258.440 696.800 258.700 ;
        RECT 924.700 258.440 924.960 258.700 ;
      LAYER met2 ;
        RECT 694.830 510.410 695.110 514.000 ;
        RECT 694.830 510.270 696.740 510.410 ;
        RECT 694.830 510.000 695.110 510.270 ;
        RECT 696.600 258.730 696.740 510.270 ;
        RECT 696.540 258.410 696.800 258.730 ;
        RECT 924.700 258.410 924.960 258.730 ;
        RECT 924.760 17.410 924.900 258.410 ;
        RECT 924.760 17.270 930.420 17.410 ;
        RECT 930.280 2.400 930.420 17.270 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.230 496.980 711.550 497.040 ;
        RECT 716.750 496.980 717.070 497.040 ;
        RECT 711.230 496.840 717.070 496.980 ;
        RECT 711.230 496.780 711.550 496.840 ;
        RECT 716.750 496.780 717.070 496.840 ;
        RECT 716.750 265.440 717.070 265.500 ;
        RECT 945.370 265.440 945.690 265.500 ;
        RECT 716.750 265.300 945.690 265.440 ;
        RECT 716.750 265.240 717.070 265.300 ;
        RECT 945.370 265.240 945.690 265.300 ;
      LAYER via ;
        RECT 711.260 496.780 711.520 497.040 ;
        RECT 716.780 496.780 717.040 497.040 ;
        RECT 716.780 265.240 717.040 265.500 ;
        RECT 945.400 265.240 945.660 265.500 ;
      LAYER met2 ;
        RECT 711.390 510.340 711.670 514.000 ;
        RECT 711.320 510.000 711.670 510.340 ;
        RECT 711.320 497.070 711.460 510.000 ;
        RECT 711.260 496.750 711.520 497.070 ;
        RECT 716.780 496.750 717.040 497.070 ;
        RECT 716.840 265.530 716.980 496.750 ;
        RECT 716.780 265.210 717.040 265.530 ;
        RECT 945.400 265.210 945.660 265.530 ;
        RECT 945.460 17.410 945.600 265.210 ;
        RECT 945.460 17.270 948.360 17.410 ;
        RECT 948.220 2.400 948.360 17.270 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 731.010 272.580 731.330 272.640 ;
        RECT 966.070 272.580 966.390 272.640 ;
        RECT 731.010 272.440 966.390 272.580 ;
        RECT 731.010 272.380 731.330 272.440 ;
        RECT 966.070 272.380 966.390 272.440 ;
      LAYER via ;
        RECT 731.040 272.380 731.300 272.640 ;
        RECT 966.100 272.380 966.360 272.640 ;
      LAYER met2 ;
        RECT 727.490 510.410 727.770 514.000 ;
        RECT 727.490 510.270 731.240 510.410 ;
        RECT 727.490 510.000 727.770 510.270 ;
        RECT 731.100 272.670 731.240 510.270 ;
        RECT 731.040 272.350 731.300 272.670 ;
        RECT 966.100 272.350 966.360 272.670 ;
        RECT 966.160 2.400 966.300 272.350 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 744.425 338.045 744.595 386.155 ;
      LAYER mcon ;
        RECT 744.425 385.985 744.595 386.155 ;
      LAYER met1 ;
        RECT 743.430 448.700 743.750 448.760 ;
        RECT 744.350 448.700 744.670 448.760 ;
        RECT 743.430 448.560 744.670 448.700 ;
        RECT 743.430 448.500 743.750 448.560 ;
        RECT 744.350 448.500 744.670 448.560 ;
        RECT 744.365 386.140 744.655 386.185 ;
        RECT 744.810 386.140 745.130 386.200 ;
        RECT 744.365 386.000 745.130 386.140 ;
        RECT 744.365 385.955 744.655 386.000 ;
        RECT 744.810 385.940 745.130 386.000 ;
        RECT 744.350 338.200 744.670 338.260 ;
        RECT 744.155 338.060 744.670 338.200 ;
        RECT 744.350 338.000 744.670 338.060 ;
        RECT 744.350 304.200 744.670 304.260 ;
        RECT 743.980 304.060 744.670 304.200 ;
        RECT 743.980 303.580 744.120 304.060 ;
        RECT 744.350 304.000 744.670 304.060 ;
        RECT 743.890 303.320 744.210 303.580 ;
        RECT 743.890 279.380 744.210 279.440 ;
        RECT 979.870 279.380 980.190 279.440 ;
        RECT 743.890 279.240 980.190 279.380 ;
        RECT 743.890 279.180 744.210 279.240 ;
        RECT 979.870 279.180 980.190 279.240 ;
      LAYER via ;
        RECT 743.460 448.500 743.720 448.760 ;
        RECT 744.380 448.500 744.640 448.760 ;
        RECT 744.840 385.940 745.100 386.200 ;
        RECT 744.380 338.000 744.640 338.260 ;
        RECT 744.380 304.000 744.640 304.260 ;
        RECT 743.920 303.320 744.180 303.580 ;
        RECT 743.920 279.180 744.180 279.440 ;
        RECT 979.900 279.180 980.160 279.440 ;
      LAYER met2 ;
        RECT 744.050 511.090 744.330 514.000 ;
        RECT 744.050 510.950 745.040 511.090 ;
        RECT 744.050 510.000 744.330 510.950 ;
        RECT 744.900 483.210 745.040 510.950 ;
        RECT 744.440 483.070 745.040 483.210 ;
        RECT 744.440 448.790 744.580 483.070 ;
        RECT 743.460 448.530 743.720 448.790 ;
        RECT 744.380 448.530 744.640 448.790 ;
        RECT 743.460 448.470 744.640 448.530 ;
        RECT 743.520 448.390 744.580 448.470 ;
        RECT 744.440 386.650 744.580 448.390 ;
        RECT 744.440 386.510 745.040 386.650 ;
        RECT 744.900 386.230 745.040 386.510 ;
        RECT 744.840 385.910 745.100 386.230 ;
        RECT 744.380 337.970 744.640 338.290 ;
        RECT 744.440 304.290 744.580 337.970 ;
        RECT 744.380 303.970 744.640 304.290 ;
        RECT 743.920 303.290 744.180 303.610 ;
        RECT 743.980 279.470 744.120 303.290 ;
        RECT 743.920 279.150 744.180 279.470 ;
        RECT 979.900 279.150 980.160 279.470 ;
        RECT 979.960 17.410 980.100 279.150 ;
        RECT 979.960 17.270 984.240 17.410 ;
        RECT 984.100 2.400 984.240 17.270 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 449.950 498.000 450.270 498.060 ;
        RECT 455.010 498.000 455.330 498.060 ;
        RECT 449.950 497.860 455.330 498.000 ;
        RECT 449.950 497.800 450.270 497.860 ;
        RECT 455.010 497.800 455.330 497.860 ;
        RECT 455.010 19.960 455.330 20.020 ;
        RECT 662.470 19.960 662.790 20.020 ;
        RECT 455.010 19.820 662.790 19.960 ;
        RECT 455.010 19.760 455.330 19.820 ;
        RECT 662.470 19.760 662.790 19.820 ;
      LAYER via ;
        RECT 449.980 497.800 450.240 498.060 ;
        RECT 455.040 497.800 455.300 498.060 ;
        RECT 455.040 19.760 455.300 20.020 ;
        RECT 662.500 19.760 662.760 20.020 ;
      LAYER met2 ;
        RECT 450.110 510.340 450.390 514.000 ;
        RECT 450.040 510.000 450.390 510.340 ;
        RECT 450.040 498.090 450.180 510.000 ;
        RECT 449.980 497.770 450.240 498.090 ;
        RECT 455.040 497.770 455.300 498.090 ;
        RECT 455.100 20.050 455.240 497.770 ;
        RECT 455.040 19.730 455.300 20.050 ;
        RECT 662.500 19.730 662.760 20.050 ;
        RECT 662.560 16.050 662.700 19.730 ;
        RECT 662.560 15.910 663.160 16.050 ;
        RECT 663.020 2.400 663.160 15.910 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 764.205 386.325 764.375 434.775 ;
      LAYER mcon ;
        RECT 764.205 434.605 764.375 434.775 ;
      LAYER met1 ;
        RECT 759.990 496.980 760.310 497.040 ;
        RECT 759.990 496.840 765.280 496.980 ;
        RECT 759.990 496.780 760.310 496.840 ;
        RECT 765.140 496.700 765.280 496.840 ;
        RECT 765.050 496.440 765.370 496.700 ;
        RECT 764.145 434.760 764.435 434.805 ;
        RECT 764.590 434.760 764.910 434.820 ;
        RECT 764.145 434.620 764.910 434.760 ;
        RECT 764.145 434.575 764.435 434.620 ;
        RECT 764.590 434.560 764.910 434.620 ;
        RECT 764.130 386.480 764.450 386.540 ;
        RECT 763.935 386.340 764.450 386.480 ;
        RECT 764.130 386.280 764.450 386.340 ;
        RECT 765.050 352.140 765.370 352.200 ;
        RECT 764.680 352.000 765.370 352.140 ;
        RECT 764.680 351.520 764.820 352.000 ;
        RECT 765.050 351.940 765.370 352.000 ;
        RECT 764.590 351.260 764.910 351.520 ;
        RECT 764.590 286.180 764.910 286.240 ;
        RECT 1000.570 286.180 1000.890 286.240 ;
        RECT 764.590 286.040 1000.890 286.180 ;
        RECT 764.590 285.980 764.910 286.040 ;
        RECT 1000.570 285.980 1000.890 286.040 ;
      LAYER via ;
        RECT 760.020 496.780 760.280 497.040 ;
        RECT 765.080 496.440 765.340 496.700 ;
        RECT 764.620 434.560 764.880 434.820 ;
        RECT 764.160 386.280 764.420 386.540 ;
        RECT 765.080 351.940 765.340 352.200 ;
        RECT 764.620 351.260 764.880 351.520 ;
        RECT 764.620 285.980 764.880 286.240 ;
        RECT 1000.600 285.980 1000.860 286.240 ;
      LAYER met2 ;
        RECT 760.150 510.340 760.430 514.000 ;
        RECT 760.080 510.000 760.430 510.340 ;
        RECT 760.080 497.070 760.220 510.000 ;
        RECT 760.020 496.750 760.280 497.070 ;
        RECT 765.080 496.410 765.340 496.730 ;
        RECT 765.140 448.530 765.280 496.410 ;
        RECT 764.680 448.390 765.280 448.530 ;
        RECT 764.680 434.850 764.820 448.390 ;
        RECT 764.620 434.530 764.880 434.850 ;
        RECT 764.160 386.250 764.420 386.570 ;
        RECT 764.220 386.085 764.360 386.250 ;
        RECT 764.150 385.715 764.430 386.085 ;
        RECT 765.070 385.715 765.350 386.085 ;
        RECT 765.140 352.230 765.280 385.715 ;
        RECT 765.080 351.910 765.340 352.230 ;
        RECT 764.620 351.230 764.880 351.550 ;
        RECT 764.680 286.270 764.820 351.230 ;
        RECT 764.620 285.950 764.880 286.270 ;
        RECT 1000.600 285.950 1000.860 286.270 ;
        RECT 1000.660 17.410 1000.800 285.950 ;
        RECT 1000.660 17.270 1002.180 17.410 ;
        RECT 1002.040 2.400 1002.180 17.270 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
      LAYER via2 ;
        RECT 764.150 385.760 764.430 386.040 ;
        RECT 765.070 385.760 765.350 386.040 ;
      LAYER met3 ;
        RECT 764.125 386.050 764.455 386.065 ;
        RECT 765.045 386.050 765.375 386.065 ;
        RECT 764.125 385.750 765.375 386.050 ;
        RECT 764.125 385.735 764.455 385.750 ;
        RECT 765.045 385.735 765.375 385.750 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 293.320 779.630 293.380 ;
        RECT 1014.370 293.320 1014.690 293.380 ;
        RECT 779.310 293.180 1014.690 293.320 ;
        RECT 779.310 293.120 779.630 293.180 ;
        RECT 1014.370 293.120 1014.690 293.180 ;
      LAYER via ;
        RECT 779.340 293.120 779.600 293.380 ;
        RECT 1014.400 293.120 1014.660 293.380 ;
      LAYER met2 ;
        RECT 776.710 510.410 776.990 514.000 ;
        RECT 776.710 510.270 779.540 510.410 ;
        RECT 776.710 510.000 776.990 510.270 ;
        RECT 779.400 293.410 779.540 510.270 ;
        RECT 779.340 293.090 779.600 293.410 ;
        RECT 1014.400 293.090 1014.660 293.410 ;
        RECT 1014.460 17.410 1014.600 293.090 ;
        RECT 1014.460 17.270 1019.660 17.410 ;
        RECT 1019.520 2.400 1019.660 17.270 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 792.650 306.920 792.970 306.980 ;
        RECT 1035.070 306.920 1035.390 306.980 ;
        RECT 792.650 306.780 1035.390 306.920 ;
        RECT 792.650 306.720 792.970 306.780 ;
        RECT 1035.070 306.720 1035.390 306.780 ;
      LAYER via ;
        RECT 792.680 306.720 792.940 306.980 ;
        RECT 1035.100 306.720 1035.360 306.980 ;
      LAYER met2 ;
        RECT 792.810 510.340 793.090 514.000 ;
        RECT 792.740 510.000 793.090 510.340 ;
        RECT 792.740 307.010 792.880 510.000 ;
        RECT 792.680 306.690 792.940 307.010 ;
        RECT 1035.100 306.690 1035.360 307.010 ;
        RECT 1035.160 17.410 1035.300 306.690 ;
        RECT 1035.160 17.270 1037.600 17.410 ;
        RECT 1037.460 2.400 1037.600 17.270 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 809.210 496.980 809.530 497.040 ;
        RECT 813.810 496.980 814.130 497.040 ;
        RECT 809.210 496.840 814.130 496.980 ;
        RECT 809.210 496.780 809.530 496.840 ;
        RECT 813.810 496.780 814.130 496.840 ;
        RECT 813.810 196.760 814.130 196.820 ;
        RECT 1048.870 196.760 1049.190 196.820 ;
        RECT 813.810 196.620 1049.190 196.760 ;
        RECT 813.810 196.560 814.130 196.620 ;
        RECT 1048.870 196.560 1049.190 196.620 ;
        RECT 1048.870 17.580 1049.190 17.640 ;
        RECT 1055.310 17.580 1055.630 17.640 ;
        RECT 1048.870 17.440 1055.630 17.580 ;
        RECT 1048.870 17.380 1049.190 17.440 ;
        RECT 1055.310 17.380 1055.630 17.440 ;
      LAYER via ;
        RECT 809.240 496.780 809.500 497.040 ;
        RECT 813.840 496.780 814.100 497.040 ;
        RECT 813.840 196.560 814.100 196.820 ;
        RECT 1048.900 196.560 1049.160 196.820 ;
        RECT 1048.900 17.380 1049.160 17.640 ;
        RECT 1055.340 17.380 1055.600 17.640 ;
      LAYER met2 ;
        RECT 809.370 510.340 809.650 514.000 ;
        RECT 809.300 510.000 809.650 510.340 ;
        RECT 809.300 497.070 809.440 510.000 ;
        RECT 809.240 496.750 809.500 497.070 ;
        RECT 813.840 496.750 814.100 497.070 ;
        RECT 813.900 196.850 814.040 496.750 ;
        RECT 813.840 196.530 814.100 196.850 ;
        RECT 1048.900 196.530 1049.160 196.850 ;
        RECT 1048.960 17.670 1049.100 196.530 ;
        RECT 1048.900 17.350 1049.160 17.670 ;
        RECT 1055.340 17.350 1055.600 17.670 ;
        RECT 1055.400 2.400 1055.540 17.350 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 210.360 827.930 210.420 ;
        RECT 1069.570 210.360 1069.890 210.420 ;
        RECT 827.610 210.220 1069.890 210.360 ;
        RECT 827.610 210.160 827.930 210.220 ;
        RECT 1069.570 210.160 1069.890 210.220 ;
      LAYER via ;
        RECT 827.640 210.160 827.900 210.420 ;
        RECT 1069.600 210.160 1069.860 210.420 ;
      LAYER met2 ;
        RECT 825.470 510.410 825.750 514.000 ;
        RECT 825.470 510.270 827.840 510.410 ;
        RECT 825.470 510.000 825.750 510.270 ;
        RECT 827.700 210.450 827.840 510.270 ;
        RECT 827.640 210.130 827.900 210.450 ;
        RECT 1069.600 210.130 1069.860 210.450 ;
        RECT 1069.660 17.410 1069.800 210.130 ;
        RECT 1069.660 17.270 1073.480 17.410 ;
        RECT 1073.340 2.400 1073.480 17.270 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.870 496.980 842.190 497.040 ;
        RECT 847.850 496.980 848.170 497.040 ;
        RECT 841.870 496.840 848.170 496.980 ;
        RECT 841.870 496.780 842.190 496.840 ;
        RECT 847.850 496.780 848.170 496.840 ;
        RECT 847.850 300.120 848.170 300.180 ;
        RECT 1090.270 300.120 1090.590 300.180 ;
        RECT 847.850 299.980 1090.590 300.120 ;
        RECT 847.850 299.920 848.170 299.980 ;
        RECT 1090.270 299.920 1090.590 299.980 ;
      LAYER via ;
        RECT 841.900 496.780 842.160 497.040 ;
        RECT 847.880 496.780 848.140 497.040 ;
        RECT 847.880 299.920 848.140 300.180 ;
        RECT 1090.300 299.920 1090.560 300.180 ;
      LAYER met2 ;
        RECT 842.030 510.340 842.310 514.000 ;
        RECT 841.960 510.000 842.310 510.340 ;
        RECT 841.960 497.070 842.100 510.000 ;
        RECT 841.900 496.750 842.160 497.070 ;
        RECT 847.880 496.750 848.140 497.070 ;
        RECT 847.940 300.210 848.080 496.750 ;
        RECT 847.880 299.890 848.140 300.210 ;
        RECT 1090.300 299.890 1090.560 300.210 ;
        RECT 1090.360 17.410 1090.500 299.890 ;
        RECT 1090.360 17.270 1090.960 17.410 ;
        RECT 1090.820 2.400 1090.960 17.270 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 857.970 496.980 858.290 497.040 ;
        RECT 862.110 496.980 862.430 497.040 ;
        RECT 857.970 496.840 862.430 496.980 ;
        RECT 857.970 496.780 858.290 496.840 ;
        RECT 862.110 496.780 862.430 496.840 ;
        RECT 862.110 314.060 862.430 314.120 ;
        RECT 1104.070 314.060 1104.390 314.120 ;
        RECT 862.110 313.920 1104.390 314.060 ;
        RECT 862.110 313.860 862.430 313.920 ;
        RECT 1104.070 313.860 1104.390 313.920 ;
      LAYER via ;
        RECT 858.000 496.780 858.260 497.040 ;
        RECT 862.140 496.780 862.400 497.040 ;
        RECT 862.140 313.860 862.400 314.120 ;
        RECT 1104.100 313.860 1104.360 314.120 ;
      LAYER met2 ;
        RECT 858.130 510.340 858.410 514.000 ;
        RECT 858.060 510.000 858.410 510.340 ;
        RECT 858.060 497.070 858.200 510.000 ;
        RECT 858.000 496.750 858.260 497.070 ;
        RECT 862.140 496.750 862.400 497.070 ;
        RECT 862.200 314.150 862.340 496.750 ;
        RECT 862.140 313.830 862.400 314.150 ;
        RECT 1104.100 313.830 1104.360 314.150 ;
        RECT 1104.160 17.410 1104.300 313.830 ;
        RECT 1104.160 17.270 1108.900 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 875.910 245.040 876.230 245.100 ;
        RECT 1124.770 245.040 1125.090 245.100 ;
        RECT 875.910 244.900 1125.090 245.040 ;
        RECT 875.910 244.840 876.230 244.900 ;
        RECT 1124.770 244.840 1125.090 244.900 ;
      LAYER via ;
        RECT 875.940 244.840 876.200 245.100 ;
        RECT 1124.800 244.840 1125.060 245.100 ;
      LAYER met2 ;
        RECT 874.690 510.410 874.970 514.000 ;
        RECT 874.690 510.270 876.140 510.410 ;
        RECT 874.690 510.000 874.970 510.270 ;
        RECT 876.000 245.130 876.140 510.270 ;
        RECT 875.940 244.810 876.200 245.130 ;
        RECT 1124.800 244.810 1125.060 245.130 ;
        RECT 1124.860 17.410 1125.000 244.810 ;
        RECT 1124.860 17.270 1126.840 17.410 ;
        RECT 1126.700 2.400 1126.840 17.270 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.630 496.980 890.950 497.040 ;
        RECT 896.150 496.980 896.470 497.040 ;
        RECT 890.630 496.840 896.470 496.980 ;
        RECT 890.630 496.780 890.950 496.840 ;
        RECT 896.150 496.780 896.470 496.840 ;
        RECT 896.150 321.200 896.470 321.260 ;
        RECT 1138.570 321.200 1138.890 321.260 ;
        RECT 896.150 321.060 1138.890 321.200 ;
        RECT 896.150 321.000 896.470 321.060 ;
        RECT 1138.570 321.000 1138.890 321.060 ;
        RECT 1138.570 17.920 1138.890 17.980 ;
        RECT 1144.550 17.920 1144.870 17.980 ;
        RECT 1138.570 17.780 1144.870 17.920 ;
        RECT 1138.570 17.720 1138.890 17.780 ;
        RECT 1144.550 17.720 1144.870 17.780 ;
      LAYER via ;
        RECT 890.660 496.780 890.920 497.040 ;
        RECT 896.180 496.780 896.440 497.040 ;
        RECT 896.180 321.000 896.440 321.260 ;
        RECT 1138.600 321.000 1138.860 321.260 ;
        RECT 1138.600 17.720 1138.860 17.980 ;
        RECT 1144.580 17.720 1144.840 17.980 ;
      LAYER met2 ;
        RECT 890.790 510.340 891.070 514.000 ;
        RECT 890.720 510.000 891.070 510.340 ;
        RECT 890.720 497.070 890.860 510.000 ;
        RECT 890.660 496.750 890.920 497.070 ;
        RECT 896.180 496.750 896.440 497.070 ;
        RECT 896.240 321.290 896.380 496.750 ;
        RECT 896.180 320.970 896.440 321.290 ;
        RECT 1138.600 320.970 1138.860 321.290 ;
        RECT 1138.660 18.010 1138.800 320.970 ;
        RECT 1138.600 17.690 1138.860 18.010 ;
        RECT 1144.580 17.690 1144.840 18.010 ;
        RECT 1144.640 2.400 1144.780 17.690 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 910.410 327.660 910.730 327.720 ;
        RECT 1159.270 327.660 1159.590 327.720 ;
        RECT 910.410 327.520 1159.590 327.660 ;
        RECT 910.410 327.460 910.730 327.520 ;
        RECT 1159.270 327.460 1159.590 327.520 ;
      LAYER via ;
        RECT 910.440 327.460 910.700 327.720 ;
        RECT 1159.300 327.460 1159.560 327.720 ;
      LAYER met2 ;
        RECT 907.350 510.410 907.630 514.000 ;
        RECT 907.350 510.270 910.640 510.410 ;
        RECT 907.350 510.000 907.630 510.270 ;
        RECT 910.500 327.750 910.640 510.270 ;
        RECT 910.440 327.430 910.700 327.750 ;
        RECT 1159.300 327.430 1159.560 327.750 ;
        RECT 1159.360 17.410 1159.500 327.430 ;
        RECT 1159.360 17.270 1162.720 17.410 ;
        RECT 1162.580 2.400 1162.720 17.270 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 468.810 19.620 469.130 19.680 ;
        RECT 680.410 19.620 680.730 19.680 ;
        RECT 468.810 19.480 680.730 19.620 ;
        RECT 468.810 19.420 469.130 19.480 ;
        RECT 680.410 19.420 680.730 19.480 ;
      LAYER via ;
        RECT 468.840 19.420 469.100 19.680 ;
        RECT 680.440 19.420 680.700 19.680 ;
      LAYER met2 ;
        RECT 466.670 510.410 466.950 514.000 ;
        RECT 466.670 510.270 469.040 510.410 ;
        RECT 466.670 510.000 466.950 510.270 ;
        RECT 468.900 19.710 469.040 510.270 ;
        RECT 468.840 19.390 469.100 19.710 ;
        RECT 680.440 19.390 680.700 19.710 ;
        RECT 680.500 2.400 680.640 19.390 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 924.210 334.460 924.530 334.520 ;
        RECT 1179.970 334.460 1180.290 334.520 ;
        RECT 924.210 334.320 1180.290 334.460 ;
        RECT 924.210 334.260 924.530 334.320 ;
        RECT 1179.970 334.260 1180.290 334.320 ;
      LAYER via ;
        RECT 924.240 334.260 924.500 334.520 ;
        RECT 1180.000 334.260 1180.260 334.520 ;
      LAYER met2 ;
        RECT 923.450 510.410 923.730 514.000 ;
        RECT 923.450 510.270 924.440 510.410 ;
        RECT 923.450 510.000 923.730 510.270 ;
        RECT 924.300 334.550 924.440 510.270 ;
        RECT 924.240 334.230 924.500 334.550 ;
        RECT 1180.000 334.230 1180.260 334.550 ;
        RECT 1180.060 2.400 1180.200 334.230 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 942.685 338.045 942.855 386.155 ;
      LAYER mcon ;
        RECT 942.685 385.985 942.855 386.155 ;
      LAYER met1 ;
        RECT 939.850 496.980 940.170 497.040 ;
        RECT 939.850 496.840 944.680 496.980 ;
        RECT 939.850 496.780 940.170 496.840 ;
        RECT 944.540 496.300 944.680 496.840 ;
        RECT 944.910 496.300 945.230 496.360 ;
        RECT 944.540 496.160 945.230 496.300 ;
        RECT 944.910 496.100 945.230 496.160 ;
        RECT 943.530 410.620 943.850 410.680 ;
        RECT 944.450 410.620 944.770 410.680 ;
        RECT 943.530 410.480 944.770 410.620 ;
        RECT 943.530 410.420 943.850 410.480 ;
        RECT 944.450 410.420 944.770 410.480 ;
        RECT 942.625 386.140 942.915 386.185 ;
        RECT 943.070 386.140 943.390 386.200 ;
        RECT 942.625 386.000 943.390 386.140 ;
        RECT 942.625 385.955 942.915 386.000 ;
        RECT 943.070 385.940 943.390 386.000 ;
        RECT 942.610 338.200 942.930 338.260 ;
        RECT 942.415 338.060 942.930 338.200 ;
        RECT 942.610 338.000 942.930 338.060 ;
        RECT 943.530 258.640 943.850 258.700 ;
        RECT 1193.770 258.640 1194.090 258.700 ;
        RECT 943.530 258.500 1194.090 258.640 ;
        RECT 943.530 258.440 943.850 258.500 ;
        RECT 1193.770 258.440 1194.090 258.500 ;
      LAYER via ;
        RECT 939.880 496.780 940.140 497.040 ;
        RECT 944.940 496.100 945.200 496.360 ;
        RECT 943.560 410.420 943.820 410.680 ;
        RECT 944.480 410.420 944.740 410.680 ;
        RECT 943.100 385.940 943.360 386.200 ;
        RECT 942.640 338.000 942.900 338.260 ;
        RECT 943.560 258.440 943.820 258.700 ;
        RECT 1193.800 258.440 1194.060 258.700 ;
      LAYER met2 ;
        RECT 940.010 510.340 940.290 514.000 ;
        RECT 939.940 510.000 940.290 510.340 ;
        RECT 939.940 497.070 940.080 510.000 ;
        RECT 939.880 496.750 940.140 497.070 ;
        RECT 944.940 496.070 945.200 496.390 ;
        RECT 945.000 468.930 945.140 496.070 ;
        RECT 944.540 468.790 945.140 468.930 ;
        RECT 944.540 448.530 944.680 468.790 ;
        RECT 943.620 448.390 944.680 448.530 ;
        RECT 943.620 410.710 943.760 448.390 ;
        RECT 943.560 410.390 943.820 410.710 ;
        RECT 944.480 410.390 944.740 410.710 ;
        RECT 944.540 386.765 944.680 410.390 ;
        RECT 943.550 386.650 943.830 386.765 ;
        RECT 943.160 386.510 943.830 386.650 ;
        RECT 943.160 386.230 943.300 386.510 ;
        RECT 943.550 386.395 943.830 386.510 ;
        RECT 944.470 386.395 944.750 386.765 ;
        RECT 943.100 385.910 943.360 386.230 ;
        RECT 942.640 337.970 942.900 338.290 ;
        RECT 942.700 303.690 942.840 337.970 ;
        RECT 942.700 303.550 943.760 303.690 ;
        RECT 943.620 258.730 943.760 303.550 ;
        RECT 943.560 258.410 943.820 258.730 ;
        RECT 1193.800 258.410 1194.060 258.730 ;
        RECT 1193.860 17.410 1194.000 258.410 ;
        RECT 1193.860 17.270 1198.140 17.410 ;
        RECT 1198.000 2.400 1198.140 17.270 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 943.550 386.440 943.830 386.720 ;
        RECT 944.470 386.440 944.750 386.720 ;
      LAYER met3 ;
        RECT 943.525 386.730 943.855 386.745 ;
        RECT 944.445 386.730 944.775 386.745 ;
        RECT 943.525 386.430 944.775 386.730 ;
        RECT 943.525 386.415 943.855 386.430 ;
        RECT 944.445 386.415 944.775 386.430 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 958.710 265.780 959.030 265.840 ;
        RECT 1214.470 265.780 1214.790 265.840 ;
        RECT 958.710 265.640 1214.790 265.780 ;
        RECT 958.710 265.580 959.030 265.640 ;
        RECT 1214.470 265.580 1214.790 265.640 ;
      LAYER via ;
        RECT 958.740 265.580 959.000 265.840 ;
        RECT 1214.500 265.580 1214.760 265.840 ;
      LAYER met2 ;
        RECT 956.110 510.410 956.390 514.000 ;
        RECT 956.110 510.270 958.940 510.410 ;
        RECT 956.110 510.000 956.390 510.270 ;
        RECT 958.800 265.870 958.940 510.270 ;
        RECT 958.740 265.550 959.000 265.870 ;
        RECT 1214.500 265.550 1214.760 265.870 ;
        RECT 1214.560 17.410 1214.700 265.550 ;
        RECT 1214.560 17.270 1216.080 17.410 ;
        RECT 1215.940 2.400 1216.080 17.270 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 272.920 972.370 272.980 ;
        RECT 1228.270 272.920 1228.590 272.980 ;
        RECT 972.050 272.780 1228.590 272.920 ;
        RECT 972.050 272.720 972.370 272.780 ;
        RECT 1228.270 272.720 1228.590 272.780 ;
      LAYER via ;
        RECT 972.080 272.720 972.340 272.980 ;
        RECT 1228.300 272.720 1228.560 272.980 ;
      LAYER met2 ;
        RECT 972.670 510.410 972.950 514.000 ;
        RECT 972.140 510.270 972.950 510.410 ;
        RECT 972.140 273.010 972.280 510.270 ;
        RECT 972.670 510.000 972.950 510.270 ;
        RECT 972.080 272.690 972.340 273.010 ;
        RECT 1228.300 272.690 1228.560 273.010 ;
        RECT 1228.360 17.410 1228.500 272.690 ;
        RECT 1228.360 17.270 1234.020 17.410 ;
        RECT 1233.880 2.400 1234.020 17.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 988.610 496.980 988.930 497.040 ;
        RECT 993.210 496.980 993.530 497.040 ;
        RECT 988.610 496.840 993.530 496.980 ;
        RECT 988.610 496.780 988.930 496.840 ;
        RECT 993.210 496.780 993.530 496.840 ;
        RECT 993.210 182.820 993.530 182.880 ;
        RECT 1248.970 182.820 1249.290 182.880 ;
        RECT 993.210 182.680 1249.290 182.820 ;
        RECT 993.210 182.620 993.530 182.680 ;
        RECT 1248.970 182.620 1249.290 182.680 ;
      LAYER via ;
        RECT 988.640 496.780 988.900 497.040 ;
        RECT 993.240 496.780 993.500 497.040 ;
        RECT 993.240 182.620 993.500 182.880 ;
        RECT 1249.000 182.620 1249.260 182.880 ;
      LAYER met2 ;
        RECT 988.770 510.340 989.050 514.000 ;
        RECT 988.700 510.000 989.050 510.340 ;
        RECT 988.700 497.070 988.840 510.000 ;
        RECT 988.640 496.750 988.900 497.070 ;
        RECT 993.240 496.750 993.500 497.070 ;
        RECT 993.300 182.910 993.440 496.750 ;
        RECT 993.240 182.590 993.500 182.910 ;
        RECT 1249.000 182.590 1249.260 182.910 ;
        RECT 1249.060 17.410 1249.200 182.590 ;
        RECT 1249.060 17.270 1251.960 17.410 ;
        RECT 1251.820 2.400 1251.960 17.270 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 279.720 1007.330 279.780 ;
        RECT 1262.770 279.720 1263.090 279.780 ;
        RECT 1007.010 279.580 1263.090 279.720 ;
        RECT 1007.010 279.520 1007.330 279.580 ;
        RECT 1262.770 279.520 1263.090 279.580 ;
        RECT 1262.770 17.580 1263.090 17.640 ;
        RECT 1269.210 17.580 1269.530 17.640 ;
        RECT 1262.770 17.440 1269.530 17.580 ;
        RECT 1262.770 17.380 1263.090 17.440 ;
        RECT 1269.210 17.380 1269.530 17.440 ;
      LAYER via ;
        RECT 1007.040 279.520 1007.300 279.780 ;
        RECT 1262.800 279.520 1263.060 279.780 ;
        RECT 1262.800 17.380 1263.060 17.640 ;
        RECT 1269.240 17.380 1269.500 17.640 ;
      LAYER met2 ;
        RECT 1005.330 510.410 1005.610 514.000 ;
        RECT 1005.330 510.270 1007.240 510.410 ;
        RECT 1005.330 510.000 1005.610 510.270 ;
        RECT 1007.100 279.810 1007.240 510.270 ;
        RECT 1007.040 279.490 1007.300 279.810 ;
        RECT 1262.800 279.490 1263.060 279.810 ;
        RECT 1262.860 17.670 1263.000 279.490 ;
        RECT 1262.800 17.350 1263.060 17.670 ;
        RECT 1269.240 17.350 1269.500 17.670 ;
        RECT 1269.300 2.400 1269.440 17.350 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.270 496.980 1021.590 497.040 ;
        RECT 1027.250 496.980 1027.570 497.040 ;
        RECT 1021.270 496.840 1027.570 496.980 ;
        RECT 1021.270 496.780 1021.590 496.840 ;
        RECT 1027.250 496.780 1027.570 496.840 ;
        RECT 1027.250 286.520 1027.570 286.580 ;
        RECT 1283.470 286.520 1283.790 286.580 ;
        RECT 1027.250 286.380 1283.790 286.520 ;
        RECT 1027.250 286.320 1027.570 286.380 ;
        RECT 1283.470 286.320 1283.790 286.380 ;
      LAYER via ;
        RECT 1021.300 496.780 1021.560 497.040 ;
        RECT 1027.280 496.780 1027.540 497.040 ;
        RECT 1027.280 286.320 1027.540 286.580 ;
        RECT 1283.500 286.320 1283.760 286.580 ;
      LAYER met2 ;
        RECT 1021.430 510.340 1021.710 514.000 ;
        RECT 1021.360 510.000 1021.710 510.340 ;
        RECT 1021.360 497.070 1021.500 510.000 ;
        RECT 1021.300 496.750 1021.560 497.070 ;
        RECT 1027.280 496.750 1027.540 497.070 ;
        RECT 1027.340 286.610 1027.480 496.750 ;
        RECT 1027.280 286.290 1027.540 286.610 ;
        RECT 1283.500 286.290 1283.760 286.610 ;
        RECT 1283.560 17.410 1283.700 286.290 ;
        RECT 1283.560 17.270 1287.380 17.410 ;
        RECT 1287.240 2.400 1287.380 17.270 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.830 496.980 1038.150 497.040 ;
        RECT 1041.510 496.980 1041.830 497.040 ;
        RECT 1037.830 496.840 1041.830 496.980 ;
        RECT 1037.830 496.780 1038.150 496.840 ;
        RECT 1041.510 496.780 1041.830 496.840 ;
        RECT 1041.510 293.320 1041.830 293.380 ;
        RECT 1304.170 293.320 1304.490 293.380 ;
        RECT 1041.510 293.180 1304.490 293.320 ;
        RECT 1041.510 293.120 1041.830 293.180 ;
        RECT 1304.170 293.120 1304.490 293.180 ;
      LAYER via ;
        RECT 1037.860 496.780 1038.120 497.040 ;
        RECT 1041.540 496.780 1041.800 497.040 ;
        RECT 1041.540 293.120 1041.800 293.380 ;
        RECT 1304.200 293.120 1304.460 293.380 ;
      LAYER met2 ;
        RECT 1037.990 510.340 1038.270 514.000 ;
        RECT 1037.920 510.000 1038.270 510.340 ;
        RECT 1037.920 497.070 1038.060 510.000 ;
        RECT 1037.860 496.750 1038.120 497.070 ;
        RECT 1041.540 496.750 1041.800 497.070 ;
        RECT 1041.600 293.410 1041.740 496.750 ;
        RECT 1041.540 293.090 1041.800 293.410 ;
        RECT 1304.200 293.090 1304.460 293.410 ;
        RECT 1304.260 17.410 1304.400 293.090 ;
        RECT 1304.260 17.270 1305.320 17.410 ;
        RECT 1305.180 2.400 1305.320 17.270 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 307.260 1055.630 307.320 ;
        RECT 1317.970 307.260 1318.290 307.320 ;
        RECT 1055.310 307.120 1318.290 307.260 ;
        RECT 1055.310 307.060 1055.630 307.120 ;
        RECT 1317.970 307.060 1318.290 307.120 ;
      LAYER via ;
        RECT 1055.340 307.060 1055.600 307.320 ;
        RECT 1318.000 307.060 1318.260 307.320 ;
      LAYER met2 ;
        RECT 1054.090 510.410 1054.370 514.000 ;
        RECT 1054.090 510.270 1055.540 510.410 ;
        RECT 1054.090 510.000 1054.370 510.270 ;
        RECT 1055.400 307.350 1055.540 510.270 ;
        RECT 1055.340 307.030 1055.600 307.350 ;
        RECT 1318.000 307.030 1318.260 307.350 ;
        RECT 1318.060 17.410 1318.200 307.030 ;
        RECT 1318.060 17.270 1323.260 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1070.030 496.980 1070.350 497.040 ;
        RECT 1075.550 496.980 1075.870 497.040 ;
        RECT 1070.030 496.840 1075.870 496.980 ;
        RECT 1070.030 496.780 1070.350 496.840 ;
        RECT 1075.550 496.780 1075.870 496.840 ;
        RECT 1075.550 341.600 1075.870 341.660 ;
        RECT 1338.670 341.600 1338.990 341.660 ;
        RECT 1075.550 341.460 1338.990 341.600 ;
        RECT 1075.550 341.400 1075.870 341.460 ;
        RECT 1338.670 341.400 1338.990 341.460 ;
      LAYER via ;
        RECT 1070.060 496.780 1070.320 497.040 ;
        RECT 1075.580 496.780 1075.840 497.040 ;
        RECT 1075.580 341.400 1075.840 341.660 ;
        RECT 1338.700 341.400 1338.960 341.660 ;
      LAYER met2 ;
        RECT 1070.190 510.340 1070.470 514.000 ;
        RECT 1070.120 510.000 1070.470 510.340 ;
        RECT 1070.120 497.070 1070.260 510.000 ;
        RECT 1070.060 496.750 1070.320 497.070 ;
        RECT 1075.580 496.750 1075.840 497.070 ;
        RECT 1075.640 341.690 1075.780 496.750 ;
        RECT 1075.580 341.370 1075.840 341.690 ;
        RECT 1338.700 341.370 1338.960 341.690 ;
        RECT 1338.760 17.410 1338.900 341.370 ;
        RECT 1338.760 17.270 1340.740 17.410 ;
        RECT 1340.600 2.400 1340.740 17.270 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 18.940 482.930 19.000 ;
        RECT 698.350 18.940 698.670 19.000 ;
        RECT 482.610 18.800 698.670 18.940 ;
        RECT 482.610 18.740 482.930 18.800 ;
        RECT 698.350 18.740 698.670 18.800 ;
      LAYER via ;
        RECT 482.640 18.740 482.900 19.000 ;
        RECT 698.380 18.740 698.640 19.000 ;
      LAYER met2 ;
        RECT 482.770 510.340 483.050 514.000 ;
        RECT 482.700 510.000 483.050 510.340 ;
        RECT 482.700 19.030 482.840 510.000 ;
        RECT 482.640 18.710 482.900 19.030 ;
        RECT 698.380 18.710 698.640 19.030 ;
        RECT 698.440 2.400 698.580 18.710 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1089.810 300.460 1090.130 300.520 ;
        RECT 1352.470 300.460 1352.790 300.520 ;
        RECT 1089.810 300.320 1352.790 300.460 ;
        RECT 1089.810 300.260 1090.130 300.320 ;
        RECT 1352.470 300.260 1352.790 300.320 ;
        RECT 1352.470 17.920 1352.790 17.980 ;
        RECT 1358.450 17.920 1358.770 17.980 ;
        RECT 1352.470 17.780 1358.770 17.920 ;
        RECT 1352.470 17.720 1352.790 17.780 ;
        RECT 1358.450 17.720 1358.770 17.780 ;
      LAYER via ;
        RECT 1089.840 300.260 1090.100 300.520 ;
        RECT 1352.500 300.260 1352.760 300.520 ;
        RECT 1352.500 17.720 1352.760 17.980 ;
        RECT 1358.480 17.720 1358.740 17.980 ;
      LAYER met2 ;
        RECT 1086.750 510.410 1087.030 514.000 ;
        RECT 1086.750 510.270 1090.040 510.410 ;
        RECT 1086.750 510.000 1087.030 510.270 ;
        RECT 1089.900 300.550 1090.040 510.270 ;
        RECT 1089.840 300.230 1090.100 300.550 ;
        RECT 1352.500 300.230 1352.760 300.550 ;
        RECT 1352.560 18.010 1352.700 300.230 ;
        RECT 1352.500 17.690 1352.760 18.010 ;
        RECT 1358.480 17.690 1358.740 18.010 ;
        RECT 1358.540 2.400 1358.680 17.690 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1102.690 496.980 1103.010 497.040 ;
        RECT 1107.290 496.980 1107.610 497.040 ;
        RECT 1102.690 496.840 1107.610 496.980 ;
        RECT 1102.690 496.780 1103.010 496.840 ;
        RECT 1107.290 496.780 1107.610 496.840 ;
        RECT 1107.290 314.060 1107.610 314.120 ;
        RECT 1373.170 314.060 1373.490 314.120 ;
        RECT 1107.290 313.920 1373.490 314.060 ;
        RECT 1107.290 313.860 1107.610 313.920 ;
        RECT 1373.170 313.860 1373.490 313.920 ;
      LAYER via ;
        RECT 1102.720 496.780 1102.980 497.040 ;
        RECT 1107.320 496.780 1107.580 497.040 ;
        RECT 1107.320 313.860 1107.580 314.120 ;
        RECT 1373.200 313.860 1373.460 314.120 ;
      LAYER met2 ;
        RECT 1102.850 510.340 1103.130 514.000 ;
        RECT 1102.780 510.000 1103.130 510.340 ;
        RECT 1102.780 497.070 1102.920 510.000 ;
        RECT 1102.720 496.750 1102.980 497.070 ;
        RECT 1107.320 496.750 1107.580 497.070 ;
        RECT 1107.380 314.150 1107.520 496.750 ;
        RECT 1107.320 313.830 1107.580 314.150 ;
        RECT 1373.200 313.830 1373.460 314.150 ;
        RECT 1373.260 17.410 1373.400 313.830 ;
        RECT 1373.260 17.270 1376.620 17.410 ;
        RECT 1376.480 2.400 1376.620 17.270 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1119.250 496.980 1119.570 497.040 ;
        RECT 1124.310 496.980 1124.630 497.040 ;
        RECT 1119.250 496.840 1124.630 496.980 ;
        RECT 1119.250 496.780 1119.570 496.840 ;
        RECT 1124.310 496.780 1124.630 496.840 ;
        RECT 1124.310 355.200 1124.630 355.260 ;
        RECT 1393.870 355.200 1394.190 355.260 ;
        RECT 1124.310 355.060 1394.190 355.200 ;
        RECT 1124.310 355.000 1124.630 355.060 ;
        RECT 1393.870 355.000 1394.190 355.060 ;
      LAYER via ;
        RECT 1119.280 496.780 1119.540 497.040 ;
        RECT 1124.340 496.780 1124.600 497.040 ;
        RECT 1124.340 355.000 1124.600 355.260 ;
        RECT 1393.900 355.000 1394.160 355.260 ;
      LAYER met2 ;
        RECT 1119.410 510.340 1119.690 514.000 ;
        RECT 1119.340 510.000 1119.690 510.340 ;
        RECT 1119.340 497.070 1119.480 510.000 ;
        RECT 1119.280 496.750 1119.540 497.070 ;
        RECT 1124.340 496.750 1124.600 497.070 ;
        RECT 1124.400 355.290 1124.540 496.750 ;
        RECT 1124.340 354.970 1124.600 355.290 ;
        RECT 1393.900 354.970 1394.160 355.290 ;
        RECT 1393.960 17.410 1394.100 354.970 ;
        RECT 1393.960 17.270 1394.560 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 320.860 1138.430 320.920 ;
        RECT 1407.670 320.860 1407.990 320.920 ;
        RECT 1138.110 320.720 1407.990 320.860 ;
        RECT 1138.110 320.660 1138.430 320.720 ;
        RECT 1407.670 320.660 1407.990 320.720 ;
      LAYER via ;
        RECT 1138.140 320.660 1138.400 320.920 ;
        RECT 1407.700 320.660 1407.960 320.920 ;
      LAYER met2 ;
        RECT 1135.510 510.410 1135.790 514.000 ;
        RECT 1135.510 510.270 1138.340 510.410 ;
        RECT 1135.510 510.000 1135.790 510.270 ;
        RECT 1138.200 320.950 1138.340 510.270 ;
        RECT 1138.140 320.630 1138.400 320.950 ;
        RECT 1407.700 320.630 1407.960 320.950 ;
        RECT 1407.760 17.410 1407.900 320.630 ;
        RECT 1407.760 17.270 1412.500 17.410 ;
        RECT 1412.360 2.400 1412.500 17.270 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.450 348.400 1151.770 348.460 ;
        RECT 1428.370 348.400 1428.690 348.460 ;
        RECT 1151.450 348.260 1428.690 348.400 ;
        RECT 1151.450 348.200 1151.770 348.260 ;
        RECT 1428.370 348.200 1428.690 348.260 ;
      LAYER via ;
        RECT 1151.480 348.200 1151.740 348.460 ;
        RECT 1428.400 348.200 1428.660 348.460 ;
      LAYER met2 ;
        RECT 1152.070 510.410 1152.350 514.000 ;
        RECT 1151.540 510.270 1152.350 510.410 ;
        RECT 1151.540 348.490 1151.680 510.270 ;
        RECT 1152.070 510.000 1152.350 510.270 ;
        RECT 1151.480 348.170 1151.740 348.490 ;
        RECT 1428.400 348.170 1428.660 348.490 ;
        RECT 1428.460 17.410 1428.600 348.170 ;
        RECT 1428.460 17.270 1429.980 17.410 ;
        RECT 1429.840 2.400 1429.980 17.270 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.010 503.440 1168.330 503.500 ;
        RECT 1172.610 503.440 1172.930 503.500 ;
        RECT 1168.010 503.300 1172.930 503.440 ;
        RECT 1168.010 503.240 1168.330 503.300 ;
        RECT 1172.610 503.240 1172.930 503.300 ;
        RECT 1172.610 327.660 1172.930 327.720 ;
        RECT 1442.170 327.660 1442.490 327.720 ;
        RECT 1172.610 327.520 1442.490 327.660 ;
        RECT 1172.610 327.460 1172.930 327.520 ;
        RECT 1442.170 327.460 1442.490 327.520 ;
      LAYER via ;
        RECT 1168.040 503.240 1168.300 503.500 ;
        RECT 1172.640 503.240 1172.900 503.500 ;
        RECT 1172.640 327.460 1172.900 327.720 ;
        RECT 1442.200 327.460 1442.460 327.720 ;
      LAYER met2 ;
        RECT 1168.170 510.340 1168.450 514.000 ;
        RECT 1168.100 510.000 1168.450 510.340 ;
        RECT 1168.100 503.530 1168.240 510.000 ;
        RECT 1168.040 503.210 1168.300 503.530 ;
        RECT 1172.640 503.210 1172.900 503.530 ;
        RECT 1172.700 327.750 1172.840 503.210 ;
        RECT 1172.640 327.430 1172.900 327.750 ;
        RECT 1442.200 327.430 1442.460 327.750 ;
        RECT 1442.260 17.410 1442.400 327.430 ;
        RECT 1442.260 17.270 1447.920 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 334.800 1186.730 334.860 ;
        RECT 1462.870 334.800 1463.190 334.860 ;
        RECT 1186.410 334.660 1463.190 334.800 ;
        RECT 1186.410 334.600 1186.730 334.660 ;
        RECT 1462.870 334.600 1463.190 334.660 ;
      LAYER via ;
        RECT 1186.440 334.600 1186.700 334.860 ;
        RECT 1462.900 334.600 1463.160 334.860 ;
      LAYER met2 ;
        RECT 1184.730 510.410 1185.010 514.000 ;
        RECT 1184.730 510.270 1186.640 510.410 ;
        RECT 1184.730 510.000 1185.010 510.270 ;
        RECT 1186.500 334.890 1186.640 510.270 ;
        RECT 1186.440 334.570 1186.700 334.890 ;
        RECT 1462.900 334.570 1463.160 334.890 ;
        RECT 1462.960 17.410 1463.100 334.570 ;
        RECT 1462.960 17.270 1465.860 17.410 ;
        RECT 1465.720 2.400 1465.860 17.270 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.670 503.100 1200.990 503.160 ;
        RECT 1206.650 503.100 1206.970 503.160 ;
        RECT 1200.670 502.960 1206.970 503.100 ;
        RECT 1200.670 502.900 1200.990 502.960 ;
        RECT 1206.650 502.900 1206.970 502.960 ;
        RECT 1206.650 265.440 1206.970 265.500 ;
        RECT 1483.570 265.440 1483.890 265.500 ;
        RECT 1206.650 265.300 1483.890 265.440 ;
        RECT 1206.650 265.240 1206.970 265.300 ;
        RECT 1483.570 265.240 1483.890 265.300 ;
      LAYER via ;
        RECT 1200.700 502.900 1200.960 503.160 ;
        RECT 1206.680 502.900 1206.940 503.160 ;
        RECT 1206.680 265.240 1206.940 265.500 ;
        RECT 1483.600 265.240 1483.860 265.500 ;
      LAYER met2 ;
        RECT 1200.830 510.340 1201.110 514.000 ;
        RECT 1200.760 510.000 1201.110 510.340 ;
        RECT 1200.760 503.190 1200.900 510.000 ;
        RECT 1200.700 502.870 1200.960 503.190 ;
        RECT 1206.680 502.870 1206.940 503.190 ;
        RECT 1206.740 265.530 1206.880 502.870 ;
        RECT 1206.680 265.210 1206.940 265.530 ;
        RECT 1483.600 265.210 1483.860 265.530 ;
        RECT 1483.660 2.400 1483.800 265.210 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1217.230 503.440 1217.550 503.500 ;
        RECT 1220.910 503.440 1221.230 503.500 ;
        RECT 1217.230 503.300 1221.230 503.440 ;
        RECT 1217.230 503.240 1217.550 503.300 ;
        RECT 1220.910 503.240 1221.230 503.300 ;
        RECT 1220.910 272.580 1221.230 272.640 ;
        RECT 1497.370 272.580 1497.690 272.640 ;
        RECT 1220.910 272.440 1497.690 272.580 ;
        RECT 1220.910 272.380 1221.230 272.440 ;
        RECT 1497.370 272.380 1497.690 272.440 ;
      LAYER via ;
        RECT 1217.260 503.240 1217.520 503.500 ;
        RECT 1220.940 503.240 1221.200 503.500 ;
        RECT 1220.940 272.380 1221.200 272.640 ;
        RECT 1497.400 272.380 1497.660 272.640 ;
      LAYER met2 ;
        RECT 1217.390 510.340 1217.670 514.000 ;
        RECT 1217.320 510.000 1217.670 510.340 ;
        RECT 1217.320 503.530 1217.460 510.000 ;
        RECT 1217.260 503.210 1217.520 503.530 ;
        RECT 1220.940 503.210 1221.200 503.530 ;
        RECT 1221.000 272.670 1221.140 503.210 ;
        RECT 1220.940 272.350 1221.200 272.670 ;
        RECT 1497.400 272.350 1497.660 272.670 ;
        RECT 1497.460 17.410 1497.600 272.350 ;
        RECT 1497.460 17.270 1501.740 17.410 ;
        RECT 1501.600 2.400 1501.740 17.270 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 362.340 1235.030 362.400 ;
        RECT 1518.070 362.340 1518.390 362.400 ;
        RECT 1234.710 362.200 1518.390 362.340 ;
        RECT 1234.710 362.140 1235.030 362.200 ;
        RECT 1518.070 362.140 1518.390 362.200 ;
      LAYER via ;
        RECT 1234.740 362.140 1235.000 362.400 ;
        RECT 1518.100 362.140 1518.360 362.400 ;
      LAYER met2 ;
        RECT 1233.490 510.410 1233.770 514.000 ;
        RECT 1233.490 510.270 1234.940 510.410 ;
        RECT 1233.490 510.000 1233.770 510.270 ;
        RECT 1234.800 362.430 1234.940 510.270 ;
        RECT 1234.740 362.110 1235.000 362.430 ;
        RECT 1518.100 362.110 1518.360 362.430 ;
        RECT 1518.160 17.410 1518.300 362.110 ;
        RECT 1518.160 17.270 1519.220 17.410 ;
        RECT 1519.080 2.400 1519.220 17.270 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 499.170 503.440 499.490 503.500 ;
        RECT 503.310 503.440 503.630 503.500 ;
        RECT 499.170 503.300 503.630 503.440 ;
        RECT 499.170 503.240 499.490 503.300 ;
        RECT 503.310 503.240 503.630 503.300 ;
        RECT 503.310 19.280 503.630 19.340 ;
        RECT 716.290 19.280 716.610 19.340 ;
        RECT 503.310 19.140 716.610 19.280 ;
        RECT 503.310 19.080 503.630 19.140 ;
        RECT 716.290 19.080 716.610 19.140 ;
      LAYER via ;
        RECT 499.200 503.240 499.460 503.500 ;
        RECT 503.340 503.240 503.600 503.500 ;
        RECT 503.340 19.080 503.600 19.340 ;
        RECT 716.320 19.080 716.580 19.340 ;
      LAYER met2 ;
        RECT 499.330 510.340 499.610 514.000 ;
        RECT 499.260 510.000 499.610 510.340 ;
        RECT 499.260 503.530 499.400 510.000 ;
        RECT 499.200 503.210 499.460 503.530 ;
        RECT 503.340 503.210 503.600 503.530 ;
        RECT 503.400 19.370 503.540 503.210 ;
        RECT 503.340 19.050 503.600 19.370 ;
        RECT 716.320 19.050 716.580 19.370 ;
        RECT 716.380 2.400 716.520 19.050 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1249.890 496.980 1250.210 497.040 ;
        RECT 1254.950 496.980 1255.270 497.040 ;
        RECT 1249.890 496.840 1255.270 496.980 ;
        RECT 1249.890 496.780 1250.210 496.840 ;
        RECT 1254.950 496.780 1255.270 496.840 ;
        RECT 1254.950 279.380 1255.270 279.440 ;
        RECT 1531.870 279.380 1532.190 279.440 ;
        RECT 1254.950 279.240 1532.190 279.380 ;
        RECT 1254.950 279.180 1255.270 279.240 ;
        RECT 1531.870 279.180 1532.190 279.240 ;
      LAYER via ;
        RECT 1249.920 496.780 1250.180 497.040 ;
        RECT 1254.980 496.780 1255.240 497.040 ;
        RECT 1254.980 279.180 1255.240 279.440 ;
        RECT 1531.900 279.180 1532.160 279.440 ;
      LAYER met2 ;
        RECT 1250.050 510.340 1250.330 514.000 ;
        RECT 1249.980 510.000 1250.330 510.340 ;
        RECT 1249.980 497.070 1250.120 510.000 ;
        RECT 1249.920 496.750 1250.180 497.070 ;
        RECT 1254.980 496.750 1255.240 497.070 ;
        RECT 1255.040 279.470 1255.180 496.750 ;
        RECT 1254.980 279.150 1255.240 279.470 ;
        RECT 1531.900 279.150 1532.160 279.470 ;
        RECT 1531.960 17.410 1532.100 279.150 ;
        RECT 1531.960 17.270 1537.160 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 286.180 1269.530 286.240 ;
        RECT 1552.570 286.180 1552.890 286.240 ;
        RECT 1269.210 286.040 1552.890 286.180 ;
        RECT 1269.210 285.980 1269.530 286.040 ;
        RECT 1552.570 285.980 1552.890 286.040 ;
      LAYER via ;
        RECT 1269.240 285.980 1269.500 286.240 ;
        RECT 1552.600 285.980 1552.860 286.240 ;
      LAYER met2 ;
        RECT 1266.150 510.410 1266.430 514.000 ;
        RECT 1266.150 510.270 1269.440 510.410 ;
        RECT 1266.150 510.000 1266.430 510.270 ;
        RECT 1269.300 286.270 1269.440 510.270 ;
        RECT 1269.240 285.950 1269.500 286.270 ;
        RECT 1552.600 285.950 1552.860 286.270 ;
        RECT 1552.660 17.410 1552.800 285.950 ;
        RECT 1552.660 17.270 1555.100 17.410 ;
        RECT 1554.960 2.400 1555.100 17.270 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1282.550 369.480 1282.870 369.540 ;
        RECT 1566.370 369.480 1566.690 369.540 ;
        RECT 1282.550 369.340 1566.690 369.480 ;
        RECT 1282.550 369.280 1282.870 369.340 ;
        RECT 1566.370 369.280 1566.690 369.340 ;
        RECT 1566.370 17.580 1566.690 17.640 ;
        RECT 1572.810 17.580 1573.130 17.640 ;
        RECT 1566.370 17.440 1573.130 17.580 ;
        RECT 1566.370 17.380 1566.690 17.440 ;
        RECT 1572.810 17.380 1573.130 17.440 ;
      LAYER via ;
        RECT 1282.580 369.280 1282.840 369.540 ;
        RECT 1566.400 369.280 1566.660 369.540 ;
        RECT 1566.400 17.380 1566.660 17.640 ;
        RECT 1572.840 17.380 1573.100 17.640 ;
      LAYER met2 ;
        RECT 1282.710 510.340 1282.990 514.000 ;
        RECT 1282.640 510.000 1282.990 510.340 ;
        RECT 1282.640 369.570 1282.780 510.000 ;
        RECT 1282.580 369.250 1282.840 369.570 ;
        RECT 1566.400 369.250 1566.660 369.570 ;
        RECT 1566.460 17.670 1566.600 369.250 ;
        RECT 1566.400 17.350 1566.660 17.670 ;
        RECT 1572.840 17.350 1573.100 17.670 ;
        RECT 1572.900 2.400 1573.040 17.350 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1298.650 496.980 1298.970 497.040 ;
        RECT 1303.710 496.980 1304.030 497.040 ;
        RECT 1298.650 496.840 1304.030 496.980 ;
        RECT 1298.650 496.780 1298.970 496.840 ;
        RECT 1303.710 496.780 1304.030 496.840 ;
        RECT 1303.710 375.940 1304.030 376.000 ;
        RECT 1587.070 375.940 1587.390 376.000 ;
        RECT 1303.710 375.800 1587.390 375.940 ;
        RECT 1303.710 375.740 1304.030 375.800 ;
        RECT 1587.070 375.740 1587.390 375.800 ;
      LAYER via ;
        RECT 1298.680 496.780 1298.940 497.040 ;
        RECT 1303.740 496.780 1304.000 497.040 ;
        RECT 1303.740 375.740 1304.000 376.000 ;
        RECT 1587.100 375.740 1587.360 376.000 ;
      LAYER met2 ;
        RECT 1298.810 510.340 1299.090 514.000 ;
        RECT 1298.740 510.000 1299.090 510.340 ;
        RECT 1298.740 497.070 1298.880 510.000 ;
        RECT 1298.680 496.750 1298.940 497.070 ;
        RECT 1303.740 496.750 1304.000 497.070 ;
        RECT 1303.800 376.030 1303.940 496.750 ;
        RECT 1303.740 375.710 1304.000 376.030 ;
        RECT 1587.100 375.710 1587.360 376.030 ;
        RECT 1587.160 16.730 1587.300 375.710 ;
        RECT 1587.160 16.590 1590.520 16.730 ;
        RECT 1590.380 2.400 1590.520 16.590 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 306.920 1317.830 306.980 ;
        RECT 1607.770 306.920 1608.090 306.980 ;
        RECT 1317.510 306.780 1608.090 306.920 ;
        RECT 1317.510 306.720 1317.830 306.780 ;
        RECT 1607.770 306.720 1608.090 306.780 ;
      LAYER via ;
        RECT 1317.540 306.720 1317.800 306.980 ;
        RECT 1607.800 306.720 1608.060 306.980 ;
      LAYER met2 ;
        RECT 1315.370 510.410 1315.650 514.000 ;
        RECT 1315.370 510.270 1317.740 510.410 ;
        RECT 1315.370 510.000 1315.650 510.270 ;
        RECT 1317.600 307.010 1317.740 510.270 ;
        RECT 1317.540 306.690 1317.800 307.010 ;
        RECT 1607.800 306.690 1608.060 307.010 ;
        RECT 1607.860 17.410 1608.000 306.690 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 107.000 1331.630 107.060 ;
        RECT 1621.570 107.000 1621.890 107.060 ;
        RECT 1331.310 106.860 1621.890 107.000 ;
        RECT 1331.310 106.800 1331.630 106.860 ;
        RECT 1621.570 106.800 1621.890 106.860 ;
      LAYER via ;
        RECT 1331.340 106.800 1331.600 107.060 ;
        RECT 1621.600 106.800 1621.860 107.060 ;
      LAYER met2 ;
        RECT 1331.470 510.340 1331.750 514.000 ;
        RECT 1331.400 510.000 1331.750 510.340 ;
        RECT 1331.400 107.090 1331.540 510.000 ;
        RECT 1331.340 106.770 1331.600 107.090 ;
        RECT 1621.600 106.770 1621.860 107.090 ;
        RECT 1621.660 16.730 1621.800 106.770 ;
        RECT 1621.660 16.590 1626.400 16.730 ;
        RECT 1626.260 2.400 1626.400 16.590 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.870 496.980 1348.190 497.040 ;
        RECT 1352.010 496.980 1352.330 497.040 ;
        RECT 1347.870 496.840 1352.330 496.980 ;
        RECT 1347.870 496.780 1348.190 496.840 ;
        RECT 1352.010 496.780 1352.330 496.840 ;
        RECT 1352.010 300.120 1352.330 300.180 ;
        RECT 1642.270 300.120 1642.590 300.180 ;
        RECT 1352.010 299.980 1642.590 300.120 ;
        RECT 1352.010 299.920 1352.330 299.980 ;
        RECT 1642.270 299.920 1642.590 299.980 ;
      LAYER via ;
        RECT 1347.900 496.780 1348.160 497.040 ;
        RECT 1352.040 496.780 1352.300 497.040 ;
        RECT 1352.040 299.920 1352.300 300.180 ;
        RECT 1642.300 299.920 1642.560 300.180 ;
      LAYER met2 ;
        RECT 1348.030 510.340 1348.310 514.000 ;
        RECT 1347.960 510.000 1348.310 510.340 ;
        RECT 1347.960 497.070 1348.100 510.000 ;
        RECT 1347.900 496.750 1348.160 497.070 ;
        RECT 1352.040 496.750 1352.300 497.070 ;
        RECT 1352.100 300.210 1352.240 496.750 ;
        RECT 1352.040 299.890 1352.300 300.210 ;
        RECT 1642.300 299.890 1642.560 300.210 ;
        RECT 1642.360 17.410 1642.500 299.890 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 341.600 1366.130 341.660 ;
        RECT 1656.070 341.600 1656.390 341.660 ;
        RECT 1365.810 341.460 1656.390 341.600 ;
        RECT 1365.810 341.400 1366.130 341.460 ;
        RECT 1656.070 341.400 1656.390 341.460 ;
        RECT 1656.070 17.920 1656.390 17.980 ;
        RECT 1662.050 17.920 1662.370 17.980 ;
        RECT 1656.070 17.780 1662.370 17.920 ;
        RECT 1656.070 17.720 1656.390 17.780 ;
        RECT 1662.050 17.720 1662.370 17.780 ;
      LAYER via ;
        RECT 1365.840 341.400 1366.100 341.660 ;
        RECT 1656.100 341.400 1656.360 341.660 ;
        RECT 1656.100 17.720 1656.360 17.980 ;
        RECT 1662.080 17.720 1662.340 17.980 ;
      LAYER met2 ;
        RECT 1364.130 510.410 1364.410 514.000 ;
        RECT 1364.130 510.270 1366.040 510.410 ;
        RECT 1364.130 510.000 1364.410 510.270 ;
        RECT 1365.900 341.690 1366.040 510.270 ;
        RECT 1365.840 341.370 1366.100 341.690 ;
        RECT 1656.100 341.370 1656.360 341.690 ;
        RECT 1656.160 18.010 1656.300 341.370 ;
        RECT 1656.100 17.690 1656.360 18.010 ;
        RECT 1662.080 17.690 1662.340 18.010 ;
        RECT 1662.140 2.400 1662.280 17.690 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.530 496.980 1380.850 497.040 ;
        RECT 1386.050 496.980 1386.370 497.040 ;
        RECT 1380.530 496.840 1386.370 496.980 ;
        RECT 1380.530 496.780 1380.850 496.840 ;
        RECT 1386.050 496.780 1386.370 496.840 ;
        RECT 1386.050 314.060 1386.370 314.120 ;
        RECT 1676.770 314.060 1677.090 314.120 ;
        RECT 1386.050 313.920 1677.090 314.060 ;
        RECT 1386.050 313.860 1386.370 313.920 ;
        RECT 1676.770 313.860 1677.090 313.920 ;
      LAYER via ;
        RECT 1380.560 496.780 1380.820 497.040 ;
        RECT 1386.080 496.780 1386.340 497.040 ;
        RECT 1386.080 313.860 1386.340 314.120 ;
        RECT 1676.800 313.860 1677.060 314.120 ;
      LAYER met2 ;
        RECT 1380.690 510.340 1380.970 514.000 ;
        RECT 1380.620 510.000 1380.970 510.340 ;
        RECT 1380.620 497.070 1380.760 510.000 ;
        RECT 1380.560 496.750 1380.820 497.070 ;
        RECT 1386.080 496.750 1386.340 497.070 ;
        RECT 1386.140 314.150 1386.280 496.750 ;
        RECT 1386.080 313.830 1386.340 314.150 ;
        RECT 1676.800 313.830 1677.060 314.150 ;
        RECT 1676.860 17.410 1677.000 313.830 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1396.630 496.980 1396.950 497.040 ;
        RECT 1400.310 496.980 1400.630 497.040 ;
        RECT 1396.630 496.840 1400.630 496.980 ;
        RECT 1396.630 496.780 1396.950 496.840 ;
        RECT 1400.310 496.780 1400.630 496.840 ;
        RECT 1400.310 355.540 1400.630 355.600 ;
        RECT 1697.470 355.540 1697.790 355.600 ;
        RECT 1400.310 355.400 1697.790 355.540 ;
        RECT 1400.310 355.340 1400.630 355.400 ;
        RECT 1697.470 355.340 1697.790 355.400 ;
      LAYER via ;
        RECT 1396.660 496.780 1396.920 497.040 ;
        RECT 1400.340 496.780 1400.600 497.040 ;
        RECT 1400.340 355.340 1400.600 355.600 ;
        RECT 1697.500 355.340 1697.760 355.600 ;
      LAYER met2 ;
        RECT 1396.790 510.340 1397.070 514.000 ;
        RECT 1396.720 510.000 1397.070 510.340 ;
        RECT 1396.720 497.070 1396.860 510.000 ;
        RECT 1396.660 496.750 1396.920 497.070 ;
        RECT 1400.340 496.750 1400.600 497.070 ;
        RECT 1400.400 355.630 1400.540 496.750 ;
        RECT 1400.340 355.310 1400.600 355.630 ;
        RECT 1697.500 355.310 1697.760 355.630 ;
        RECT 1697.560 2.400 1697.700 355.310 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 18.600 517.430 18.660 ;
        RECT 734.230 18.600 734.550 18.660 ;
        RECT 517.110 18.460 734.550 18.600 ;
        RECT 517.110 18.400 517.430 18.460 ;
        RECT 734.230 18.400 734.550 18.460 ;
      LAYER via ;
        RECT 517.140 18.400 517.400 18.660 ;
        RECT 734.260 18.400 734.520 18.660 ;
      LAYER met2 ;
        RECT 515.430 510.410 515.710 514.000 ;
        RECT 515.430 510.270 517.340 510.410 ;
        RECT 515.430 510.000 515.710 510.270 ;
        RECT 517.200 18.690 517.340 510.270 ;
        RECT 517.140 18.370 517.400 18.690 ;
        RECT 734.260 18.370 734.520 18.690 ;
        RECT 734.320 2.400 734.460 18.370 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 320.860 1414.430 320.920 ;
        RECT 1711.270 320.860 1711.590 320.920 ;
        RECT 1414.110 320.720 1711.590 320.860 ;
        RECT 1414.110 320.660 1414.430 320.720 ;
        RECT 1711.270 320.660 1711.590 320.720 ;
      LAYER via ;
        RECT 1414.140 320.660 1414.400 320.920 ;
        RECT 1711.300 320.660 1711.560 320.920 ;
      LAYER met2 ;
        RECT 1413.350 510.410 1413.630 514.000 ;
        RECT 1413.350 510.270 1414.340 510.410 ;
        RECT 1413.350 510.000 1413.630 510.270 ;
        RECT 1414.200 320.950 1414.340 510.270 ;
        RECT 1414.140 320.630 1414.400 320.950 ;
        RECT 1711.300 320.630 1711.560 320.950 ;
        RECT 1711.360 17.410 1711.500 320.630 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.290 496.980 1429.610 497.040 ;
        RECT 1434.810 496.980 1435.130 497.040 ;
        RECT 1429.290 496.840 1435.130 496.980 ;
        RECT 1429.290 496.780 1429.610 496.840 ;
        RECT 1434.810 496.780 1435.130 496.840 ;
        RECT 1434.810 348.400 1435.130 348.460 ;
        RECT 1731.970 348.400 1732.290 348.460 ;
        RECT 1434.810 348.260 1732.290 348.400 ;
        RECT 1434.810 348.200 1435.130 348.260 ;
        RECT 1731.970 348.200 1732.290 348.260 ;
      LAYER via ;
        RECT 1429.320 496.780 1429.580 497.040 ;
        RECT 1434.840 496.780 1435.100 497.040 ;
        RECT 1434.840 348.200 1435.100 348.460 ;
        RECT 1732.000 348.200 1732.260 348.460 ;
      LAYER met2 ;
        RECT 1429.450 510.340 1429.730 514.000 ;
        RECT 1429.380 510.000 1429.730 510.340 ;
        RECT 1429.380 497.070 1429.520 510.000 ;
        RECT 1429.320 496.750 1429.580 497.070 ;
        RECT 1434.840 496.750 1435.100 497.070 ;
        RECT 1434.900 348.490 1435.040 496.750 ;
        RECT 1434.840 348.170 1435.100 348.490 ;
        RECT 1732.000 348.170 1732.260 348.490 ;
        RECT 1732.060 17.410 1732.200 348.170 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 327.660 1448.930 327.720 ;
        RECT 1745.770 327.660 1746.090 327.720 ;
        RECT 1448.610 327.520 1746.090 327.660 ;
        RECT 1448.610 327.460 1448.930 327.520 ;
        RECT 1745.770 327.460 1746.090 327.520 ;
      LAYER via ;
        RECT 1448.640 327.460 1448.900 327.720 ;
        RECT 1745.800 327.460 1746.060 327.720 ;
      LAYER met2 ;
        RECT 1446.010 510.410 1446.290 514.000 ;
        RECT 1446.010 510.270 1448.840 510.410 ;
        RECT 1446.010 510.000 1446.290 510.270 ;
        RECT 1448.700 327.750 1448.840 510.270 ;
        RECT 1448.640 327.430 1448.900 327.750 ;
        RECT 1745.800 327.430 1746.060 327.750 ;
        RECT 1745.860 17.410 1746.000 327.430 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1766.545 241.485 1766.715 289.595 ;
      LAYER mcon ;
        RECT 1766.545 289.425 1766.715 289.595 ;
      LAYER met1 ;
        RECT 1461.950 334.460 1462.270 334.520 ;
        RECT 1766.930 334.460 1767.250 334.520 ;
        RECT 1461.950 334.320 1767.250 334.460 ;
        RECT 1461.950 334.260 1462.270 334.320 ;
        RECT 1766.930 334.260 1767.250 334.320 ;
        RECT 1766.470 289.580 1766.790 289.640 ;
        RECT 1766.275 289.440 1766.790 289.580 ;
        RECT 1766.470 289.380 1766.790 289.440 ;
        RECT 1766.470 241.640 1766.790 241.700 ;
        RECT 1766.275 241.500 1766.790 241.640 ;
        RECT 1766.470 241.440 1766.790 241.500 ;
        RECT 1766.470 193.020 1766.790 193.080 ;
        RECT 1766.930 193.020 1767.250 193.080 ;
        RECT 1766.470 192.880 1767.250 193.020 ;
        RECT 1766.470 192.820 1766.790 192.880 ;
        RECT 1766.930 192.820 1767.250 192.880 ;
        RECT 1766.470 137.940 1766.790 138.000 ;
        RECT 1769.230 137.940 1769.550 138.000 ;
        RECT 1766.470 137.800 1769.550 137.940 ;
        RECT 1766.470 137.740 1766.790 137.800 ;
        RECT 1769.230 137.740 1769.550 137.800 ;
        RECT 1768.770 47.980 1769.090 48.240 ;
        RECT 1768.860 47.560 1769.000 47.980 ;
        RECT 1768.770 47.300 1769.090 47.560 ;
      LAYER via ;
        RECT 1461.980 334.260 1462.240 334.520 ;
        RECT 1766.960 334.260 1767.220 334.520 ;
        RECT 1766.500 289.380 1766.760 289.640 ;
        RECT 1766.500 241.440 1766.760 241.700 ;
        RECT 1766.500 192.820 1766.760 193.080 ;
        RECT 1766.960 192.820 1767.220 193.080 ;
        RECT 1766.500 137.740 1766.760 138.000 ;
        RECT 1769.260 137.740 1769.520 138.000 ;
        RECT 1768.800 47.980 1769.060 48.240 ;
        RECT 1768.800 47.300 1769.060 47.560 ;
      LAYER met2 ;
        RECT 1462.110 510.340 1462.390 514.000 ;
        RECT 1462.040 510.000 1462.390 510.340 ;
        RECT 1462.040 334.550 1462.180 510.000 ;
        RECT 1461.980 334.230 1462.240 334.550 ;
        RECT 1766.960 334.230 1767.220 334.550 ;
        RECT 1767.020 290.090 1767.160 334.230 ;
        RECT 1766.560 289.950 1767.160 290.090 ;
        RECT 1766.560 289.670 1766.700 289.950 ;
        RECT 1766.500 289.350 1766.760 289.670 ;
        RECT 1766.500 241.410 1766.760 241.730 ;
        RECT 1766.560 194.210 1766.700 241.410 ;
        RECT 1766.560 194.070 1767.160 194.210 ;
        RECT 1767.020 193.530 1767.160 194.070 ;
        RECT 1766.560 193.390 1767.160 193.530 ;
        RECT 1766.560 193.110 1766.700 193.390 ;
        RECT 1766.500 192.790 1766.760 193.110 ;
        RECT 1766.960 192.790 1767.220 193.110 ;
        RECT 1767.020 145.250 1767.160 192.790 ;
        RECT 1766.560 145.110 1767.160 145.250 ;
        RECT 1766.560 138.030 1766.700 145.110 ;
        RECT 1766.500 137.710 1766.760 138.030 ;
        RECT 1769.260 137.710 1769.520 138.030 ;
        RECT 1769.320 61.610 1769.460 137.710 ;
        RECT 1768.860 61.470 1769.460 61.610 ;
        RECT 1768.860 48.270 1769.000 61.470 ;
        RECT 1768.800 47.950 1769.060 48.270 ;
        RECT 1768.800 47.270 1769.060 47.590 ;
        RECT 1768.860 2.400 1769.000 47.270 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1478.050 501.060 1478.370 501.120 ;
        RECT 1483.110 501.060 1483.430 501.120 ;
        RECT 1478.050 500.920 1483.430 501.060 ;
        RECT 1478.050 500.860 1478.370 500.920 ;
        RECT 1483.110 500.860 1483.430 500.920 ;
        RECT 1483.110 382.740 1483.430 382.800 ;
        RECT 1780.270 382.740 1780.590 382.800 ;
        RECT 1483.110 382.600 1780.590 382.740 ;
        RECT 1483.110 382.540 1483.430 382.600 ;
        RECT 1780.270 382.540 1780.590 382.600 ;
        RECT 1780.270 37.980 1780.590 38.040 ;
        RECT 1786.710 37.980 1787.030 38.040 ;
        RECT 1780.270 37.840 1787.030 37.980 ;
        RECT 1780.270 37.780 1780.590 37.840 ;
        RECT 1786.710 37.780 1787.030 37.840 ;
      LAYER via ;
        RECT 1478.080 500.860 1478.340 501.120 ;
        RECT 1483.140 500.860 1483.400 501.120 ;
        RECT 1483.140 382.540 1483.400 382.800 ;
        RECT 1780.300 382.540 1780.560 382.800 ;
        RECT 1780.300 37.780 1780.560 38.040 ;
        RECT 1786.740 37.780 1787.000 38.040 ;
      LAYER met2 ;
        RECT 1478.210 510.340 1478.490 514.000 ;
        RECT 1478.140 510.000 1478.490 510.340 ;
        RECT 1478.140 501.150 1478.280 510.000 ;
        RECT 1478.080 500.830 1478.340 501.150 ;
        RECT 1483.140 500.830 1483.400 501.150 ;
        RECT 1483.200 382.830 1483.340 500.830 ;
        RECT 1483.140 382.510 1483.400 382.830 ;
        RECT 1780.300 382.510 1780.560 382.830 ;
        RECT 1780.360 38.070 1780.500 382.510 ;
        RECT 1780.300 37.750 1780.560 38.070 ;
        RECT 1786.740 37.750 1787.000 38.070 ;
        RECT 1786.800 2.400 1786.940 37.750 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 389.880 1497.230 389.940 ;
        RECT 1800.970 389.880 1801.290 389.940 ;
        RECT 1496.910 389.740 1801.290 389.880 ;
        RECT 1496.910 389.680 1497.230 389.740 ;
        RECT 1800.970 389.680 1801.290 389.740 ;
      LAYER via ;
        RECT 1496.940 389.680 1497.200 389.940 ;
        RECT 1801.000 389.680 1801.260 389.940 ;
      LAYER met2 ;
        RECT 1494.770 510.410 1495.050 514.000 ;
        RECT 1494.770 510.270 1497.140 510.410 ;
        RECT 1494.770 510.000 1495.050 510.270 ;
        RECT 1497.000 389.970 1497.140 510.270 ;
        RECT 1496.940 389.650 1497.200 389.970 ;
        RECT 1801.000 389.650 1801.260 389.970 ;
        RECT 1801.060 17.410 1801.200 389.650 ;
        RECT 1801.060 17.270 1804.880 17.410 ;
        RECT 1804.740 2.400 1804.880 17.270 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.250 397.020 1510.570 397.080 ;
        RECT 1821.670 397.020 1821.990 397.080 ;
        RECT 1510.250 396.880 1821.990 397.020 ;
        RECT 1510.250 396.820 1510.570 396.880 ;
        RECT 1821.670 396.820 1821.990 396.880 ;
      LAYER via ;
        RECT 1510.280 396.820 1510.540 397.080 ;
        RECT 1821.700 396.820 1821.960 397.080 ;
      LAYER met2 ;
        RECT 1510.870 510.410 1511.150 514.000 ;
        RECT 1510.340 510.270 1511.150 510.410 ;
        RECT 1510.340 397.110 1510.480 510.270 ;
        RECT 1510.870 510.000 1511.150 510.270 ;
        RECT 1510.280 396.790 1510.540 397.110 ;
        RECT 1821.700 396.790 1821.960 397.110 ;
        RECT 1821.760 16.730 1821.900 396.790 ;
        RECT 1821.760 16.590 1822.820 16.730 ;
        RECT 1822.680 2.400 1822.820 16.590 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1527.270 496.980 1527.590 497.040 ;
        RECT 1531.410 496.980 1531.730 497.040 ;
        RECT 1527.270 496.840 1531.730 496.980 ;
        RECT 1527.270 496.780 1527.590 496.840 ;
        RECT 1531.410 496.780 1531.730 496.840 ;
        RECT 1531.410 286.520 1531.730 286.580 ;
        RECT 1835.470 286.520 1835.790 286.580 ;
        RECT 1531.410 286.380 1835.790 286.520 ;
        RECT 1531.410 286.320 1531.730 286.380 ;
        RECT 1835.470 286.320 1835.790 286.380 ;
      LAYER via ;
        RECT 1527.300 496.780 1527.560 497.040 ;
        RECT 1531.440 496.780 1531.700 497.040 ;
        RECT 1531.440 286.320 1531.700 286.580 ;
        RECT 1835.500 286.320 1835.760 286.580 ;
      LAYER met2 ;
        RECT 1527.430 510.340 1527.710 514.000 ;
        RECT 1527.360 510.000 1527.710 510.340 ;
        RECT 1527.360 497.070 1527.500 510.000 ;
        RECT 1527.300 496.750 1527.560 497.070 ;
        RECT 1531.440 496.750 1531.700 497.070 ;
        RECT 1531.500 286.610 1531.640 496.750 ;
        RECT 1531.440 286.290 1531.700 286.610 ;
        RECT 1835.500 286.290 1835.760 286.610 ;
        RECT 1835.560 16.730 1835.700 286.290 ;
        RECT 1835.560 16.590 1840.300 16.730 ;
        RECT 1840.160 2.400 1840.300 16.590 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1856.245 282.965 1856.415 331.075 ;
        RECT 1856.245 186.405 1856.415 234.515 ;
        RECT 1856.245 89.845 1856.415 137.955 ;
      LAYER mcon ;
        RECT 1856.245 330.905 1856.415 331.075 ;
        RECT 1856.245 234.345 1856.415 234.515 ;
        RECT 1856.245 137.785 1856.415 137.955 ;
      LAYER met1 ;
        RECT 1545.210 362.340 1545.530 362.400 ;
        RECT 1856.170 362.340 1856.490 362.400 ;
        RECT 1545.210 362.200 1856.490 362.340 ;
        RECT 1545.210 362.140 1545.530 362.200 ;
        RECT 1856.170 362.140 1856.490 362.200 ;
        RECT 1856.170 331.060 1856.490 331.120 ;
        RECT 1855.975 330.920 1856.490 331.060 ;
        RECT 1856.170 330.860 1856.490 330.920 ;
        RECT 1856.170 283.120 1856.490 283.180 ;
        RECT 1855.975 282.980 1856.490 283.120 ;
        RECT 1856.170 282.920 1856.490 282.980 ;
        RECT 1856.170 234.500 1856.490 234.560 ;
        RECT 1855.975 234.360 1856.490 234.500 ;
        RECT 1856.170 234.300 1856.490 234.360 ;
        RECT 1856.170 186.560 1856.490 186.620 ;
        RECT 1855.975 186.420 1856.490 186.560 ;
        RECT 1856.170 186.360 1856.490 186.420 ;
        RECT 1856.170 137.940 1856.490 138.000 ;
        RECT 1855.975 137.800 1856.490 137.940 ;
        RECT 1856.170 137.740 1856.490 137.800 ;
        RECT 1856.170 90.000 1856.490 90.060 ;
        RECT 1855.975 89.860 1856.490 90.000 ;
        RECT 1856.170 89.800 1856.490 89.860 ;
        RECT 1856.170 62.260 1856.490 62.520 ;
        RECT 1856.260 61.780 1856.400 62.260 ;
        RECT 1858.010 61.780 1858.330 61.840 ;
        RECT 1856.260 61.640 1858.330 61.780 ;
        RECT 1858.010 61.580 1858.330 61.640 ;
      LAYER via ;
        RECT 1545.240 362.140 1545.500 362.400 ;
        RECT 1856.200 362.140 1856.460 362.400 ;
        RECT 1856.200 330.860 1856.460 331.120 ;
        RECT 1856.200 282.920 1856.460 283.180 ;
        RECT 1856.200 234.300 1856.460 234.560 ;
        RECT 1856.200 186.360 1856.460 186.620 ;
        RECT 1856.200 137.740 1856.460 138.000 ;
        RECT 1856.200 89.800 1856.460 90.060 ;
        RECT 1856.200 62.260 1856.460 62.520 ;
        RECT 1858.040 61.580 1858.300 61.840 ;
      LAYER met2 ;
        RECT 1543.530 510.410 1543.810 514.000 ;
        RECT 1543.530 510.270 1545.440 510.410 ;
        RECT 1543.530 510.000 1543.810 510.270 ;
        RECT 1545.300 362.430 1545.440 510.270 ;
        RECT 1545.240 362.110 1545.500 362.430 ;
        RECT 1856.200 362.110 1856.460 362.430 ;
        RECT 1856.260 331.150 1856.400 362.110 ;
        RECT 1856.200 330.830 1856.460 331.150 ;
        RECT 1856.200 282.890 1856.460 283.210 ;
        RECT 1856.260 234.590 1856.400 282.890 ;
        RECT 1856.200 234.270 1856.460 234.590 ;
        RECT 1856.200 186.330 1856.460 186.650 ;
        RECT 1856.260 138.030 1856.400 186.330 ;
        RECT 1856.200 137.710 1856.460 138.030 ;
        RECT 1856.200 89.770 1856.460 90.090 ;
        RECT 1856.260 62.550 1856.400 89.770 ;
        RECT 1856.200 62.230 1856.460 62.550 ;
        RECT 1858.040 61.550 1858.300 61.870 ;
        RECT 1858.100 2.400 1858.240 61.550 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.930 496.980 1560.250 497.040 ;
        RECT 1565.450 496.980 1565.770 497.040 ;
        RECT 1559.930 496.840 1565.770 496.980 ;
        RECT 1559.930 496.780 1560.250 496.840 ;
        RECT 1565.450 496.780 1565.770 496.840 ;
        RECT 1565.450 369.140 1565.770 369.200 ;
        RECT 1869.970 369.140 1870.290 369.200 ;
        RECT 1565.450 369.000 1870.290 369.140 ;
        RECT 1565.450 368.940 1565.770 369.000 ;
        RECT 1869.970 368.940 1870.290 369.000 ;
        RECT 1869.970 37.980 1870.290 38.040 ;
        RECT 1875.950 37.980 1876.270 38.040 ;
        RECT 1869.970 37.840 1876.270 37.980 ;
        RECT 1869.970 37.780 1870.290 37.840 ;
        RECT 1875.950 37.780 1876.270 37.840 ;
      LAYER via ;
        RECT 1559.960 496.780 1560.220 497.040 ;
        RECT 1565.480 496.780 1565.740 497.040 ;
        RECT 1565.480 368.940 1565.740 369.200 ;
        RECT 1870.000 368.940 1870.260 369.200 ;
        RECT 1870.000 37.780 1870.260 38.040 ;
        RECT 1875.980 37.780 1876.240 38.040 ;
      LAYER met2 ;
        RECT 1560.090 510.340 1560.370 514.000 ;
        RECT 1560.020 510.000 1560.370 510.340 ;
        RECT 1560.020 497.070 1560.160 510.000 ;
        RECT 1559.960 496.750 1560.220 497.070 ;
        RECT 1565.480 496.750 1565.740 497.070 ;
        RECT 1565.540 369.230 1565.680 496.750 ;
        RECT 1565.480 368.910 1565.740 369.230 ;
        RECT 1870.000 368.910 1870.260 369.230 ;
        RECT 1870.060 38.070 1870.200 368.910 ;
        RECT 1870.000 37.750 1870.260 38.070 ;
        RECT 1875.980 37.750 1876.240 38.070 ;
        RECT 1876.040 2.400 1876.180 37.750 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 503.440 532.150 503.500 ;
        RECT 537.810 503.440 538.130 503.500 ;
        RECT 531.830 503.300 538.130 503.440 ;
        RECT 531.830 503.240 532.150 503.300 ;
        RECT 537.810 503.240 538.130 503.300 ;
        RECT 537.810 18.260 538.130 18.320 ;
        RECT 752.170 18.260 752.490 18.320 ;
        RECT 537.810 18.120 752.490 18.260 ;
        RECT 537.810 18.060 538.130 18.120 ;
        RECT 752.170 18.060 752.490 18.120 ;
      LAYER via ;
        RECT 531.860 503.240 532.120 503.500 ;
        RECT 537.840 503.240 538.100 503.500 ;
        RECT 537.840 18.060 538.100 18.320 ;
        RECT 752.200 18.060 752.460 18.320 ;
      LAYER met2 ;
        RECT 531.990 510.340 532.270 514.000 ;
        RECT 531.920 510.000 532.270 510.340 ;
        RECT 531.920 503.530 532.060 510.000 ;
        RECT 531.860 503.210 532.120 503.530 ;
        RECT 537.840 503.210 538.100 503.530 ;
        RECT 537.900 18.350 538.040 503.210 ;
        RECT 537.840 18.030 538.100 18.350 ;
        RECT 752.200 18.030 752.460 18.350 ;
        RECT 752.260 2.400 752.400 18.030 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1890.745 338.385 1890.915 386.155 ;
        RECT 1890.745 289.765 1890.915 337.875 ;
        RECT 1890.745 241.485 1890.915 289.255 ;
        RECT 1890.745 145.265 1890.915 193.035 ;
        RECT 1890.745 48.365 1890.915 96.475 ;
      LAYER mcon ;
        RECT 1890.745 385.985 1890.915 386.155 ;
        RECT 1890.745 337.705 1890.915 337.875 ;
        RECT 1890.745 289.085 1890.915 289.255 ;
        RECT 1890.745 192.865 1890.915 193.035 ;
        RECT 1890.745 96.305 1890.915 96.475 ;
      LAYER met1 ;
        RECT 1576.030 496.980 1576.350 497.040 ;
        RECT 1579.710 496.980 1580.030 497.040 ;
        RECT 1576.030 496.840 1580.030 496.980 ;
        RECT 1576.030 496.780 1576.350 496.840 ;
        RECT 1579.710 496.780 1580.030 496.840 ;
        RECT 1579.710 403.820 1580.030 403.880 ;
        RECT 1891.130 403.820 1891.450 403.880 ;
        RECT 1579.710 403.680 1891.450 403.820 ;
        RECT 1579.710 403.620 1580.030 403.680 ;
        RECT 1891.130 403.620 1891.450 403.680 ;
        RECT 1890.670 386.140 1890.990 386.200 ;
        RECT 1890.475 386.000 1890.990 386.140 ;
        RECT 1890.670 385.940 1890.990 386.000 ;
        RECT 1890.670 338.540 1890.990 338.600 ;
        RECT 1890.475 338.400 1890.990 338.540 ;
        RECT 1890.670 338.340 1890.990 338.400 ;
        RECT 1890.670 337.860 1890.990 337.920 ;
        RECT 1890.475 337.720 1890.990 337.860 ;
        RECT 1890.670 337.660 1890.990 337.720 ;
        RECT 1890.670 289.920 1890.990 289.980 ;
        RECT 1890.475 289.780 1890.990 289.920 ;
        RECT 1890.670 289.720 1890.990 289.780 ;
        RECT 1890.670 289.240 1890.990 289.300 ;
        RECT 1890.475 289.100 1890.990 289.240 ;
        RECT 1890.670 289.040 1890.990 289.100 ;
        RECT 1890.670 241.640 1890.990 241.700 ;
        RECT 1890.475 241.500 1890.990 241.640 ;
        RECT 1890.670 241.440 1890.990 241.500 ;
        RECT 1890.670 193.020 1890.990 193.080 ;
        RECT 1890.475 192.880 1890.990 193.020 ;
        RECT 1890.670 192.820 1890.990 192.880 ;
        RECT 1890.670 145.420 1890.990 145.480 ;
        RECT 1890.475 145.280 1890.990 145.420 ;
        RECT 1890.670 145.220 1890.990 145.280 ;
        RECT 1890.670 144.740 1890.990 144.800 ;
        RECT 1891.130 144.740 1891.450 144.800 ;
        RECT 1890.670 144.600 1891.450 144.740 ;
        RECT 1890.670 144.540 1890.990 144.600 ;
        RECT 1891.130 144.540 1891.450 144.600 ;
        RECT 1890.670 96.460 1890.990 96.520 ;
        RECT 1890.475 96.320 1890.990 96.460 ;
        RECT 1890.670 96.260 1890.990 96.320 ;
        RECT 1890.685 48.520 1890.975 48.565 ;
        RECT 1893.890 48.520 1894.210 48.580 ;
        RECT 1890.685 48.380 1894.210 48.520 ;
        RECT 1890.685 48.335 1890.975 48.380 ;
        RECT 1893.890 48.320 1894.210 48.380 ;
      LAYER via ;
        RECT 1576.060 496.780 1576.320 497.040 ;
        RECT 1579.740 496.780 1580.000 497.040 ;
        RECT 1579.740 403.620 1580.000 403.880 ;
        RECT 1891.160 403.620 1891.420 403.880 ;
        RECT 1890.700 385.940 1890.960 386.200 ;
        RECT 1890.700 338.340 1890.960 338.600 ;
        RECT 1890.700 337.660 1890.960 337.920 ;
        RECT 1890.700 289.720 1890.960 289.980 ;
        RECT 1890.700 289.040 1890.960 289.300 ;
        RECT 1890.700 241.440 1890.960 241.700 ;
        RECT 1890.700 192.820 1890.960 193.080 ;
        RECT 1890.700 145.220 1890.960 145.480 ;
        RECT 1890.700 144.540 1890.960 144.800 ;
        RECT 1891.160 144.540 1891.420 144.800 ;
        RECT 1890.700 96.260 1890.960 96.520 ;
        RECT 1893.920 48.320 1894.180 48.580 ;
      LAYER met2 ;
        RECT 1576.190 510.340 1576.470 514.000 ;
        RECT 1576.120 510.000 1576.470 510.340 ;
        RECT 1576.120 497.070 1576.260 510.000 ;
        RECT 1576.060 496.750 1576.320 497.070 ;
        RECT 1579.740 496.750 1580.000 497.070 ;
        RECT 1579.800 403.910 1579.940 496.750 ;
        RECT 1579.740 403.590 1580.000 403.910 ;
        RECT 1891.160 403.590 1891.420 403.910 ;
        RECT 1891.220 386.650 1891.360 403.590 ;
        RECT 1890.760 386.510 1891.360 386.650 ;
        RECT 1890.760 386.230 1890.900 386.510 ;
        RECT 1890.700 385.910 1890.960 386.230 ;
        RECT 1890.700 338.310 1890.960 338.630 ;
        RECT 1890.760 337.950 1890.900 338.310 ;
        RECT 1890.700 337.630 1890.960 337.950 ;
        RECT 1890.700 289.690 1890.960 290.010 ;
        RECT 1890.760 289.330 1890.900 289.690 ;
        RECT 1890.700 289.010 1890.960 289.330 ;
        RECT 1890.700 241.410 1890.960 241.730 ;
        RECT 1890.760 194.210 1890.900 241.410 ;
        RECT 1890.760 194.070 1891.360 194.210 ;
        RECT 1891.220 193.530 1891.360 194.070 ;
        RECT 1890.760 193.390 1891.360 193.530 ;
        RECT 1890.760 193.110 1890.900 193.390 ;
        RECT 1890.700 192.790 1890.960 193.110 ;
        RECT 1890.700 145.190 1890.960 145.510 ;
        RECT 1890.760 144.830 1890.900 145.190 ;
        RECT 1890.700 144.510 1890.960 144.830 ;
        RECT 1891.160 144.510 1891.420 144.830 ;
        RECT 1891.220 96.970 1891.360 144.510 ;
        RECT 1890.760 96.830 1891.360 96.970 ;
        RECT 1890.760 96.550 1890.900 96.830 ;
        RECT 1890.700 96.230 1890.960 96.550 ;
        RECT 1893.920 48.290 1894.180 48.610 ;
        RECT 1893.980 2.400 1894.120 48.290 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 375.940 1593.830 376.000 ;
        RECT 1911.370 375.940 1911.690 376.000 ;
        RECT 1593.510 375.800 1911.690 375.940 ;
        RECT 1593.510 375.740 1593.830 375.800 ;
        RECT 1911.370 375.740 1911.690 375.800 ;
      LAYER via ;
        RECT 1593.540 375.740 1593.800 376.000 ;
        RECT 1911.400 375.740 1911.660 376.000 ;
      LAYER met2 ;
        RECT 1592.750 510.410 1593.030 514.000 ;
        RECT 1592.750 510.270 1593.740 510.410 ;
        RECT 1592.750 510.000 1593.030 510.270 ;
        RECT 1593.600 376.030 1593.740 510.270 ;
        RECT 1593.540 375.710 1593.800 376.030 ;
        RECT 1911.400 375.710 1911.660 376.030 ;
        RECT 1911.460 17.410 1911.600 375.710 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1608.690 503.440 1609.010 503.500 ;
        RECT 1613.750 503.440 1614.070 503.500 ;
        RECT 1608.690 503.300 1614.070 503.440 ;
        RECT 1608.690 503.240 1609.010 503.300 ;
        RECT 1613.750 503.240 1614.070 503.300 ;
        RECT 1613.750 417.420 1614.070 417.480 ;
        RECT 1925.170 417.420 1925.490 417.480 ;
        RECT 1613.750 417.280 1925.490 417.420 ;
        RECT 1613.750 417.220 1614.070 417.280 ;
        RECT 1925.170 417.220 1925.490 417.280 ;
      LAYER via ;
        RECT 1608.720 503.240 1608.980 503.500 ;
        RECT 1613.780 503.240 1614.040 503.500 ;
        RECT 1613.780 417.220 1614.040 417.480 ;
        RECT 1925.200 417.220 1925.460 417.480 ;
      LAYER met2 ;
        RECT 1608.850 510.340 1609.130 514.000 ;
        RECT 1608.780 510.000 1609.130 510.340 ;
        RECT 1608.780 503.530 1608.920 510.000 ;
        RECT 1608.720 503.210 1608.980 503.530 ;
        RECT 1613.780 503.210 1614.040 503.530 ;
        RECT 1613.840 417.510 1613.980 503.210 ;
        RECT 1613.780 417.190 1614.040 417.510 ;
        RECT 1925.200 417.190 1925.460 417.510 ;
        RECT 1925.260 16.730 1925.400 417.190 ;
        RECT 1925.260 16.590 1929.540 16.730 ;
        RECT 1929.400 2.400 1929.540 16.590 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1625.250 500.380 1625.570 500.440 ;
        RECT 1686.890 500.380 1687.210 500.440 ;
        RECT 1625.250 500.240 1687.210 500.380 ;
        RECT 1625.250 500.180 1625.570 500.240 ;
        RECT 1686.890 500.180 1687.210 500.240 ;
        RECT 1686.890 168.880 1687.210 168.940 ;
        RECT 1945.870 168.880 1946.190 168.940 ;
        RECT 1686.890 168.740 1946.190 168.880 ;
        RECT 1686.890 168.680 1687.210 168.740 ;
        RECT 1945.870 168.680 1946.190 168.740 ;
        RECT 1945.870 96.460 1946.190 96.520 ;
        RECT 1946.790 96.460 1947.110 96.520 ;
        RECT 1945.870 96.320 1947.110 96.460 ;
        RECT 1945.870 96.260 1946.190 96.320 ;
        RECT 1946.790 96.260 1947.110 96.320 ;
        RECT 1947.250 47.980 1947.570 48.240 ;
        RECT 1947.340 47.560 1947.480 47.980 ;
        RECT 1947.250 47.300 1947.570 47.560 ;
      LAYER via ;
        RECT 1625.280 500.180 1625.540 500.440 ;
        RECT 1686.920 500.180 1687.180 500.440 ;
        RECT 1686.920 168.680 1687.180 168.940 ;
        RECT 1945.900 168.680 1946.160 168.940 ;
        RECT 1945.900 96.260 1946.160 96.520 ;
        RECT 1946.820 96.260 1947.080 96.520 ;
        RECT 1947.280 47.980 1947.540 48.240 ;
        RECT 1947.280 47.300 1947.540 47.560 ;
      LAYER met2 ;
        RECT 1625.410 510.340 1625.690 514.000 ;
        RECT 1625.340 510.000 1625.690 510.340 ;
        RECT 1625.340 500.470 1625.480 510.000 ;
        RECT 1625.280 500.150 1625.540 500.470 ;
        RECT 1686.920 500.150 1687.180 500.470 ;
        RECT 1686.980 168.970 1687.120 500.150 ;
        RECT 1686.920 168.650 1687.180 168.970 ;
        RECT 1945.900 168.650 1946.160 168.970 ;
        RECT 1945.960 96.550 1946.100 168.650 ;
        RECT 1945.900 96.230 1946.160 96.550 ;
        RECT 1946.820 96.230 1947.080 96.550 ;
        RECT 1946.880 48.690 1947.020 96.230 ;
        RECT 1946.880 48.550 1947.480 48.690 ;
        RECT 1947.340 48.270 1947.480 48.550 ;
        RECT 1947.280 47.950 1947.540 48.270 ;
        RECT 1947.280 47.270 1947.540 47.590 ;
        RECT 1947.340 2.400 1947.480 47.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.810 410.620 1642.130 410.680 ;
        RECT 1959.670 410.620 1959.990 410.680 ;
        RECT 1641.810 410.480 1959.990 410.620 ;
        RECT 1641.810 410.420 1642.130 410.480 ;
        RECT 1959.670 410.420 1959.990 410.480 ;
        RECT 1959.670 62.120 1959.990 62.180 ;
        RECT 1965.190 62.120 1965.510 62.180 ;
        RECT 1959.670 61.980 1965.510 62.120 ;
        RECT 1959.670 61.920 1959.990 61.980 ;
        RECT 1965.190 61.920 1965.510 61.980 ;
      LAYER via ;
        RECT 1641.840 410.420 1642.100 410.680 ;
        RECT 1959.700 410.420 1959.960 410.680 ;
        RECT 1959.700 61.920 1959.960 62.180 ;
        RECT 1965.220 61.920 1965.480 62.180 ;
      LAYER met2 ;
        RECT 1641.510 511.090 1641.790 514.000 ;
        RECT 1640.520 510.950 1641.790 511.090 ;
        RECT 1640.520 483.325 1640.660 510.950 ;
        RECT 1641.510 510.000 1641.790 510.950 ;
        RECT 1640.450 482.955 1640.730 483.325 ;
        RECT 1641.830 482.955 1642.110 483.325 ;
        RECT 1641.900 410.710 1642.040 482.955 ;
        RECT 1641.840 410.390 1642.100 410.710 ;
        RECT 1959.700 410.390 1959.960 410.710 ;
        RECT 1959.760 62.210 1959.900 410.390 ;
        RECT 1959.700 61.890 1959.960 62.210 ;
        RECT 1965.220 61.890 1965.480 62.210 ;
        RECT 1965.280 2.400 1965.420 61.890 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 1640.450 483.000 1640.730 483.280 ;
        RECT 1641.830 483.000 1642.110 483.280 ;
      LAYER met3 ;
        RECT 1640.425 483.290 1640.755 483.305 ;
        RECT 1641.805 483.290 1642.135 483.305 ;
        RECT 1640.425 482.990 1642.135 483.290 ;
        RECT 1640.425 482.975 1640.755 482.990 ;
        RECT 1641.805 482.975 1642.135 482.990 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1657.910 503.440 1658.230 503.500 ;
        RECT 1662.510 503.440 1662.830 503.500 ;
        RECT 1657.910 503.300 1662.830 503.440 ;
        RECT 1657.910 503.240 1658.230 503.300 ;
        RECT 1662.510 503.240 1662.830 503.300 ;
        RECT 1662.510 341.600 1662.830 341.660 ;
        RECT 1980.370 341.600 1980.690 341.660 ;
        RECT 1662.510 341.460 1980.690 341.600 ;
        RECT 1662.510 341.400 1662.830 341.460 ;
        RECT 1980.370 341.400 1980.690 341.460 ;
        RECT 1980.370 62.120 1980.690 62.180 ;
        RECT 1983.130 62.120 1983.450 62.180 ;
        RECT 1980.370 61.980 1983.450 62.120 ;
        RECT 1980.370 61.920 1980.690 61.980 ;
        RECT 1983.130 61.920 1983.450 61.980 ;
      LAYER via ;
        RECT 1657.940 503.240 1658.200 503.500 ;
        RECT 1662.540 503.240 1662.800 503.500 ;
        RECT 1662.540 341.400 1662.800 341.660 ;
        RECT 1980.400 341.400 1980.660 341.660 ;
        RECT 1980.400 61.920 1980.660 62.180 ;
        RECT 1983.160 61.920 1983.420 62.180 ;
      LAYER met2 ;
        RECT 1658.070 510.340 1658.350 514.000 ;
        RECT 1658.000 510.000 1658.350 510.340 ;
        RECT 1658.000 503.530 1658.140 510.000 ;
        RECT 1657.940 503.210 1658.200 503.530 ;
        RECT 1662.540 503.210 1662.800 503.530 ;
        RECT 1662.600 341.690 1662.740 503.210 ;
        RECT 1662.540 341.370 1662.800 341.690 ;
        RECT 1980.400 341.370 1980.660 341.690 ;
        RECT 1980.460 62.210 1980.600 341.370 ;
        RECT 1980.400 61.890 1980.660 62.210 ;
        RECT 1983.160 61.890 1983.420 62.210 ;
        RECT 1983.220 2.400 1983.360 61.890 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.310 355.200 1676.630 355.260 ;
        RECT 2001.070 355.200 2001.390 355.260 ;
        RECT 1676.310 355.060 2001.390 355.200 ;
        RECT 1676.310 355.000 1676.630 355.060 ;
        RECT 2001.070 355.000 2001.390 355.060 ;
      LAYER via ;
        RECT 1676.340 355.000 1676.600 355.260 ;
        RECT 2001.100 355.000 2001.360 355.260 ;
      LAYER met2 ;
        RECT 1674.170 510.410 1674.450 514.000 ;
        RECT 1674.170 510.270 1676.540 510.410 ;
        RECT 1674.170 510.000 1674.450 510.270 ;
        RECT 1676.400 355.290 1676.540 510.270 ;
        RECT 1676.340 354.970 1676.600 355.290 ;
        RECT 2001.100 354.970 2001.360 355.290 ;
        RECT 2001.160 2.400 2001.300 354.970 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.570 503.440 1690.890 503.500 ;
        RECT 1696.550 503.440 1696.870 503.500 ;
        RECT 1690.570 503.300 1696.870 503.440 ;
        RECT 1690.570 503.240 1690.890 503.300 ;
        RECT 1696.550 503.240 1696.870 503.300 ;
        RECT 1696.550 424.220 1696.870 424.280 ;
        RECT 2014.870 424.220 2015.190 424.280 ;
        RECT 1696.550 424.080 2015.190 424.220 ;
        RECT 1696.550 424.020 1696.870 424.080 ;
        RECT 2014.870 424.020 2015.190 424.080 ;
      LAYER via ;
        RECT 1690.600 503.240 1690.860 503.500 ;
        RECT 1696.580 503.240 1696.840 503.500 ;
        RECT 1696.580 424.020 1696.840 424.280 ;
        RECT 2014.900 424.020 2015.160 424.280 ;
      LAYER met2 ;
        RECT 1690.730 510.340 1691.010 514.000 ;
        RECT 1690.660 510.000 1691.010 510.340 ;
        RECT 1690.660 503.530 1690.800 510.000 ;
        RECT 1690.600 503.210 1690.860 503.530 ;
        RECT 1696.580 503.210 1696.840 503.530 ;
        RECT 1696.640 424.310 1696.780 503.210 ;
        RECT 1696.580 423.990 1696.840 424.310 ;
        RECT 2014.900 423.990 2015.160 424.310 ;
        RECT 2014.960 17.410 2015.100 423.990 ;
        RECT 2014.960 17.270 2018.780 17.410 ;
        RECT 2018.640 2.400 2018.780 17.270 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1706.670 496.980 1706.990 497.040 ;
        RECT 1710.810 496.980 1711.130 497.040 ;
        RECT 1706.670 496.840 1711.130 496.980 ;
        RECT 1706.670 496.780 1706.990 496.840 ;
        RECT 1710.810 496.780 1711.130 496.840 ;
        RECT 1710.810 431.360 1711.130 431.420 ;
        RECT 2035.570 431.360 2035.890 431.420 ;
        RECT 1710.810 431.220 2035.890 431.360 ;
        RECT 1710.810 431.160 1711.130 431.220 ;
        RECT 2035.570 431.160 2035.890 431.220 ;
      LAYER via ;
        RECT 1706.700 496.780 1706.960 497.040 ;
        RECT 1710.840 496.780 1711.100 497.040 ;
        RECT 1710.840 431.160 1711.100 431.420 ;
        RECT 2035.600 431.160 2035.860 431.420 ;
      LAYER met2 ;
        RECT 1706.830 510.340 1707.110 514.000 ;
        RECT 1706.760 510.000 1707.110 510.340 ;
        RECT 1706.760 497.070 1706.900 510.000 ;
        RECT 1706.700 496.750 1706.960 497.070 ;
        RECT 1710.840 496.750 1711.100 497.070 ;
        RECT 1710.900 431.450 1711.040 496.750 ;
        RECT 1710.840 431.130 1711.100 431.450 ;
        RECT 2035.600 431.130 2035.860 431.450 ;
        RECT 2035.660 17.410 2035.800 431.130 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 51.580 1724.930 51.640 ;
        RECT 2053.970 51.580 2054.290 51.640 ;
        RECT 1724.610 51.440 2054.290 51.580 ;
        RECT 1724.610 51.380 1724.930 51.440 ;
        RECT 2053.970 51.380 2054.290 51.440 ;
      LAYER via ;
        RECT 1724.640 51.380 1724.900 51.640 ;
        RECT 2054.000 51.380 2054.260 51.640 ;
      LAYER met2 ;
        RECT 1723.390 510.410 1723.670 514.000 ;
        RECT 1723.390 510.270 1724.840 510.410 ;
        RECT 1723.390 510.000 1723.670 510.270 ;
        RECT 1724.700 51.670 1724.840 510.270 ;
        RECT 1724.640 51.350 1724.900 51.670 ;
        RECT 2054.000 51.350 2054.260 51.670 ;
        RECT 2054.060 20.810 2054.200 51.350 ;
        RECT 2054.060 20.670 2054.660 20.810 ;
        RECT 2054.520 2.400 2054.660 20.670 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 17.920 551.930 17.980 ;
        RECT 769.650 17.920 769.970 17.980 ;
        RECT 551.610 17.780 769.970 17.920 ;
        RECT 551.610 17.720 551.930 17.780 ;
        RECT 769.650 17.720 769.970 17.780 ;
      LAYER via ;
        RECT 551.640 17.720 551.900 17.980 ;
        RECT 769.680 17.720 769.940 17.980 ;
      LAYER met2 ;
        RECT 548.090 510.410 548.370 514.000 ;
        RECT 548.090 510.270 551.840 510.410 ;
        RECT 548.090 510.000 548.370 510.270 ;
        RECT 551.700 18.010 551.840 510.270 ;
        RECT 551.640 17.690 551.900 18.010 ;
        RECT 769.680 17.690 769.940 18.010 ;
        RECT 769.740 2.400 769.880 17.690 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 496.980 1739.650 497.040 ;
        RECT 1744.850 496.980 1745.170 497.040 ;
        RECT 1739.330 496.840 1745.170 496.980 ;
        RECT 1739.330 496.780 1739.650 496.840 ;
        RECT 1744.850 496.780 1745.170 496.840 ;
        RECT 1744.850 210.700 1745.170 210.760 ;
        RECT 2070.070 210.700 2070.390 210.760 ;
        RECT 1744.850 210.560 2070.390 210.700 ;
        RECT 1744.850 210.500 1745.170 210.560 ;
        RECT 2070.070 210.500 2070.390 210.560 ;
        RECT 2070.070 96.460 2070.390 96.520 ;
        RECT 2072.370 96.460 2072.690 96.520 ;
        RECT 2070.070 96.320 2072.690 96.460 ;
        RECT 2070.070 96.260 2070.390 96.320 ;
        RECT 2072.370 96.260 2072.690 96.320 ;
      LAYER via ;
        RECT 1739.360 496.780 1739.620 497.040 ;
        RECT 1744.880 496.780 1745.140 497.040 ;
        RECT 1744.880 210.500 1745.140 210.760 ;
        RECT 2070.100 210.500 2070.360 210.760 ;
        RECT 2070.100 96.260 2070.360 96.520 ;
        RECT 2072.400 96.260 2072.660 96.520 ;
      LAYER met2 ;
        RECT 1739.490 510.340 1739.770 514.000 ;
        RECT 1739.420 510.000 1739.770 510.340 ;
        RECT 1739.420 497.070 1739.560 510.000 ;
        RECT 1739.360 496.750 1739.620 497.070 ;
        RECT 1744.880 496.750 1745.140 497.070 ;
        RECT 1744.940 210.790 1745.080 496.750 ;
        RECT 1744.880 210.470 1745.140 210.790 ;
        RECT 2070.100 210.470 2070.360 210.790 ;
        RECT 2070.160 96.550 2070.300 210.470 ;
        RECT 2070.100 96.230 2070.360 96.550 ;
        RECT 2072.400 96.230 2072.660 96.550 ;
        RECT 2072.460 2.400 2072.600 96.230 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 438.160 1759.430 438.220 ;
        RECT 2083.870 438.160 2084.190 438.220 ;
        RECT 1759.110 438.020 2084.190 438.160 ;
        RECT 1759.110 437.960 1759.430 438.020 ;
        RECT 2083.870 437.960 2084.190 438.020 ;
        RECT 2083.870 37.980 2084.190 38.040 ;
        RECT 2089.850 37.980 2090.170 38.040 ;
        RECT 2083.870 37.840 2090.170 37.980 ;
        RECT 2083.870 37.780 2084.190 37.840 ;
        RECT 2089.850 37.780 2090.170 37.840 ;
      LAYER via ;
        RECT 1759.140 437.960 1759.400 438.220 ;
        RECT 2083.900 437.960 2084.160 438.220 ;
        RECT 2083.900 37.780 2084.160 38.040 ;
        RECT 2089.880 37.780 2090.140 38.040 ;
      LAYER met2 ;
        RECT 1756.050 510.410 1756.330 514.000 ;
        RECT 1756.050 510.270 1759.340 510.410 ;
        RECT 1756.050 510.000 1756.330 510.270 ;
        RECT 1759.200 438.250 1759.340 510.270 ;
        RECT 1759.140 437.930 1759.400 438.250 ;
        RECT 2083.900 437.930 2084.160 438.250 ;
        RECT 2083.960 38.070 2084.100 437.930 ;
        RECT 2083.900 37.750 2084.160 38.070 ;
        RECT 2089.880 37.750 2090.140 38.070 ;
        RECT 2089.940 2.400 2090.080 37.750 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 458.900 1773.230 458.960 ;
        RECT 2104.570 458.900 2104.890 458.960 ;
        RECT 1772.910 458.760 2104.890 458.900 ;
        RECT 1772.910 458.700 1773.230 458.760 ;
        RECT 2104.570 458.700 2104.890 458.760 ;
      LAYER via ;
        RECT 1772.940 458.700 1773.200 458.960 ;
        RECT 2104.600 458.700 2104.860 458.960 ;
      LAYER met2 ;
        RECT 1772.150 510.410 1772.430 514.000 ;
        RECT 1772.150 510.270 1773.140 510.410 ;
        RECT 1772.150 510.000 1772.430 510.270 ;
        RECT 1773.000 458.990 1773.140 510.270 ;
        RECT 1772.940 458.670 1773.200 458.990 ;
        RECT 2104.600 458.670 2104.860 458.990 ;
        RECT 2104.660 17.410 2104.800 458.670 ;
        RECT 2104.660 17.270 2108.020 17.410 ;
        RECT 2107.880 2.400 2108.020 17.270 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1788.550 496.980 1788.870 497.040 ;
        RECT 1793.150 496.980 1793.470 497.040 ;
        RECT 1788.550 496.840 1793.470 496.980 ;
        RECT 1788.550 496.780 1788.870 496.840 ;
        RECT 1793.150 496.780 1793.470 496.840 ;
        RECT 1793.150 382.740 1793.470 382.800 ;
        RECT 2125.270 382.740 2125.590 382.800 ;
        RECT 1793.150 382.600 2125.590 382.740 ;
        RECT 1793.150 382.540 1793.470 382.600 ;
        RECT 2125.270 382.540 2125.590 382.600 ;
      LAYER via ;
        RECT 1788.580 496.780 1788.840 497.040 ;
        RECT 1793.180 496.780 1793.440 497.040 ;
        RECT 1793.180 382.540 1793.440 382.800 ;
        RECT 2125.300 382.540 2125.560 382.800 ;
      LAYER met2 ;
        RECT 1788.710 510.340 1788.990 514.000 ;
        RECT 1788.640 510.000 1788.990 510.340 ;
        RECT 1788.640 497.070 1788.780 510.000 ;
        RECT 1788.580 496.750 1788.840 497.070 ;
        RECT 1793.180 496.750 1793.440 497.070 ;
        RECT 1793.240 382.830 1793.380 496.750 ;
        RECT 1793.180 382.510 1793.440 382.830 ;
        RECT 2125.300 382.510 2125.560 382.830 ;
        RECT 2125.360 17.410 2125.500 382.510 ;
        RECT 2125.360 17.270 2125.960 17.410 ;
        RECT 2125.820 2.400 2125.960 17.270 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.410 389.880 1807.730 389.940 ;
        RECT 2139.070 389.880 2139.390 389.940 ;
        RECT 1807.410 389.740 2139.390 389.880 ;
        RECT 1807.410 389.680 1807.730 389.740 ;
        RECT 2139.070 389.680 2139.390 389.740 ;
      LAYER via ;
        RECT 1807.440 389.680 1807.700 389.940 ;
        RECT 2139.100 389.680 2139.360 389.940 ;
      LAYER met2 ;
        RECT 1804.810 510.410 1805.090 514.000 ;
        RECT 1804.810 510.270 1807.640 510.410 ;
        RECT 1804.810 510.000 1805.090 510.270 ;
        RECT 1807.500 389.970 1807.640 510.270 ;
        RECT 1807.440 389.650 1807.700 389.970 ;
        RECT 2139.100 389.650 2139.360 389.970 ;
        RECT 2139.160 17.410 2139.300 389.650 ;
        RECT 2139.160 17.270 2143.900 17.410 ;
        RECT 2143.760 2.400 2143.900 17.270 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 396.680 1821.530 396.740 ;
        RECT 2159.770 396.680 2160.090 396.740 ;
        RECT 1821.210 396.540 2160.090 396.680 ;
        RECT 1821.210 396.480 1821.530 396.540 ;
        RECT 2159.770 396.480 2160.090 396.540 ;
      LAYER via ;
        RECT 1821.240 396.480 1821.500 396.740 ;
        RECT 2159.800 396.480 2160.060 396.740 ;
      LAYER met2 ;
        RECT 1821.370 510.340 1821.650 514.000 ;
        RECT 1821.300 510.000 1821.650 510.340 ;
        RECT 1821.300 396.770 1821.440 510.000 ;
        RECT 1821.240 396.450 1821.500 396.770 ;
        RECT 2159.800 396.450 2160.060 396.770 ;
        RECT 2159.860 17.410 2160.000 396.450 ;
        RECT 2159.860 17.270 2161.840 17.410 ;
        RECT 2161.700 2.400 2161.840 17.270 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1837.310 496.980 1837.630 497.040 ;
        RECT 1841.910 496.980 1842.230 497.040 ;
        RECT 1837.310 496.840 1842.230 496.980 ;
        RECT 1837.310 496.780 1837.630 496.840 ;
        RECT 1841.910 496.780 1842.230 496.840 ;
        RECT 1841.910 465.700 1842.230 465.760 ;
        RECT 2173.570 465.700 2173.890 465.760 ;
        RECT 1841.910 465.560 2173.890 465.700 ;
        RECT 1841.910 465.500 1842.230 465.560 ;
        RECT 2173.570 465.500 2173.890 465.560 ;
      LAYER via ;
        RECT 1837.340 496.780 1837.600 497.040 ;
        RECT 1841.940 496.780 1842.200 497.040 ;
        RECT 1841.940 465.500 1842.200 465.760 ;
        RECT 2173.600 465.500 2173.860 465.760 ;
      LAYER met2 ;
        RECT 1837.470 510.340 1837.750 514.000 ;
        RECT 1837.400 510.000 1837.750 510.340 ;
        RECT 1837.400 497.070 1837.540 510.000 ;
        RECT 1837.340 496.750 1837.600 497.070 ;
        RECT 1841.940 496.750 1842.200 497.070 ;
        RECT 1842.000 465.790 1842.140 496.750 ;
        RECT 1841.940 465.470 1842.200 465.790 ;
        RECT 2173.600 465.470 2173.860 465.790 ;
        RECT 2173.660 17.410 2173.800 465.470 ;
        RECT 2173.660 17.270 2179.320 17.410 ;
        RECT 2179.180 2.400 2179.320 17.270 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1853.870 479.640 1854.190 479.700 ;
        RECT 2194.270 479.640 2194.590 479.700 ;
        RECT 1853.870 479.500 2194.590 479.640 ;
        RECT 1853.870 479.440 1854.190 479.500 ;
        RECT 2194.270 479.440 2194.590 479.500 ;
      LAYER via ;
        RECT 1853.900 479.440 1854.160 479.700 ;
        RECT 2194.300 479.440 2194.560 479.700 ;
      LAYER met2 ;
        RECT 1854.030 510.340 1854.310 514.000 ;
        RECT 1853.960 510.000 1854.310 510.340 ;
        RECT 1853.960 479.730 1854.100 510.000 ;
        RECT 1853.900 479.410 1854.160 479.730 ;
        RECT 2194.300 479.410 2194.560 479.730 ;
        RECT 2194.360 17.410 2194.500 479.410 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.970 496.980 1870.290 497.040 ;
        RECT 1875.950 496.980 1876.270 497.040 ;
        RECT 1869.970 496.840 1876.270 496.980 ;
        RECT 1869.970 496.780 1870.290 496.840 ;
        RECT 1875.950 496.780 1876.270 496.840 ;
        RECT 1875.950 403.480 1876.270 403.540 ;
        RECT 2214.970 403.480 2215.290 403.540 ;
        RECT 1875.950 403.340 2215.290 403.480 ;
        RECT 1875.950 403.280 1876.270 403.340 ;
        RECT 2214.970 403.280 2215.290 403.340 ;
      LAYER via ;
        RECT 1870.000 496.780 1870.260 497.040 ;
        RECT 1875.980 496.780 1876.240 497.040 ;
        RECT 1875.980 403.280 1876.240 403.540 ;
        RECT 2215.000 403.280 2215.260 403.540 ;
      LAYER met2 ;
        RECT 1870.130 510.340 1870.410 514.000 ;
        RECT 1870.060 510.000 1870.410 510.340 ;
        RECT 1870.060 497.070 1870.200 510.000 ;
        RECT 1870.000 496.750 1870.260 497.070 ;
        RECT 1875.980 496.750 1876.240 497.070 ;
        RECT 1876.040 403.570 1876.180 496.750 ;
        RECT 1875.980 403.250 1876.240 403.570 ;
        RECT 2215.000 403.250 2215.260 403.570 ;
        RECT 2215.060 2.400 2215.200 403.250 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1886.070 496.980 1886.390 497.040 ;
        RECT 1890.210 496.980 1890.530 497.040 ;
        RECT 1886.070 496.840 1890.530 496.980 ;
        RECT 1886.070 496.780 1886.390 496.840 ;
        RECT 1890.210 496.780 1890.530 496.840 ;
        RECT 1890.210 20.300 1890.530 20.360 ;
        RECT 2232.910 20.300 2233.230 20.360 ;
        RECT 1890.210 20.160 2233.230 20.300 ;
        RECT 1890.210 20.100 1890.530 20.160 ;
        RECT 2232.910 20.100 2233.230 20.160 ;
      LAYER via ;
        RECT 1886.100 496.780 1886.360 497.040 ;
        RECT 1890.240 496.780 1890.500 497.040 ;
        RECT 1890.240 20.100 1890.500 20.360 ;
        RECT 2232.940 20.100 2233.200 20.360 ;
      LAYER met2 ;
        RECT 1886.230 510.340 1886.510 514.000 ;
        RECT 1886.160 510.000 1886.510 510.340 ;
        RECT 1886.160 497.070 1886.300 510.000 ;
        RECT 1886.100 496.750 1886.360 497.070 ;
        RECT 1890.240 496.750 1890.500 497.070 ;
        RECT 1890.300 20.390 1890.440 496.750 ;
        RECT 1890.240 20.070 1890.500 20.390 ;
        RECT 2232.940 20.070 2233.200 20.390 ;
        RECT 2233.000 2.400 2233.140 20.070 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 17.240 565.730 17.300 ;
        RECT 787.590 17.240 787.910 17.300 ;
        RECT 565.410 17.100 787.910 17.240 ;
        RECT 565.410 17.040 565.730 17.100 ;
        RECT 787.590 17.040 787.910 17.100 ;
      LAYER via ;
        RECT 565.440 17.040 565.700 17.300 ;
        RECT 787.620 17.040 787.880 17.300 ;
      LAYER met2 ;
        RECT 564.650 510.410 564.930 514.000 ;
        RECT 564.650 510.270 565.640 510.410 ;
        RECT 564.650 510.000 564.930 510.270 ;
        RECT 565.500 17.330 565.640 510.270 ;
        RECT 565.440 17.010 565.700 17.330 ;
        RECT 787.620 17.010 787.880 17.330 ;
        RECT 787.680 2.400 787.820 17.010 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 18.940 1904.330 19.000 ;
        RECT 2250.850 18.940 2251.170 19.000 ;
        RECT 1904.010 18.800 2251.170 18.940 ;
        RECT 1904.010 18.740 1904.330 18.800 ;
        RECT 2250.850 18.740 2251.170 18.800 ;
      LAYER via ;
        RECT 1904.040 18.740 1904.300 19.000 ;
        RECT 2250.880 18.740 2251.140 19.000 ;
      LAYER met2 ;
        RECT 1902.790 510.410 1903.070 514.000 ;
        RECT 1902.790 510.270 1904.240 510.410 ;
        RECT 1902.790 510.000 1903.070 510.270 ;
        RECT 1904.100 19.030 1904.240 510.270 ;
        RECT 1904.040 18.710 1904.300 19.030 ;
        RECT 2250.880 18.710 2251.140 19.030 ;
        RECT 2250.940 2.400 2251.080 18.710 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1918.730 496.980 1919.050 497.040 ;
        RECT 1924.710 496.980 1925.030 497.040 ;
        RECT 1918.730 496.840 1925.030 496.980 ;
        RECT 1918.730 496.780 1919.050 496.840 ;
        RECT 1924.710 496.780 1925.030 496.840 ;
        RECT 1924.710 20.640 1925.030 20.700 ;
        RECT 2268.330 20.640 2268.650 20.700 ;
        RECT 1924.710 20.500 2268.650 20.640 ;
        RECT 1924.710 20.440 1925.030 20.500 ;
        RECT 2268.330 20.440 2268.650 20.500 ;
      LAYER via ;
        RECT 1918.760 496.780 1919.020 497.040 ;
        RECT 1924.740 496.780 1925.000 497.040 ;
        RECT 1924.740 20.440 1925.000 20.700 ;
        RECT 2268.360 20.440 2268.620 20.700 ;
      LAYER met2 ;
        RECT 1918.890 510.340 1919.170 514.000 ;
        RECT 1918.820 510.000 1919.170 510.340 ;
        RECT 1918.820 497.070 1918.960 510.000 ;
        RECT 1918.760 496.750 1919.020 497.070 ;
        RECT 1924.740 496.750 1925.000 497.070 ;
        RECT 1924.800 20.730 1924.940 496.750 ;
        RECT 1924.740 20.410 1925.000 20.730 ;
        RECT 2268.360 20.410 2268.620 20.730 ;
        RECT 2268.420 2.400 2268.560 20.410 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 19.280 1938.830 19.340 ;
        RECT 2286.270 19.280 2286.590 19.340 ;
        RECT 1938.510 19.140 2286.590 19.280 ;
        RECT 1938.510 19.080 1938.830 19.140 ;
        RECT 2286.270 19.080 2286.590 19.140 ;
      LAYER via ;
        RECT 1938.540 19.080 1938.800 19.340 ;
        RECT 2286.300 19.080 2286.560 19.340 ;
      LAYER met2 ;
        RECT 1935.450 510.410 1935.730 514.000 ;
        RECT 1935.450 510.270 1938.740 510.410 ;
        RECT 1935.450 510.000 1935.730 510.270 ;
        RECT 1938.600 19.370 1938.740 510.270 ;
        RECT 1938.540 19.050 1938.800 19.370 ;
        RECT 2286.300 19.050 2286.560 19.370 ;
        RECT 2286.360 2.400 2286.500 19.050 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 19.620 1952.630 19.680 ;
        RECT 2304.210 19.620 2304.530 19.680 ;
        RECT 1952.310 19.480 2304.530 19.620 ;
        RECT 1952.310 19.420 1952.630 19.480 ;
        RECT 2304.210 19.420 2304.530 19.480 ;
      LAYER via ;
        RECT 1952.340 19.420 1952.600 19.680 ;
        RECT 2304.240 19.420 2304.500 19.680 ;
      LAYER met2 ;
        RECT 1951.550 510.410 1951.830 514.000 ;
        RECT 1951.550 510.270 1952.540 510.410 ;
        RECT 1951.550 510.000 1951.830 510.270 ;
        RECT 1952.400 19.710 1952.540 510.270 ;
        RECT 1952.340 19.390 1952.600 19.710 ;
        RECT 2304.240 19.390 2304.500 19.710 ;
        RECT 2304.300 2.400 2304.440 19.390 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.950 498.680 1968.270 498.740 ;
        RECT 1973.010 498.680 1973.330 498.740 ;
        RECT 1967.950 498.540 1973.330 498.680 ;
        RECT 1967.950 498.480 1968.270 498.540 ;
        RECT 1973.010 498.480 1973.330 498.540 ;
        RECT 1973.010 19.960 1973.330 20.020 ;
        RECT 2322.150 19.960 2322.470 20.020 ;
        RECT 1973.010 19.820 2322.470 19.960 ;
        RECT 1973.010 19.760 1973.330 19.820 ;
        RECT 2322.150 19.760 2322.470 19.820 ;
      LAYER via ;
        RECT 1967.980 498.480 1968.240 498.740 ;
        RECT 1973.040 498.480 1973.300 498.740 ;
        RECT 1973.040 19.760 1973.300 20.020 ;
        RECT 2322.180 19.760 2322.440 20.020 ;
      LAYER met2 ;
        RECT 1968.110 510.340 1968.390 514.000 ;
        RECT 1968.040 510.000 1968.390 510.340 ;
        RECT 1968.040 498.770 1968.180 510.000 ;
        RECT 1967.980 498.450 1968.240 498.770 ;
        RECT 1973.040 498.450 1973.300 498.770 ;
        RECT 1973.100 20.050 1973.240 498.450 ;
        RECT 1973.040 19.730 1973.300 20.050 ;
        RECT 2322.180 19.730 2322.440 20.050 ;
        RECT 2322.240 2.400 2322.380 19.730 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.810 18.600 1987.130 18.660 ;
        RECT 2339.170 18.600 2339.490 18.660 ;
        RECT 1986.810 18.460 2339.490 18.600 ;
        RECT 1986.810 18.400 1987.130 18.460 ;
        RECT 2339.170 18.400 2339.490 18.460 ;
      LAYER via ;
        RECT 1986.840 18.400 1987.100 18.660 ;
        RECT 2339.200 18.400 2339.460 18.660 ;
      LAYER met2 ;
        RECT 1984.210 510.410 1984.490 514.000 ;
        RECT 1984.210 510.270 1987.040 510.410 ;
        RECT 1984.210 510.000 1984.490 510.270 ;
        RECT 1986.900 18.690 1987.040 510.270 ;
        RECT 1986.840 18.370 1987.100 18.690 ;
        RECT 2339.200 18.370 2339.460 18.690 ;
        RECT 2339.260 16.050 2339.400 18.370 ;
        RECT 2339.260 15.910 2339.860 16.050 ;
        RECT 2339.720 2.400 2339.860 15.910 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.610 17.920 2000.930 17.980 ;
        RECT 2357.570 17.920 2357.890 17.980 ;
        RECT 2000.610 17.780 2357.890 17.920 ;
        RECT 2000.610 17.720 2000.930 17.780 ;
        RECT 2357.570 17.720 2357.890 17.780 ;
      LAYER via ;
        RECT 2000.640 17.720 2000.900 17.980 ;
        RECT 2357.600 17.720 2357.860 17.980 ;
      LAYER met2 ;
        RECT 2000.770 510.340 2001.050 514.000 ;
        RECT 2000.700 510.000 2001.050 510.340 ;
        RECT 2000.700 18.010 2000.840 510.000 ;
        RECT 2000.640 17.690 2000.900 18.010 ;
        RECT 2357.600 17.690 2357.860 18.010 ;
        RECT 2357.660 2.400 2357.800 17.690 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.710 496.980 2017.030 497.040 ;
        RECT 2021.310 496.980 2021.630 497.040 ;
        RECT 2016.710 496.840 2021.630 496.980 ;
        RECT 2016.710 496.780 2017.030 496.840 ;
        RECT 2021.310 496.780 2021.630 496.840 ;
        RECT 2021.310 18.260 2021.630 18.320 ;
        RECT 2375.510 18.260 2375.830 18.320 ;
        RECT 2021.310 18.120 2375.830 18.260 ;
        RECT 2021.310 18.060 2021.630 18.120 ;
        RECT 2375.510 18.060 2375.830 18.120 ;
      LAYER via ;
        RECT 2016.740 496.780 2017.000 497.040 ;
        RECT 2021.340 496.780 2021.600 497.040 ;
        RECT 2021.340 18.060 2021.600 18.320 ;
        RECT 2375.540 18.060 2375.800 18.320 ;
      LAYER met2 ;
        RECT 2016.870 510.340 2017.150 514.000 ;
        RECT 2016.800 510.000 2017.150 510.340 ;
        RECT 2016.800 497.070 2016.940 510.000 ;
        RECT 2016.740 496.750 2017.000 497.070 ;
        RECT 2021.340 496.750 2021.600 497.070 ;
        RECT 2021.400 18.350 2021.540 496.750 ;
        RECT 2021.340 18.030 2021.600 18.350 ;
        RECT 2375.540 18.030 2375.800 18.350 ;
        RECT 2375.600 2.400 2375.740 18.030 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2035.110 17.240 2035.430 17.300 ;
        RECT 2393.450 17.240 2393.770 17.300 ;
        RECT 2035.110 17.100 2393.770 17.240 ;
        RECT 2035.110 17.040 2035.430 17.100 ;
        RECT 2393.450 17.040 2393.770 17.100 ;
      LAYER via ;
        RECT 2035.140 17.040 2035.400 17.300 ;
        RECT 2393.480 17.040 2393.740 17.300 ;
      LAYER met2 ;
        RECT 2033.430 510.410 2033.710 514.000 ;
        RECT 2033.430 510.270 2035.340 510.410 ;
        RECT 2033.430 510.000 2033.710 510.270 ;
        RECT 2035.200 17.330 2035.340 510.270 ;
        RECT 2035.140 17.010 2035.400 17.330 ;
        RECT 2393.480 17.010 2393.740 17.330 ;
        RECT 2393.540 2.400 2393.680 17.010 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2049.370 499.020 2049.690 499.080 ;
        RECT 2055.810 499.020 2056.130 499.080 ;
        RECT 2049.370 498.880 2056.130 499.020 ;
        RECT 2049.370 498.820 2049.690 498.880 ;
        RECT 2055.810 498.820 2056.130 498.880 ;
        RECT 2055.810 17.580 2056.130 17.640 ;
        RECT 2411.390 17.580 2411.710 17.640 ;
        RECT 2055.810 17.440 2411.710 17.580 ;
        RECT 2055.810 17.380 2056.130 17.440 ;
        RECT 2411.390 17.380 2411.710 17.440 ;
      LAYER via ;
        RECT 2049.400 498.820 2049.660 499.080 ;
        RECT 2055.840 498.820 2056.100 499.080 ;
        RECT 2055.840 17.380 2056.100 17.640 ;
        RECT 2411.420 17.380 2411.680 17.640 ;
      LAYER met2 ;
        RECT 2049.530 510.340 2049.810 514.000 ;
        RECT 2049.460 510.000 2049.810 510.340 ;
        RECT 2049.460 499.110 2049.600 510.000 ;
        RECT 2049.400 498.790 2049.660 499.110 ;
        RECT 2055.840 498.790 2056.100 499.110 ;
        RECT 2055.900 17.670 2056.040 498.790 ;
        RECT 2055.840 17.350 2056.100 17.670 ;
        RECT 2411.420 17.350 2411.680 17.670 ;
        RECT 2411.480 2.400 2411.620 17.350 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.590 496.980 580.910 497.040 ;
        RECT 586.110 496.980 586.430 497.040 ;
        RECT 580.590 496.840 586.430 496.980 ;
        RECT 580.590 496.780 580.910 496.840 ;
        RECT 586.110 496.780 586.430 496.840 ;
        RECT 586.110 17.580 586.430 17.640 ;
        RECT 586.110 17.440 788.280 17.580 ;
        RECT 586.110 17.380 586.430 17.440 ;
        RECT 788.140 17.240 788.280 17.440 ;
        RECT 805.530 17.240 805.850 17.300 ;
        RECT 788.140 17.100 805.850 17.240 ;
        RECT 805.530 17.040 805.850 17.100 ;
      LAYER via ;
        RECT 580.620 496.780 580.880 497.040 ;
        RECT 586.140 496.780 586.400 497.040 ;
        RECT 586.140 17.380 586.400 17.640 ;
        RECT 805.560 17.040 805.820 17.300 ;
      LAYER met2 ;
        RECT 580.750 510.340 581.030 514.000 ;
        RECT 580.680 510.000 581.030 510.340 ;
        RECT 580.680 497.070 580.820 510.000 ;
        RECT 580.620 496.750 580.880 497.070 ;
        RECT 586.140 496.750 586.400 497.070 ;
        RECT 586.200 17.670 586.340 496.750 ;
        RECT 586.140 17.350 586.400 17.670 ;
        RECT 805.560 17.010 805.820 17.330 ;
        RECT 805.620 2.400 805.760 17.010 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 407.170 17.580 407.490 17.640 ;
        RECT 2.830 17.440 407.490 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 407.170 17.380 407.490 17.440 ;
      LAYER via ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 407.200 17.380 407.460 17.640 ;
      LAYER met2 ;
        RECT 412.390 510.410 412.670 514.000 ;
        RECT 407.260 510.270 412.670 510.410 ;
        RECT 407.260 17.670 407.400 510.270 ;
        RECT 412.390 510.000 412.670 510.270 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 407.200 17.350 407.460 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.240 8.670 17.300 ;
        RECT 414.070 17.240 414.390 17.300 ;
        RECT 8.350 17.100 414.390 17.240 ;
        RECT 8.350 17.040 8.670 17.100 ;
        RECT 414.070 17.040 414.390 17.100 ;
      LAYER via ;
        RECT 8.380 17.040 8.640 17.300 ;
        RECT 414.100 17.040 414.360 17.300 ;
      LAYER met2 ;
        RECT 417.450 510.410 417.730 514.000 ;
        RECT 414.160 510.270 417.730 510.410 ;
        RECT 414.160 17.330 414.300 510.270 ;
        RECT 417.450 510.000 417.730 510.270 ;
        RECT 8.380 17.010 8.640 17.330 ;
        RECT 414.100 17.010 414.360 17.330 ;
        RECT 8.440 2.400 8.580 17.010 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 3010.000 547.020 3528.900 ;
        RECT 724.020 3010.000 727.020 3528.900 ;
        RECT 904.020 3010.000 907.020 3528.900 ;
        RECT 1084.020 3010.000 1087.020 3528.900 ;
        RECT 1264.020 3010.000 1267.020 3528.900 ;
        RECT 1444.020 3010.000 1447.020 3528.900 ;
        RECT 1624.020 3010.000 1627.020 3528.900 ;
        RECT 1804.020 3010.000 1807.020 3528.900 ;
        RECT 1984.020 3010.000 1987.020 3528.900 ;
        RECT 2164.020 3010.000 2167.020 3528.900 ;
        RECT 2344.020 3010.000 2347.020 3528.900 ;
        RECT 544.020 -9.220 547.020 510.000 ;
        RECT 724.020 -9.220 727.020 510.000 ;
        RECT 904.020 -9.220 907.020 510.000 ;
        RECT 1084.020 -9.220 1087.020 510.000 ;
        RECT 1264.020 -9.220 1267.020 510.000 ;
        RECT 1444.020 -9.220 1447.020 510.000 ;
        RECT 1624.020 -9.220 1627.020 510.000 ;
        RECT 1804.020 -9.220 1807.020 510.000 ;
        RECT 1984.020 -9.220 1987.020 510.000 ;
        RECT 2164.020 -9.220 2167.020 510.000 ;
        RECT 2344.020 -9.220 2347.020 510.000 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3010.000 457.020 3528.900 ;
        RECT 634.020 3010.000 637.020 3528.900 ;
        RECT 814.020 3010.000 817.020 3528.900 ;
        RECT 994.020 3010.000 997.020 3528.900 ;
        RECT 1174.020 3010.000 1177.020 3528.900 ;
        RECT 1354.020 3010.000 1357.020 3528.900 ;
        RECT 1534.020 3010.000 1537.020 3528.900 ;
        RECT 1714.020 3010.000 1717.020 3528.900 ;
        RECT 1894.020 3010.000 1897.020 3528.900 ;
        RECT 2074.020 3010.000 2077.020 3528.900 ;
        RECT 2254.020 3010.000 2257.020 3528.900 ;
        RECT 2434.020 3010.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 510.000 ;
        RECT 634.020 -9.220 637.020 510.000 ;
        RECT 814.020 -9.220 817.020 510.000 ;
        RECT 994.020 -9.220 997.020 510.000 ;
        RECT 1174.020 -9.220 1177.020 510.000 ;
        RECT 1354.020 -9.220 1357.020 510.000 ;
        RECT 1534.020 -9.220 1537.020 510.000 ;
        RECT 1714.020 -9.220 1717.020 510.000 ;
        RECT 1894.020 -9.220 1897.020 510.000 ;
        RECT 2074.020 -9.220 2077.020 510.000 ;
        RECT 2254.020 -9.220 2257.020 510.000 ;
        RECT 2434.020 -9.220 2437.020 510.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 3010.000 565.020 3538.100 ;
        RECT 742.020 3010.000 745.020 3538.100 ;
        RECT 922.020 3010.000 925.020 3538.100 ;
        RECT 1102.020 3010.000 1105.020 3538.100 ;
        RECT 1282.020 3010.000 1285.020 3538.100 ;
        RECT 1462.020 3010.000 1465.020 3538.100 ;
        RECT 1642.020 3010.000 1645.020 3538.100 ;
        RECT 1822.020 3010.000 1825.020 3538.100 ;
        RECT 2002.020 3010.000 2005.020 3538.100 ;
        RECT 2182.020 3010.000 2185.020 3538.100 ;
        RECT 2362.020 3010.000 2365.020 3538.100 ;
        RECT 562.020 -18.420 565.020 510.000 ;
        RECT 742.020 -18.420 745.020 510.000 ;
        RECT 922.020 -18.420 925.020 510.000 ;
        RECT 1102.020 -18.420 1105.020 510.000 ;
        RECT 1282.020 -18.420 1285.020 510.000 ;
        RECT 1462.020 -18.420 1465.020 510.000 ;
        RECT 1642.020 -18.420 1645.020 510.000 ;
        RECT 1822.020 -18.420 1825.020 510.000 ;
        RECT 2002.020 -18.420 2005.020 510.000 ;
        RECT 2182.020 -18.420 2185.020 510.000 ;
        RECT 2362.020 -18.420 2365.020 510.000 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3010.000 475.020 3538.100 ;
        RECT 652.020 3010.000 655.020 3538.100 ;
        RECT 832.020 3010.000 835.020 3538.100 ;
        RECT 1012.020 3010.000 1015.020 3538.100 ;
        RECT 1192.020 3010.000 1195.020 3538.100 ;
        RECT 1372.020 3010.000 1375.020 3538.100 ;
        RECT 1552.020 3010.000 1555.020 3538.100 ;
        RECT 1732.020 3010.000 1735.020 3538.100 ;
        RECT 1912.020 3010.000 1915.020 3538.100 ;
        RECT 2092.020 3010.000 2095.020 3538.100 ;
        RECT 2272.020 3010.000 2275.020 3538.100 ;
        RECT 2452.020 3010.000 2455.020 3538.100 ;
        RECT 472.020 -18.420 475.020 510.000 ;
        RECT 652.020 -18.420 655.020 510.000 ;
        RECT 832.020 -18.420 835.020 510.000 ;
        RECT 1012.020 -18.420 1015.020 510.000 ;
        RECT 1192.020 -18.420 1195.020 510.000 ;
        RECT 1372.020 -18.420 1375.020 510.000 ;
        RECT 1552.020 -18.420 1555.020 510.000 ;
        RECT 1732.020 -18.420 1735.020 510.000 ;
        RECT 1912.020 -18.420 1915.020 510.000 ;
        RECT 2092.020 -18.420 2095.020 510.000 ;
        RECT 2272.020 -18.420 2275.020 510.000 ;
        RECT 2452.020 -18.420 2455.020 510.000 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 3010.000 583.020 3547.300 ;
        RECT 760.020 3010.000 763.020 3547.300 ;
        RECT 940.020 3010.000 943.020 3547.300 ;
        RECT 1120.020 3010.000 1123.020 3547.300 ;
        RECT 1300.020 3010.000 1303.020 3547.300 ;
        RECT 1480.020 3010.000 1483.020 3547.300 ;
        RECT 1660.020 3010.000 1663.020 3547.300 ;
        RECT 1840.020 3010.000 1843.020 3547.300 ;
        RECT 2020.020 3010.000 2023.020 3547.300 ;
        RECT 2200.020 3010.000 2203.020 3547.300 ;
        RECT 2380.020 3010.000 2383.020 3547.300 ;
        RECT 580.020 -27.620 583.020 510.000 ;
        RECT 760.020 -27.620 763.020 510.000 ;
        RECT 940.020 -27.620 943.020 510.000 ;
        RECT 1120.020 -27.620 1123.020 510.000 ;
        RECT 1300.020 -27.620 1303.020 510.000 ;
        RECT 1480.020 -27.620 1483.020 510.000 ;
        RECT 1660.020 -27.620 1663.020 510.000 ;
        RECT 1840.020 -27.620 1843.020 510.000 ;
        RECT 2020.020 -27.620 2023.020 510.000 ;
        RECT 2200.020 -27.620 2203.020 510.000 ;
        RECT 2380.020 -27.620 2383.020 510.000 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 3010.000 493.020 3547.300 ;
        RECT 670.020 3010.000 673.020 3547.300 ;
        RECT 850.020 3010.000 853.020 3547.300 ;
        RECT 1030.020 3010.000 1033.020 3547.300 ;
        RECT 1210.020 3010.000 1213.020 3547.300 ;
        RECT 1390.020 3010.000 1393.020 3547.300 ;
        RECT 1570.020 3010.000 1573.020 3547.300 ;
        RECT 1750.020 3010.000 1753.020 3547.300 ;
        RECT 1930.020 3010.000 1933.020 3547.300 ;
        RECT 2110.020 3010.000 2113.020 3547.300 ;
        RECT 2290.020 3010.000 2293.020 3547.300 ;
        RECT 2470.020 3010.000 2473.020 3547.300 ;
        RECT 490.020 -27.620 493.020 510.000 ;
        RECT 670.020 -27.620 673.020 510.000 ;
        RECT 850.020 -27.620 853.020 510.000 ;
        RECT 1030.020 -27.620 1033.020 510.000 ;
        RECT 1210.020 -27.620 1213.020 510.000 ;
        RECT 1390.020 -27.620 1393.020 510.000 ;
        RECT 1570.020 -27.620 1573.020 510.000 ;
        RECT 1750.020 -27.620 1753.020 510.000 ;
        RECT 1930.020 -27.620 1933.020 510.000 ;
        RECT 2110.020 -27.620 2113.020 510.000 ;
        RECT 2290.020 -27.620 2293.020 510.000 ;
        RECT 2470.020 -27.620 2473.020 510.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3010.000 421.020 3556.500 ;
        RECT 598.020 3010.000 601.020 3556.500 ;
        RECT 778.020 3010.000 781.020 3556.500 ;
        RECT 958.020 3010.000 961.020 3556.500 ;
        RECT 1138.020 3010.000 1141.020 3556.500 ;
        RECT 1318.020 3010.000 1321.020 3556.500 ;
        RECT 1498.020 3010.000 1501.020 3556.500 ;
        RECT 1678.020 3010.000 1681.020 3556.500 ;
        RECT 1858.020 3010.000 1861.020 3556.500 ;
        RECT 2038.020 3010.000 2041.020 3556.500 ;
        RECT 2218.020 3010.000 2221.020 3556.500 ;
        RECT 2398.020 3010.000 2401.020 3556.500 ;
        RECT 418.020 -36.820 421.020 510.000 ;
        RECT 598.020 -36.820 601.020 510.000 ;
        RECT 778.020 -36.820 781.020 510.000 ;
        RECT 958.020 -36.820 961.020 510.000 ;
        RECT 1138.020 -36.820 1141.020 510.000 ;
        RECT 1318.020 -36.820 1321.020 510.000 ;
        RECT 1498.020 -36.820 1501.020 510.000 ;
        RECT 1678.020 -36.820 1681.020 510.000 ;
        RECT 1858.020 -36.820 1861.020 510.000 ;
        RECT 2038.020 -36.820 2041.020 510.000 ;
        RECT 2218.020 -36.820 2221.020 510.000 ;
        RECT 2398.020 -36.820 2401.020 510.000 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 3010.000 511.020 3556.500 ;
        RECT 688.020 3010.000 691.020 3556.500 ;
        RECT 868.020 3010.000 871.020 3556.500 ;
        RECT 1048.020 3010.000 1051.020 3556.500 ;
        RECT 1228.020 3010.000 1231.020 3556.500 ;
        RECT 1408.020 3010.000 1411.020 3556.500 ;
        RECT 1588.020 3010.000 1591.020 3556.500 ;
        RECT 1768.020 3010.000 1771.020 3556.500 ;
        RECT 1948.020 3010.000 1951.020 3556.500 ;
        RECT 2128.020 3010.000 2131.020 3556.500 ;
        RECT 2308.020 3010.000 2311.020 3556.500 ;
        RECT 2488.020 3010.000 2491.020 3556.500 ;
        RECT 508.020 -36.820 511.020 510.000 ;
        RECT 688.020 -36.820 691.020 510.000 ;
        RECT 868.020 -36.820 871.020 510.000 ;
        RECT 1048.020 -36.820 1051.020 510.000 ;
        RECT 1228.020 -36.820 1231.020 510.000 ;
        RECT 1408.020 -36.820 1411.020 510.000 ;
        RECT 1588.020 -36.820 1591.020 510.000 ;
        RECT 1768.020 -36.820 1771.020 510.000 ;
        RECT 1948.020 -36.820 1951.020 510.000 ;
        RECT 2128.020 -36.820 2131.020 510.000 ;
        RECT 2308.020 -36.820 2311.020 510.000 ;
        RECT 2488.020 -36.820 2491.020 510.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 415.520 520.795 2504.380 2998.885 ;
      LAYER met1 ;
        RECT 412.370 514.460 2504.380 2999.040 ;
      LAYER met2 ;
        RECT 412.400 3005.720 448.450 3006.010 ;
        RECT 449.290 3005.720 526.190 3006.010 ;
        RECT 527.030 3005.720 603.930 3006.010 ;
        RECT 604.770 3005.720 681.670 3006.010 ;
        RECT 682.510 3005.720 759.410 3006.010 ;
        RECT 760.250 3005.720 837.150 3006.010 ;
        RECT 837.990 3005.720 914.890 3006.010 ;
        RECT 915.730 3005.720 992.630 3006.010 ;
        RECT 993.470 3005.720 1070.370 3006.010 ;
        RECT 1071.210 3005.720 1148.110 3006.010 ;
        RECT 1148.950 3005.720 1225.850 3006.010 ;
        RECT 1226.690 3005.720 1303.590 3006.010 ;
        RECT 1304.430 3005.720 1381.330 3006.010 ;
        RECT 1382.170 3005.720 1459.070 3006.010 ;
        RECT 1459.910 3005.720 1537.270 3006.010 ;
        RECT 1538.110 3005.720 1615.010 3006.010 ;
        RECT 1615.850 3005.720 1692.750 3006.010 ;
        RECT 1693.590 3005.720 1770.490 3006.010 ;
        RECT 1771.330 3005.720 1848.230 3006.010 ;
        RECT 1849.070 3005.720 1925.970 3006.010 ;
        RECT 1926.810 3005.720 2003.710 3006.010 ;
        RECT 2004.550 3005.720 2081.450 3006.010 ;
        RECT 2082.290 3005.720 2159.190 3006.010 ;
        RECT 2160.030 3005.720 2236.930 3006.010 ;
        RECT 2237.770 3005.720 2314.670 3006.010 ;
        RECT 2315.510 3005.720 2392.410 3006.010 ;
        RECT 2393.250 3005.720 2470.150 3006.010 ;
        RECT 2470.990 3005.720 2501.520 3006.010 ;
        RECT 412.400 514.280 2501.520 3005.720 ;
        RECT 412.950 514.000 417.170 514.280 ;
        RECT 418.010 514.000 422.690 514.280 ;
        RECT 423.530 514.000 428.210 514.280 ;
        RECT 429.050 514.000 433.730 514.280 ;
        RECT 434.570 514.000 439.250 514.280 ;
        RECT 440.090 514.000 444.310 514.280 ;
        RECT 445.150 514.000 449.830 514.280 ;
        RECT 450.670 514.000 455.350 514.280 ;
        RECT 456.190 514.000 460.870 514.280 ;
        RECT 461.710 514.000 466.390 514.280 ;
        RECT 467.230 514.000 471.910 514.280 ;
        RECT 472.750 514.000 476.970 514.280 ;
        RECT 477.810 514.000 482.490 514.280 ;
        RECT 483.330 514.000 488.010 514.280 ;
        RECT 488.850 514.000 493.530 514.280 ;
        RECT 494.370 514.000 499.050 514.280 ;
        RECT 499.890 514.000 504.570 514.280 ;
        RECT 505.410 514.000 509.630 514.280 ;
        RECT 510.470 514.000 515.150 514.280 ;
        RECT 515.990 514.000 520.670 514.280 ;
        RECT 521.510 514.000 526.190 514.280 ;
        RECT 527.030 514.000 531.710 514.280 ;
        RECT 532.550 514.000 537.230 514.280 ;
        RECT 538.070 514.000 542.290 514.280 ;
        RECT 543.130 514.000 547.810 514.280 ;
        RECT 548.650 514.000 553.330 514.280 ;
        RECT 554.170 514.000 558.850 514.280 ;
        RECT 559.690 514.000 564.370 514.280 ;
        RECT 565.210 514.000 569.430 514.280 ;
        RECT 570.270 514.000 574.950 514.280 ;
        RECT 575.790 514.000 580.470 514.280 ;
        RECT 581.310 514.000 585.990 514.280 ;
        RECT 586.830 514.000 591.510 514.280 ;
        RECT 592.350 514.000 597.030 514.280 ;
        RECT 597.870 514.000 602.090 514.280 ;
        RECT 602.930 514.000 607.610 514.280 ;
        RECT 608.450 514.000 613.130 514.280 ;
        RECT 613.970 514.000 618.650 514.280 ;
        RECT 619.490 514.000 624.170 514.280 ;
        RECT 625.010 514.000 629.690 514.280 ;
        RECT 630.530 514.000 634.750 514.280 ;
        RECT 635.590 514.000 640.270 514.280 ;
        RECT 641.110 514.000 645.790 514.280 ;
        RECT 646.630 514.000 651.310 514.280 ;
        RECT 652.150 514.000 656.830 514.280 ;
        RECT 657.670 514.000 662.350 514.280 ;
        RECT 663.190 514.000 667.410 514.280 ;
        RECT 668.250 514.000 672.930 514.280 ;
        RECT 673.770 514.000 678.450 514.280 ;
        RECT 679.290 514.000 683.970 514.280 ;
        RECT 684.810 514.000 689.490 514.280 ;
        RECT 690.330 514.000 694.550 514.280 ;
        RECT 695.390 514.000 700.070 514.280 ;
        RECT 700.910 514.000 705.590 514.280 ;
        RECT 706.430 514.000 711.110 514.280 ;
        RECT 711.950 514.000 716.630 514.280 ;
        RECT 717.470 514.000 722.150 514.280 ;
        RECT 722.990 514.000 727.210 514.280 ;
        RECT 728.050 514.000 732.730 514.280 ;
        RECT 733.570 514.000 738.250 514.280 ;
        RECT 739.090 514.000 743.770 514.280 ;
        RECT 744.610 514.000 749.290 514.280 ;
        RECT 750.130 514.000 754.810 514.280 ;
        RECT 755.650 514.000 759.870 514.280 ;
        RECT 760.710 514.000 765.390 514.280 ;
        RECT 766.230 514.000 770.910 514.280 ;
        RECT 771.750 514.000 776.430 514.280 ;
        RECT 777.270 514.000 781.950 514.280 ;
        RECT 782.790 514.000 787.470 514.280 ;
        RECT 788.310 514.000 792.530 514.280 ;
        RECT 793.370 514.000 798.050 514.280 ;
        RECT 798.890 514.000 803.570 514.280 ;
        RECT 804.410 514.000 809.090 514.280 ;
        RECT 809.930 514.000 814.610 514.280 ;
        RECT 815.450 514.000 819.670 514.280 ;
        RECT 820.510 514.000 825.190 514.280 ;
        RECT 826.030 514.000 830.710 514.280 ;
        RECT 831.550 514.000 836.230 514.280 ;
        RECT 837.070 514.000 841.750 514.280 ;
        RECT 842.590 514.000 847.270 514.280 ;
        RECT 848.110 514.000 852.330 514.280 ;
        RECT 853.170 514.000 857.850 514.280 ;
        RECT 858.690 514.000 863.370 514.280 ;
        RECT 864.210 514.000 868.890 514.280 ;
        RECT 869.730 514.000 874.410 514.280 ;
        RECT 875.250 514.000 879.930 514.280 ;
        RECT 880.770 514.000 884.990 514.280 ;
        RECT 885.830 514.000 890.510 514.280 ;
        RECT 891.350 514.000 896.030 514.280 ;
        RECT 896.870 514.000 901.550 514.280 ;
        RECT 902.390 514.000 907.070 514.280 ;
        RECT 907.910 514.000 912.590 514.280 ;
        RECT 913.430 514.000 917.650 514.280 ;
        RECT 918.490 514.000 923.170 514.280 ;
        RECT 924.010 514.000 928.690 514.280 ;
        RECT 929.530 514.000 934.210 514.280 ;
        RECT 935.050 514.000 939.730 514.280 ;
        RECT 940.570 514.000 944.790 514.280 ;
        RECT 945.630 514.000 950.310 514.280 ;
        RECT 951.150 514.000 955.830 514.280 ;
        RECT 956.670 514.000 961.350 514.280 ;
        RECT 962.190 514.000 966.870 514.280 ;
        RECT 967.710 514.000 972.390 514.280 ;
        RECT 973.230 514.000 977.450 514.280 ;
        RECT 978.290 514.000 982.970 514.280 ;
        RECT 983.810 514.000 988.490 514.280 ;
        RECT 989.330 514.000 994.010 514.280 ;
        RECT 994.850 514.000 999.530 514.280 ;
        RECT 1000.370 514.000 1005.050 514.280 ;
        RECT 1005.890 514.000 1010.110 514.280 ;
        RECT 1010.950 514.000 1015.630 514.280 ;
        RECT 1016.470 514.000 1021.150 514.280 ;
        RECT 1021.990 514.000 1026.670 514.280 ;
        RECT 1027.510 514.000 1032.190 514.280 ;
        RECT 1033.030 514.000 1037.710 514.280 ;
        RECT 1038.550 514.000 1042.770 514.280 ;
        RECT 1043.610 514.000 1048.290 514.280 ;
        RECT 1049.130 514.000 1053.810 514.280 ;
        RECT 1054.650 514.000 1059.330 514.280 ;
        RECT 1060.170 514.000 1064.850 514.280 ;
        RECT 1065.690 514.000 1069.910 514.280 ;
        RECT 1070.750 514.000 1075.430 514.280 ;
        RECT 1076.270 514.000 1080.950 514.280 ;
        RECT 1081.790 514.000 1086.470 514.280 ;
        RECT 1087.310 514.000 1091.990 514.280 ;
        RECT 1092.830 514.000 1097.510 514.280 ;
        RECT 1098.350 514.000 1102.570 514.280 ;
        RECT 1103.410 514.000 1108.090 514.280 ;
        RECT 1108.930 514.000 1113.610 514.280 ;
        RECT 1114.450 514.000 1119.130 514.280 ;
        RECT 1119.970 514.000 1124.650 514.280 ;
        RECT 1125.490 514.000 1130.170 514.280 ;
        RECT 1131.010 514.000 1135.230 514.280 ;
        RECT 1136.070 514.000 1140.750 514.280 ;
        RECT 1141.590 514.000 1146.270 514.280 ;
        RECT 1147.110 514.000 1151.790 514.280 ;
        RECT 1152.630 514.000 1157.310 514.280 ;
        RECT 1158.150 514.000 1162.830 514.280 ;
        RECT 1163.670 514.000 1167.890 514.280 ;
        RECT 1168.730 514.000 1173.410 514.280 ;
        RECT 1174.250 514.000 1178.930 514.280 ;
        RECT 1179.770 514.000 1184.450 514.280 ;
        RECT 1185.290 514.000 1189.970 514.280 ;
        RECT 1190.810 514.000 1195.490 514.280 ;
        RECT 1196.330 514.000 1200.550 514.280 ;
        RECT 1201.390 514.000 1206.070 514.280 ;
        RECT 1206.910 514.000 1211.590 514.280 ;
        RECT 1212.430 514.000 1217.110 514.280 ;
        RECT 1217.950 514.000 1222.630 514.280 ;
        RECT 1223.470 514.000 1227.690 514.280 ;
        RECT 1228.530 514.000 1233.210 514.280 ;
        RECT 1234.050 514.000 1238.730 514.280 ;
        RECT 1239.570 514.000 1244.250 514.280 ;
        RECT 1245.090 514.000 1249.770 514.280 ;
        RECT 1250.610 514.000 1255.290 514.280 ;
        RECT 1256.130 514.000 1260.350 514.280 ;
        RECT 1261.190 514.000 1265.870 514.280 ;
        RECT 1266.710 514.000 1271.390 514.280 ;
        RECT 1272.230 514.000 1276.910 514.280 ;
        RECT 1277.750 514.000 1282.430 514.280 ;
        RECT 1283.270 514.000 1287.950 514.280 ;
        RECT 1288.790 514.000 1293.010 514.280 ;
        RECT 1293.850 514.000 1298.530 514.280 ;
        RECT 1299.370 514.000 1304.050 514.280 ;
        RECT 1304.890 514.000 1309.570 514.280 ;
        RECT 1310.410 514.000 1315.090 514.280 ;
        RECT 1315.930 514.000 1320.610 514.280 ;
        RECT 1321.450 514.000 1325.670 514.280 ;
        RECT 1326.510 514.000 1331.190 514.280 ;
        RECT 1332.030 514.000 1336.710 514.280 ;
        RECT 1337.550 514.000 1342.230 514.280 ;
        RECT 1343.070 514.000 1347.750 514.280 ;
        RECT 1348.590 514.000 1352.810 514.280 ;
        RECT 1353.650 514.000 1358.330 514.280 ;
        RECT 1359.170 514.000 1363.850 514.280 ;
        RECT 1364.690 514.000 1369.370 514.280 ;
        RECT 1370.210 514.000 1374.890 514.280 ;
        RECT 1375.730 514.000 1380.410 514.280 ;
        RECT 1381.250 514.000 1385.470 514.280 ;
        RECT 1386.310 514.000 1390.990 514.280 ;
        RECT 1391.830 514.000 1396.510 514.280 ;
        RECT 1397.350 514.000 1402.030 514.280 ;
        RECT 1402.870 514.000 1407.550 514.280 ;
        RECT 1408.390 514.000 1413.070 514.280 ;
        RECT 1413.910 514.000 1418.130 514.280 ;
        RECT 1418.970 514.000 1423.650 514.280 ;
        RECT 1424.490 514.000 1429.170 514.280 ;
        RECT 1430.010 514.000 1434.690 514.280 ;
        RECT 1435.530 514.000 1440.210 514.280 ;
        RECT 1441.050 514.000 1445.730 514.280 ;
        RECT 1446.570 514.000 1450.790 514.280 ;
        RECT 1451.630 514.000 1456.310 514.280 ;
        RECT 1457.150 514.000 1461.830 514.280 ;
        RECT 1462.670 514.000 1467.350 514.280 ;
        RECT 1468.190 514.000 1472.870 514.280 ;
        RECT 1473.710 514.000 1477.930 514.280 ;
        RECT 1478.770 514.000 1483.450 514.280 ;
        RECT 1484.290 514.000 1488.970 514.280 ;
        RECT 1489.810 514.000 1494.490 514.280 ;
        RECT 1495.330 514.000 1500.010 514.280 ;
        RECT 1500.850 514.000 1505.530 514.280 ;
        RECT 1506.370 514.000 1510.590 514.280 ;
        RECT 1511.430 514.000 1516.110 514.280 ;
        RECT 1516.950 514.000 1521.630 514.280 ;
        RECT 1522.470 514.000 1527.150 514.280 ;
        RECT 1527.990 514.000 1532.670 514.280 ;
        RECT 1533.510 514.000 1538.190 514.280 ;
        RECT 1539.030 514.000 1543.250 514.280 ;
        RECT 1544.090 514.000 1548.770 514.280 ;
        RECT 1549.610 514.000 1554.290 514.280 ;
        RECT 1555.130 514.000 1559.810 514.280 ;
        RECT 1560.650 514.000 1565.330 514.280 ;
        RECT 1566.170 514.000 1570.850 514.280 ;
        RECT 1571.690 514.000 1575.910 514.280 ;
        RECT 1576.750 514.000 1581.430 514.280 ;
        RECT 1582.270 514.000 1586.950 514.280 ;
        RECT 1587.790 514.000 1592.470 514.280 ;
        RECT 1593.310 514.000 1597.990 514.280 ;
        RECT 1598.830 514.000 1603.050 514.280 ;
        RECT 1603.890 514.000 1608.570 514.280 ;
        RECT 1609.410 514.000 1614.090 514.280 ;
        RECT 1614.930 514.000 1619.610 514.280 ;
        RECT 1620.450 514.000 1625.130 514.280 ;
        RECT 1625.970 514.000 1630.650 514.280 ;
        RECT 1631.490 514.000 1635.710 514.280 ;
        RECT 1636.550 514.000 1641.230 514.280 ;
        RECT 1642.070 514.000 1646.750 514.280 ;
        RECT 1647.590 514.000 1652.270 514.280 ;
        RECT 1653.110 514.000 1657.790 514.280 ;
        RECT 1658.630 514.000 1663.310 514.280 ;
        RECT 1664.150 514.000 1668.370 514.280 ;
        RECT 1669.210 514.000 1673.890 514.280 ;
        RECT 1674.730 514.000 1679.410 514.280 ;
        RECT 1680.250 514.000 1684.930 514.280 ;
        RECT 1685.770 514.000 1690.450 514.280 ;
        RECT 1691.290 514.000 1695.970 514.280 ;
        RECT 1696.810 514.000 1701.030 514.280 ;
        RECT 1701.870 514.000 1706.550 514.280 ;
        RECT 1707.390 514.000 1712.070 514.280 ;
        RECT 1712.910 514.000 1717.590 514.280 ;
        RECT 1718.430 514.000 1723.110 514.280 ;
        RECT 1723.950 514.000 1728.170 514.280 ;
        RECT 1729.010 514.000 1733.690 514.280 ;
        RECT 1734.530 514.000 1739.210 514.280 ;
        RECT 1740.050 514.000 1744.730 514.280 ;
        RECT 1745.570 514.000 1750.250 514.280 ;
        RECT 1751.090 514.000 1755.770 514.280 ;
        RECT 1756.610 514.000 1760.830 514.280 ;
        RECT 1761.670 514.000 1766.350 514.280 ;
        RECT 1767.190 514.000 1771.870 514.280 ;
        RECT 1772.710 514.000 1777.390 514.280 ;
        RECT 1778.230 514.000 1782.910 514.280 ;
        RECT 1783.750 514.000 1788.430 514.280 ;
        RECT 1789.270 514.000 1793.490 514.280 ;
        RECT 1794.330 514.000 1799.010 514.280 ;
        RECT 1799.850 514.000 1804.530 514.280 ;
        RECT 1805.370 514.000 1810.050 514.280 ;
        RECT 1810.890 514.000 1815.570 514.280 ;
        RECT 1816.410 514.000 1821.090 514.280 ;
        RECT 1821.930 514.000 1826.150 514.280 ;
        RECT 1826.990 514.000 1831.670 514.280 ;
        RECT 1832.510 514.000 1837.190 514.280 ;
        RECT 1838.030 514.000 1842.710 514.280 ;
        RECT 1843.550 514.000 1848.230 514.280 ;
        RECT 1849.070 514.000 1853.750 514.280 ;
        RECT 1854.590 514.000 1858.810 514.280 ;
        RECT 1859.650 514.000 1864.330 514.280 ;
        RECT 1865.170 514.000 1869.850 514.280 ;
        RECT 1870.690 514.000 1875.370 514.280 ;
        RECT 1876.210 514.000 1880.890 514.280 ;
        RECT 1881.730 514.000 1885.950 514.280 ;
        RECT 1886.790 514.000 1891.470 514.280 ;
        RECT 1892.310 514.000 1896.990 514.280 ;
        RECT 1897.830 514.000 1902.510 514.280 ;
        RECT 1903.350 514.000 1908.030 514.280 ;
        RECT 1908.870 514.000 1913.550 514.280 ;
        RECT 1914.390 514.000 1918.610 514.280 ;
        RECT 1919.450 514.000 1924.130 514.280 ;
        RECT 1924.970 514.000 1929.650 514.280 ;
        RECT 1930.490 514.000 1935.170 514.280 ;
        RECT 1936.010 514.000 1940.690 514.280 ;
        RECT 1941.530 514.000 1946.210 514.280 ;
        RECT 1947.050 514.000 1951.270 514.280 ;
        RECT 1952.110 514.000 1956.790 514.280 ;
        RECT 1957.630 514.000 1962.310 514.280 ;
        RECT 1963.150 514.000 1967.830 514.280 ;
        RECT 1968.670 514.000 1973.350 514.280 ;
        RECT 1974.190 514.000 1978.870 514.280 ;
        RECT 1979.710 514.000 1983.930 514.280 ;
        RECT 1984.770 514.000 1989.450 514.280 ;
        RECT 1990.290 514.000 1994.970 514.280 ;
        RECT 1995.810 514.000 2000.490 514.280 ;
        RECT 2001.330 514.000 2006.010 514.280 ;
        RECT 2006.850 514.000 2011.070 514.280 ;
        RECT 2011.910 514.000 2016.590 514.280 ;
        RECT 2017.430 514.000 2022.110 514.280 ;
        RECT 2022.950 514.000 2027.630 514.280 ;
        RECT 2028.470 514.000 2033.150 514.280 ;
        RECT 2033.990 514.000 2038.670 514.280 ;
        RECT 2039.510 514.000 2043.730 514.280 ;
        RECT 2044.570 514.000 2049.250 514.280 ;
        RECT 2050.090 514.000 2054.770 514.280 ;
        RECT 2055.610 514.000 2060.290 514.280 ;
        RECT 2061.130 514.000 2065.810 514.280 ;
        RECT 2066.650 514.000 2071.330 514.280 ;
        RECT 2072.170 514.000 2076.390 514.280 ;
        RECT 2077.230 514.000 2081.910 514.280 ;
        RECT 2082.750 514.000 2087.430 514.280 ;
        RECT 2088.270 514.000 2092.950 514.280 ;
        RECT 2093.790 514.000 2098.470 514.280 ;
        RECT 2099.310 514.000 2103.990 514.280 ;
        RECT 2104.830 514.000 2109.050 514.280 ;
        RECT 2109.890 514.000 2114.570 514.280 ;
        RECT 2115.410 514.000 2120.090 514.280 ;
        RECT 2120.930 514.000 2125.610 514.280 ;
        RECT 2126.450 514.000 2131.130 514.280 ;
        RECT 2131.970 514.000 2136.190 514.280 ;
        RECT 2137.030 514.000 2141.710 514.280 ;
        RECT 2142.550 514.000 2147.230 514.280 ;
        RECT 2148.070 514.000 2152.750 514.280 ;
        RECT 2153.590 514.000 2158.270 514.280 ;
        RECT 2159.110 514.000 2163.790 514.280 ;
        RECT 2164.630 514.000 2168.850 514.280 ;
        RECT 2169.690 514.000 2174.370 514.280 ;
        RECT 2175.210 514.000 2179.890 514.280 ;
        RECT 2180.730 514.000 2185.410 514.280 ;
        RECT 2186.250 514.000 2190.930 514.280 ;
        RECT 2191.770 514.000 2196.450 514.280 ;
        RECT 2197.290 514.000 2201.510 514.280 ;
        RECT 2202.350 514.000 2207.030 514.280 ;
        RECT 2207.870 514.000 2212.550 514.280 ;
        RECT 2213.390 514.000 2218.070 514.280 ;
        RECT 2218.910 514.000 2223.590 514.280 ;
        RECT 2224.430 514.000 2229.110 514.280 ;
        RECT 2229.950 514.000 2234.170 514.280 ;
        RECT 2235.010 514.000 2239.690 514.280 ;
        RECT 2240.530 514.000 2245.210 514.280 ;
        RECT 2246.050 514.000 2250.730 514.280 ;
        RECT 2251.570 514.000 2256.250 514.280 ;
        RECT 2257.090 514.000 2261.310 514.280 ;
        RECT 2262.150 514.000 2266.830 514.280 ;
        RECT 2267.670 514.000 2272.350 514.280 ;
        RECT 2273.190 514.000 2277.870 514.280 ;
        RECT 2278.710 514.000 2283.390 514.280 ;
        RECT 2284.230 514.000 2288.910 514.280 ;
        RECT 2289.750 514.000 2293.970 514.280 ;
        RECT 2294.810 514.000 2299.490 514.280 ;
        RECT 2300.330 514.000 2305.010 514.280 ;
        RECT 2305.850 514.000 2310.530 514.280 ;
        RECT 2311.370 514.000 2316.050 514.280 ;
        RECT 2316.890 514.000 2321.570 514.280 ;
        RECT 2322.410 514.000 2326.630 514.280 ;
        RECT 2327.470 514.000 2332.150 514.280 ;
        RECT 2332.990 514.000 2337.670 514.280 ;
        RECT 2338.510 514.000 2343.190 514.280 ;
        RECT 2344.030 514.000 2348.710 514.280 ;
        RECT 2349.550 514.000 2354.230 514.280 ;
        RECT 2355.070 514.000 2359.290 514.280 ;
        RECT 2360.130 514.000 2364.810 514.280 ;
        RECT 2365.650 514.000 2370.330 514.280 ;
        RECT 2371.170 514.000 2375.850 514.280 ;
        RECT 2376.690 514.000 2381.370 514.280 ;
        RECT 2382.210 514.000 2386.430 514.280 ;
        RECT 2387.270 514.000 2391.950 514.280 ;
        RECT 2392.790 514.000 2397.470 514.280 ;
        RECT 2398.310 514.000 2402.990 514.280 ;
        RECT 2403.830 514.000 2408.510 514.280 ;
        RECT 2409.350 514.000 2414.030 514.280 ;
        RECT 2414.870 514.000 2419.090 514.280 ;
        RECT 2419.930 514.000 2424.610 514.280 ;
        RECT 2425.450 514.000 2430.130 514.280 ;
        RECT 2430.970 514.000 2435.650 514.280 ;
        RECT 2436.490 514.000 2441.170 514.280 ;
        RECT 2442.010 514.000 2446.690 514.280 ;
        RECT 2447.530 514.000 2451.750 514.280 ;
        RECT 2452.590 514.000 2457.270 514.280 ;
        RECT 2458.110 514.000 2462.790 514.280 ;
        RECT 2463.630 514.000 2468.310 514.280 ;
        RECT 2469.150 514.000 2473.830 514.280 ;
        RECT 2474.670 514.000 2479.350 514.280 ;
        RECT 2480.190 514.000 2484.410 514.280 ;
        RECT 2485.250 514.000 2489.930 514.280 ;
        RECT 2490.770 514.000 2495.450 514.280 ;
        RECT 2496.290 514.000 2500.970 514.280 ;
      LAYER met3 ;
        RECT 414.000 2982.160 2506.000 2998.965 ;
        RECT 414.000 2980.760 2505.600 2982.160 ;
        RECT 414.000 2980.120 2506.000 2980.760 ;
        RECT 414.400 2978.720 2506.000 2980.120 ;
        RECT 414.000 2926.400 2506.000 2978.720 ;
        RECT 414.000 2925.000 2505.600 2926.400 ;
        RECT 414.000 2920.280 2506.000 2925.000 ;
        RECT 414.400 2918.880 2506.000 2920.280 ;
        RECT 414.000 2870.640 2506.000 2918.880 ;
        RECT 414.000 2869.240 2505.600 2870.640 ;
        RECT 414.000 2861.120 2506.000 2869.240 ;
        RECT 414.400 2859.720 2506.000 2861.120 ;
        RECT 414.000 2815.560 2506.000 2859.720 ;
        RECT 414.000 2814.160 2505.600 2815.560 ;
        RECT 414.000 2801.280 2506.000 2814.160 ;
        RECT 414.400 2799.880 2506.000 2801.280 ;
        RECT 414.000 2759.800 2506.000 2799.880 ;
        RECT 414.000 2758.400 2505.600 2759.800 ;
        RECT 414.000 2742.120 2506.000 2758.400 ;
        RECT 414.400 2740.720 2506.000 2742.120 ;
        RECT 414.000 2704.040 2506.000 2740.720 ;
        RECT 414.000 2702.640 2505.600 2704.040 ;
        RECT 414.000 2682.280 2506.000 2702.640 ;
        RECT 414.400 2680.880 2506.000 2682.280 ;
        RECT 414.000 2648.960 2506.000 2680.880 ;
        RECT 414.000 2647.560 2505.600 2648.960 ;
        RECT 414.000 2623.120 2506.000 2647.560 ;
        RECT 414.400 2621.720 2506.000 2623.120 ;
        RECT 414.000 2593.200 2506.000 2621.720 ;
        RECT 414.000 2591.800 2505.600 2593.200 ;
        RECT 414.000 2563.280 2506.000 2591.800 ;
        RECT 414.400 2561.880 2506.000 2563.280 ;
        RECT 414.000 2537.440 2506.000 2561.880 ;
        RECT 414.000 2536.040 2505.600 2537.440 ;
        RECT 414.000 2504.120 2506.000 2536.040 ;
        RECT 414.400 2502.720 2506.000 2504.120 ;
        RECT 414.000 2482.360 2506.000 2502.720 ;
        RECT 414.000 2480.960 2505.600 2482.360 ;
        RECT 414.000 2444.280 2506.000 2480.960 ;
        RECT 414.400 2442.880 2506.000 2444.280 ;
        RECT 414.000 2426.600 2506.000 2442.880 ;
        RECT 414.000 2425.200 2505.600 2426.600 ;
        RECT 414.000 2385.120 2506.000 2425.200 ;
        RECT 414.400 2383.720 2506.000 2385.120 ;
        RECT 414.000 2370.840 2506.000 2383.720 ;
        RECT 414.000 2369.440 2505.600 2370.840 ;
        RECT 414.000 2325.280 2506.000 2369.440 ;
        RECT 414.400 2323.880 2506.000 2325.280 ;
        RECT 414.000 2315.760 2506.000 2323.880 ;
        RECT 414.000 2314.360 2505.600 2315.760 ;
        RECT 414.000 2266.120 2506.000 2314.360 ;
        RECT 414.400 2264.720 2506.000 2266.120 ;
        RECT 414.000 2260.000 2506.000 2264.720 ;
        RECT 414.000 2258.600 2505.600 2260.000 ;
        RECT 414.000 2206.280 2506.000 2258.600 ;
        RECT 414.400 2204.880 2506.000 2206.280 ;
        RECT 414.000 2204.240 2506.000 2204.880 ;
        RECT 414.000 2202.840 2505.600 2204.240 ;
        RECT 414.000 2148.480 2506.000 2202.840 ;
        RECT 414.000 2147.120 2505.600 2148.480 ;
        RECT 414.400 2147.080 2505.600 2147.120 ;
        RECT 414.400 2145.720 2506.000 2147.080 ;
        RECT 414.000 2093.400 2506.000 2145.720 ;
        RECT 414.000 2092.000 2505.600 2093.400 ;
        RECT 414.000 2087.280 2506.000 2092.000 ;
        RECT 414.400 2085.880 2506.000 2087.280 ;
        RECT 414.000 2037.640 2506.000 2085.880 ;
        RECT 414.000 2036.240 2505.600 2037.640 ;
        RECT 414.000 2028.120 2506.000 2036.240 ;
        RECT 414.400 2026.720 2506.000 2028.120 ;
        RECT 414.000 1981.880 2506.000 2026.720 ;
        RECT 414.000 1980.480 2505.600 1981.880 ;
        RECT 414.000 1968.280 2506.000 1980.480 ;
        RECT 414.400 1966.880 2506.000 1968.280 ;
        RECT 414.000 1926.800 2506.000 1966.880 ;
        RECT 414.000 1925.400 2505.600 1926.800 ;
        RECT 414.000 1909.120 2506.000 1925.400 ;
        RECT 414.400 1907.720 2506.000 1909.120 ;
        RECT 414.000 1871.040 2506.000 1907.720 ;
        RECT 414.000 1869.640 2505.600 1871.040 ;
        RECT 414.000 1849.280 2506.000 1869.640 ;
        RECT 414.400 1847.880 2506.000 1849.280 ;
        RECT 414.000 1815.280 2506.000 1847.880 ;
        RECT 414.000 1813.880 2505.600 1815.280 ;
        RECT 414.000 1790.120 2506.000 1813.880 ;
        RECT 414.400 1788.720 2506.000 1790.120 ;
        RECT 414.000 1760.200 2506.000 1788.720 ;
        RECT 414.000 1758.800 2505.600 1760.200 ;
        RECT 414.000 1730.280 2506.000 1758.800 ;
        RECT 414.400 1728.880 2506.000 1730.280 ;
        RECT 414.000 1704.440 2506.000 1728.880 ;
        RECT 414.000 1703.040 2505.600 1704.440 ;
        RECT 414.000 1670.440 2506.000 1703.040 ;
        RECT 414.400 1669.040 2506.000 1670.440 ;
        RECT 414.000 1648.680 2506.000 1669.040 ;
        RECT 414.000 1647.280 2505.600 1648.680 ;
        RECT 414.000 1611.280 2506.000 1647.280 ;
        RECT 414.400 1609.880 2506.000 1611.280 ;
        RECT 414.000 1593.600 2506.000 1609.880 ;
        RECT 414.000 1592.200 2505.600 1593.600 ;
        RECT 414.000 1551.440 2506.000 1592.200 ;
        RECT 414.400 1550.040 2506.000 1551.440 ;
        RECT 414.000 1537.840 2506.000 1550.040 ;
        RECT 414.000 1536.440 2505.600 1537.840 ;
        RECT 414.000 1492.280 2506.000 1536.440 ;
        RECT 414.400 1490.880 2506.000 1492.280 ;
        RECT 414.000 1482.080 2506.000 1490.880 ;
        RECT 414.000 1480.680 2505.600 1482.080 ;
        RECT 414.000 1432.440 2506.000 1480.680 ;
        RECT 414.400 1431.040 2506.000 1432.440 ;
        RECT 414.000 1427.000 2506.000 1431.040 ;
        RECT 414.000 1425.600 2505.600 1427.000 ;
        RECT 414.000 1373.280 2506.000 1425.600 ;
        RECT 414.400 1371.880 2506.000 1373.280 ;
        RECT 414.000 1371.240 2506.000 1371.880 ;
        RECT 414.000 1369.840 2505.600 1371.240 ;
        RECT 414.000 1315.480 2506.000 1369.840 ;
        RECT 414.000 1314.080 2505.600 1315.480 ;
        RECT 414.000 1313.440 2506.000 1314.080 ;
        RECT 414.400 1312.040 2506.000 1313.440 ;
        RECT 414.000 1259.720 2506.000 1312.040 ;
        RECT 414.000 1258.320 2505.600 1259.720 ;
        RECT 414.000 1254.280 2506.000 1258.320 ;
        RECT 414.400 1252.880 2506.000 1254.280 ;
        RECT 414.000 1204.640 2506.000 1252.880 ;
        RECT 414.000 1203.240 2505.600 1204.640 ;
        RECT 414.000 1194.440 2506.000 1203.240 ;
        RECT 414.400 1193.040 2506.000 1194.440 ;
        RECT 414.000 1148.880 2506.000 1193.040 ;
        RECT 414.000 1147.480 2505.600 1148.880 ;
        RECT 414.000 1135.280 2506.000 1147.480 ;
        RECT 414.400 1133.880 2506.000 1135.280 ;
        RECT 414.000 1093.120 2506.000 1133.880 ;
        RECT 414.000 1091.720 2505.600 1093.120 ;
        RECT 414.000 1075.440 2506.000 1091.720 ;
        RECT 414.400 1074.040 2506.000 1075.440 ;
        RECT 414.000 1038.040 2506.000 1074.040 ;
        RECT 414.000 1036.640 2505.600 1038.040 ;
        RECT 414.000 1016.280 2506.000 1036.640 ;
        RECT 414.400 1014.880 2506.000 1016.280 ;
        RECT 414.000 982.280 2506.000 1014.880 ;
        RECT 414.000 980.880 2505.600 982.280 ;
        RECT 414.000 956.440 2506.000 980.880 ;
        RECT 414.400 955.040 2506.000 956.440 ;
        RECT 414.000 926.520 2506.000 955.040 ;
        RECT 414.000 925.120 2505.600 926.520 ;
        RECT 414.000 897.280 2506.000 925.120 ;
        RECT 414.400 895.880 2506.000 897.280 ;
        RECT 414.000 871.440 2506.000 895.880 ;
        RECT 414.000 870.040 2505.600 871.440 ;
        RECT 414.000 837.440 2506.000 870.040 ;
        RECT 414.400 836.040 2506.000 837.440 ;
        RECT 414.000 815.680 2506.000 836.040 ;
        RECT 414.000 814.280 2505.600 815.680 ;
        RECT 414.000 778.280 2506.000 814.280 ;
        RECT 414.400 776.880 2506.000 778.280 ;
        RECT 414.000 759.920 2506.000 776.880 ;
        RECT 414.000 758.520 2505.600 759.920 ;
        RECT 414.000 718.440 2506.000 758.520 ;
        RECT 414.400 717.040 2506.000 718.440 ;
        RECT 414.000 704.840 2506.000 717.040 ;
        RECT 414.000 703.440 2505.600 704.840 ;
        RECT 414.000 659.280 2506.000 703.440 ;
        RECT 414.400 657.880 2506.000 659.280 ;
        RECT 414.000 649.080 2506.000 657.880 ;
        RECT 414.000 647.680 2505.600 649.080 ;
        RECT 414.000 599.440 2506.000 647.680 ;
        RECT 414.400 598.040 2506.000 599.440 ;
        RECT 414.000 593.320 2506.000 598.040 ;
        RECT 414.000 591.920 2505.600 593.320 ;
        RECT 414.000 540.280 2506.000 591.920 ;
        RECT 414.400 538.880 2506.000 540.280 ;
        RECT 414.000 538.240 2506.000 538.880 ;
        RECT 414.000 536.840 2505.600 538.240 ;
        RECT 414.000 514.255 2506.000 536.840 ;
      LAYER met4 ;
        RECT 431.040 520.640 432.640 2999.040 ;
      LAYER met4 ;
        RECT 476.535 520.640 507.440 2999.040 ;
      LAYER met4 ;
        RECT 507.840 520.640 509.440 2999.040 ;
      LAYER met4 ;
        RECT 509.840 520.640 2487.065 2999.040 ;
  END
END user_project_wrapper
END LIBRARY

