magic
tech sky130A
magscale 1 2
timestamp 1607488137
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 348709 685899 348743 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 412649 683247 412683 692733
rect 218989 666587 219023 676141
rect 348709 666587 348743 676141
rect 413017 666587 413051 683077
rect 429577 666587 429611 683077
rect 542737 666587 542771 683077
rect 559297 666587 559331 683077
rect 72985 647275 73019 656829
rect 219265 647275 219299 656829
rect 348985 647275 349019 656829
rect 72801 627963 72835 637517
rect 219081 627963 219115 637517
rect 348801 627963 348835 637517
rect 172897 89675 172931 96577
rect 178141 87091 178175 96577
rect 86141 77299 86175 86921
rect 88533 77299 88567 86921
rect 110521 77299 110555 86921
rect 124229 77299 124263 86921
rect 129841 77299 129875 86921
rect 142169 77299 142203 86921
rect 31677 67643 31711 75157
rect 85773 66283 85807 67745
rect 31677 48331 31711 57885
rect 87153 56627 87187 66181
rect 88349 56627 88383 66181
rect 95525 64923 95559 74477
rect 136741 67643 136775 77197
rect 142169 70363 142203 77129
rect 154773 67643 154807 80733
rect 160201 75939 160235 85493
rect 164433 75939 164467 85493
rect 169953 75939 169987 85493
rect 172621 75939 172655 80733
rect 178141 75939 178175 85493
rect 184029 80019 184063 86921
rect 195989 77299 196023 86921
rect 200313 77299 200347 86921
rect 230857 85595 230891 86989
rect 164341 67643 164375 72437
rect 85773 47039 85807 56525
rect 110705 48331 110739 57885
rect 111901 56627 111935 66181
rect 124413 57987 124447 60809
rect 160201 57987 160235 67541
rect 183753 66283 183787 77197
rect 215401 75939 215435 85493
rect 218161 75939 218195 85493
rect 224877 75939 224911 85493
rect 226533 75939 226567 85493
rect 251465 84235 251499 93789
rect 248889 77299 248923 80121
rect 252661 77299 252695 86921
rect 258273 84235 258307 93789
rect 272073 77299 272107 80189
rect 287345 77299 287379 80189
rect 290013 77299 290047 86921
rect 310161 80019 310195 86921
rect 408233 85595 408267 95081
rect 415041 82875 415075 92429
rect 422125 82943 422159 92429
rect 468861 89675 468895 96509
rect 350181 75939 350215 80121
rect 212733 67643 212767 70465
rect 248613 67643 248647 70397
rect 124321 48331 124355 51085
rect 136833 48331 136867 57885
rect 121653 38675 121687 48229
rect 172897 46971 172931 57885
rect 178417 56627 178451 66181
rect 212733 53839 212767 66181
rect 226625 48331 226659 63937
rect 229385 48331 229419 66181
rect 283113 57987 283147 67541
rect 328009 66283 328043 75837
rect 408141 66283 408175 75837
rect 410901 70023 410935 74477
rect 147965 38675 147999 41429
rect 208501 38675 208535 48229
rect 252477 46971 252511 48433
rect 258181 46971 258215 56457
rect 260849 48331 260883 57885
rect 266461 48331 266495 57885
rect 287253 56627 287287 66181
rect 310253 59211 310287 63461
rect 321109 55267 321143 64821
rect 328009 56627 328043 66113
rect 332333 56627 332367 66181
rect 350181 63903 350215 66181
rect 356989 56627 357023 66181
rect 422033 63563 422067 81345
rect 428841 67643 428875 80733
rect 439973 67643 440007 77197
rect 468953 67643 468987 85493
rect 31677 29019 31711 38573
rect 153485 29087 153519 31773
rect 158821 29019 158855 38573
rect 112085 11883 112119 19261
rect 153301 18003 153335 27557
rect 161673 19363 161707 28917
rect 171149 19363 171183 28917
rect 176761 27659 176795 34629
rect 207029 29019 207063 38573
rect 212825 28883 212859 44081
rect 223589 37315 223623 38709
rect 224969 37315 225003 46869
rect 226625 29019 226659 38573
rect 229385 29019 229419 38573
rect 248981 37315 249015 46869
rect 260849 38743 260883 48161
rect 287253 39831 287287 48229
rect 332333 46971 332367 48365
rect 386153 48331 386187 55981
rect 310253 40715 310287 45509
rect 284493 29087 284527 38573
rect 212917 19295 212951 26197
rect 224969 19431 225003 28917
rect 229385 21403 229419 22185
rect 230673 19363 230707 22117
rect 176761 10319 176795 12461
rect 213469 9707 213503 17221
rect 220553 9707 220587 14433
rect 224969 9707 225003 19261
rect 248613 10319 248647 19261
rect 255421 18003 255455 27557
rect 271981 19363 272015 28917
rect 284493 19363 284527 28917
rect 287253 19363 287287 28917
rect 321109 27659 321143 37213
rect 260849 9707 260883 19261
rect 310253 12359 310287 27489
rect 327917 26367 327951 31705
rect 350365 31671 350399 44081
rect 390201 38675 390235 48229
rect 357081 31739 357115 37213
rect 386245 29631 386279 38573
rect 415317 35955 415351 48909
rect 426265 48331 426299 57885
rect 427829 56627 427863 57205
rect 428841 48331 428875 51833
rect 439881 48331 439915 57817
rect 431969 37315 432003 46869
rect 439881 38675 439915 41429
rect 429025 27727 429059 31841
rect 321109 18003 321143 22117
rect 328101 21947 328135 26197
rect 357173 18003 357207 27557
rect 395445 9707 395479 18581
rect 408233 18003 408267 27557
rect 408417 9707 408451 16813
rect 422309 9707 422343 27557
rect 431969 18003 432003 27557
rect 9689 3179 9723 3349
rect 22201 3315 22235 3349
rect 22051 3281 22235 3315
rect 19257 3179 19291 3281
rect 31493 595 31527 9605
rect 85773 3451 85807 9605
rect 102241 3383 102275 3553
rect 31711 3349 31861 3383
rect 151553 595 151587 9605
rect 167009 3927 167043 4097
rect 157349 3655 157383 3893
rect 224877 3315 224911 3485
rect 224969 3315 225003 3485
rect 233525 3315 233559 3417
rect 271981 3179 272015 9605
rect 321109 6171 321143 9537
rect 347697 3383 347731 3553
rect 177773 595 177807 2805
rect 358553 595 358587 9605
rect 359749 595 359783 9605
rect 406117 595 406151 9605
rect 407313 595 407347 9605
rect 414489 595 414523 9605
rect 428933 4811 428967 9605
rect 431141 595 431175 9605
rect 432337 595 432371 9605
rect 568773 3383 568807 3553
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 348709 695453 348743 695487
rect 348709 685865 348743 685899
rect 412649 692733 412683 692767
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 412649 683213 412683 683247
rect 284033 676209 284067 676243
rect 413017 683077 413051 683111
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 348709 676141 348743 676175
rect 348709 666553 348743 666587
rect 413017 666553 413051 666587
rect 429577 683077 429611 683111
rect 429577 666553 429611 666587
rect 542737 683077 542771 683111
rect 542737 666553 542771 666587
rect 559297 683077 559331 683111
rect 559297 666553 559331 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 348985 656829 349019 656863
rect 348985 647241 349019 647275
rect 72801 637517 72835 637551
rect 72801 627929 72835 627963
rect 219081 637517 219115 637551
rect 219081 627929 219115 627963
rect 348801 637517 348835 637551
rect 348801 627929 348835 627963
rect 172897 96577 172931 96611
rect 172897 89641 172931 89675
rect 178141 96577 178175 96611
rect 468861 96509 468895 96543
rect 408233 95081 408267 95115
rect 178141 87057 178175 87091
rect 251465 93789 251499 93823
rect 230857 86989 230891 87023
rect 86141 86921 86175 86955
rect 86141 77265 86175 77299
rect 88533 86921 88567 86955
rect 88533 77265 88567 77299
rect 110521 86921 110555 86955
rect 110521 77265 110555 77299
rect 124229 86921 124263 86955
rect 124229 77265 124263 77299
rect 129841 86921 129875 86955
rect 129841 77265 129875 77299
rect 142169 86921 142203 86955
rect 184029 86921 184063 86955
rect 160201 85493 160235 85527
rect 142169 77265 142203 77299
rect 154773 80733 154807 80767
rect 136741 77197 136775 77231
rect 31677 75157 31711 75191
rect 95525 74477 95559 74511
rect 31677 67609 31711 67643
rect 85773 67745 85807 67779
rect 85773 66249 85807 66283
rect 87153 66181 87187 66215
rect 31677 57885 31711 57919
rect 87153 56593 87187 56627
rect 88349 66181 88383 66215
rect 142169 77129 142203 77163
rect 142169 70329 142203 70363
rect 136741 67609 136775 67643
rect 160201 75905 160235 75939
rect 164433 85493 164467 85527
rect 164433 75905 164467 75939
rect 169953 85493 169987 85527
rect 178141 85493 178175 85527
rect 169953 75905 169987 75939
rect 172621 80733 172655 80767
rect 172621 75905 172655 75939
rect 184029 79985 184063 80019
rect 195989 86921 196023 86955
rect 195989 77265 196023 77299
rect 200313 86921 200347 86955
rect 230857 85561 230891 85595
rect 200313 77265 200347 77299
rect 215401 85493 215435 85527
rect 178141 75905 178175 75939
rect 183753 77197 183787 77231
rect 154773 67609 154807 67643
rect 164341 72437 164375 72471
rect 164341 67609 164375 67643
rect 160201 67541 160235 67575
rect 95525 64889 95559 64923
rect 111901 66181 111935 66215
rect 88349 56593 88383 56627
rect 110705 57885 110739 57919
rect 31677 48297 31711 48331
rect 85773 56525 85807 56559
rect 124413 60809 124447 60843
rect 124413 57953 124447 57987
rect 215401 75905 215435 75939
rect 218161 85493 218195 85527
rect 218161 75905 218195 75939
rect 224877 85493 224911 85527
rect 224877 75905 224911 75939
rect 226533 85493 226567 85527
rect 258273 93789 258307 93823
rect 251465 84201 251499 84235
rect 252661 86921 252695 86955
rect 248889 80121 248923 80155
rect 248889 77265 248923 77299
rect 258273 84201 258307 84235
rect 290013 86921 290047 86955
rect 252661 77265 252695 77299
rect 272073 80189 272107 80223
rect 272073 77265 272107 77299
rect 287345 80189 287379 80223
rect 287345 77265 287379 77299
rect 310161 86921 310195 86955
rect 408233 85561 408267 85595
rect 415041 92429 415075 92463
rect 422125 92429 422159 92463
rect 468861 89641 468895 89675
rect 422125 82909 422159 82943
rect 468953 85493 468987 85527
rect 415041 82841 415075 82875
rect 422033 81345 422067 81379
rect 310161 79985 310195 80019
rect 350181 80121 350215 80155
rect 290013 77265 290047 77299
rect 226533 75905 226567 75939
rect 350181 75905 350215 75939
rect 328009 75837 328043 75871
rect 212733 70465 212767 70499
rect 212733 67609 212767 67643
rect 248613 70397 248647 70431
rect 248613 67609 248647 67643
rect 183753 66249 183787 66283
rect 283113 67541 283147 67575
rect 160201 57953 160235 57987
rect 178417 66181 178451 66215
rect 111901 56593 111935 56627
rect 136833 57885 136867 57919
rect 110705 48297 110739 48331
rect 124321 51085 124355 51119
rect 124321 48297 124355 48331
rect 136833 48297 136867 48331
rect 172897 57885 172931 57919
rect 85773 47005 85807 47039
rect 121653 48229 121687 48263
rect 178417 56593 178451 56627
rect 212733 66181 212767 66215
rect 229385 66181 229419 66215
rect 212733 53805 212767 53839
rect 226625 63937 226659 63971
rect 226625 48297 226659 48331
rect 328009 66249 328043 66283
rect 408141 75837 408175 75871
rect 410901 74477 410935 74511
rect 410901 69989 410935 70023
rect 408141 66249 408175 66283
rect 283113 57953 283147 57987
rect 287253 66181 287287 66215
rect 260849 57885 260883 57919
rect 258181 56457 258215 56491
rect 229385 48297 229419 48331
rect 252477 48433 252511 48467
rect 172897 46937 172931 46971
rect 208501 48229 208535 48263
rect 121653 38641 121687 38675
rect 147965 41429 147999 41463
rect 147965 38641 147999 38675
rect 252477 46937 252511 46971
rect 260849 48297 260883 48331
rect 266461 57885 266495 57919
rect 332333 66181 332367 66215
rect 328009 66113 328043 66147
rect 321109 64821 321143 64855
rect 310253 63461 310287 63495
rect 310253 59177 310287 59211
rect 287253 56593 287287 56627
rect 328009 56593 328043 56627
rect 350181 66181 350215 66215
rect 350181 63869 350215 63903
rect 356989 66181 357023 66215
rect 332333 56593 332367 56627
rect 428841 80733 428875 80767
rect 428841 67609 428875 67643
rect 439973 77197 440007 77231
rect 439973 67609 440007 67643
rect 468953 67609 468987 67643
rect 422033 63529 422067 63563
rect 356989 56593 357023 56627
rect 426265 57885 426299 57919
rect 321109 55233 321143 55267
rect 386153 55981 386187 56015
rect 266461 48297 266495 48331
rect 332333 48365 332367 48399
rect 287253 48229 287287 48263
rect 258181 46937 258215 46971
rect 260849 48161 260883 48195
rect 224969 46869 225003 46903
rect 208501 38641 208535 38675
rect 212825 44081 212859 44115
rect 31677 38573 31711 38607
rect 158821 38573 158855 38607
rect 153485 31773 153519 31807
rect 153485 29053 153519 29087
rect 31677 28985 31711 29019
rect 207029 38573 207063 38607
rect 158821 28985 158855 29019
rect 176761 34629 176795 34663
rect 161673 28917 161707 28951
rect 153301 27557 153335 27591
rect 112085 19261 112119 19295
rect 161673 19329 161707 19363
rect 171149 28917 171183 28951
rect 207029 28985 207063 29019
rect 223589 38709 223623 38743
rect 223589 37281 223623 37315
rect 248981 46869 249015 46903
rect 224969 37281 225003 37315
rect 226625 38573 226659 38607
rect 226625 28985 226659 29019
rect 229385 38573 229419 38607
rect 386153 48297 386187 48331
rect 415317 48909 415351 48943
rect 332333 46937 332367 46971
rect 390201 48229 390235 48263
rect 310253 45509 310287 45543
rect 310253 40681 310287 40715
rect 350365 44081 350399 44115
rect 287253 39797 287287 39831
rect 260849 38709 260883 38743
rect 248981 37281 249015 37315
rect 284493 38573 284527 38607
rect 284493 29053 284527 29087
rect 321109 37213 321143 37247
rect 229385 28985 229419 29019
rect 212825 28849 212859 28883
rect 224969 28917 225003 28951
rect 176761 27625 176795 27659
rect 171149 19329 171183 19363
rect 212917 26197 212951 26231
rect 271981 28917 272015 28951
rect 255421 27557 255455 27591
rect 229385 22185 229419 22219
rect 229385 21369 229419 21403
rect 230673 22117 230707 22151
rect 224969 19397 225003 19431
rect 230673 19329 230707 19363
rect 212917 19261 212951 19295
rect 224969 19261 225003 19295
rect 153301 17969 153335 18003
rect 213469 17221 213503 17255
rect 112085 11849 112119 11883
rect 176761 12461 176795 12495
rect 176761 10285 176795 10319
rect 213469 9673 213503 9707
rect 220553 14433 220587 14467
rect 220553 9673 220587 9707
rect 248613 19261 248647 19295
rect 271981 19329 272015 19363
rect 284493 28917 284527 28951
rect 284493 19329 284527 19363
rect 287253 28917 287287 28951
rect 321109 27625 321143 27659
rect 327917 31705 327951 31739
rect 287253 19329 287287 19363
rect 310253 27489 310287 27523
rect 255421 17969 255455 18003
rect 260849 19261 260883 19295
rect 248613 10285 248647 10319
rect 224969 9673 225003 9707
rect 390201 38641 390235 38675
rect 386245 38573 386279 38607
rect 357081 37213 357115 37247
rect 357081 31705 357115 31739
rect 350365 31637 350399 31671
rect 439881 57817 439915 57851
rect 427829 57205 427863 57239
rect 427829 56593 427863 56627
rect 426265 48297 426299 48331
rect 428841 51833 428875 51867
rect 428841 48297 428875 48331
rect 439881 48297 439915 48331
rect 431969 46869 432003 46903
rect 439881 41429 439915 41463
rect 439881 38641 439915 38675
rect 431969 37281 432003 37315
rect 415317 35921 415351 35955
rect 386245 29597 386279 29631
rect 429025 31841 429059 31875
rect 429025 27693 429059 27727
rect 327917 26333 327951 26367
rect 357173 27557 357207 27591
rect 328101 26197 328135 26231
rect 321109 22117 321143 22151
rect 328101 21913 328135 21947
rect 321109 17969 321143 18003
rect 408233 27557 408267 27591
rect 357173 17969 357207 18003
rect 395445 18581 395479 18615
rect 310253 12325 310287 12359
rect 260849 9673 260883 9707
rect 408233 17969 408267 18003
rect 422309 27557 422343 27591
rect 395445 9673 395479 9707
rect 408417 16813 408451 16847
rect 408417 9673 408451 9707
rect 431969 27557 432003 27591
rect 431969 17969 432003 18003
rect 422309 9673 422343 9707
rect 31493 9605 31527 9639
rect 9689 3349 9723 3383
rect 22201 3349 22235 3383
rect 9689 3145 9723 3179
rect 19257 3281 19291 3315
rect 22017 3281 22051 3315
rect 19257 3145 19291 3179
rect 85773 9605 85807 9639
rect 151553 9605 151587 9639
rect 85773 3417 85807 3451
rect 102241 3553 102275 3587
rect 31677 3349 31711 3383
rect 31861 3349 31895 3383
rect 102241 3349 102275 3383
rect 31493 561 31527 595
rect 271981 9605 272015 9639
rect 167009 4097 167043 4131
rect 157349 3893 157383 3927
rect 167009 3893 167043 3927
rect 157349 3621 157383 3655
rect 224877 3485 224911 3519
rect 224877 3281 224911 3315
rect 224969 3485 225003 3519
rect 224969 3281 225003 3315
rect 233525 3417 233559 3451
rect 233525 3281 233559 3315
rect 358553 9605 358587 9639
rect 321109 9537 321143 9571
rect 321109 6137 321143 6171
rect 347697 3553 347731 3587
rect 347697 3349 347731 3383
rect 271981 3145 272015 3179
rect 151553 561 151587 595
rect 177773 2805 177807 2839
rect 177773 561 177807 595
rect 358553 561 358587 595
rect 359749 9605 359783 9639
rect 359749 561 359783 595
rect 406117 9605 406151 9639
rect 406117 561 406151 595
rect 407313 9605 407347 9639
rect 407313 561 407347 595
rect 414489 9605 414523 9639
rect 428933 9605 428967 9639
rect 428933 4777 428967 4811
rect 431141 9605 431175 9639
rect 414489 561 414523 595
rect 431141 561 431175 595
rect 432337 9605 432371 9639
rect 568773 3553 568807 3587
rect 568773 3349 568807 3383
rect 432337 561 432371 595
<< metal1 >>
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 365622 699700 365628 699712
rect 365036 699672 365628 699700
rect 365036 699660 365042 699672
rect 365622 699660 365628 699672
rect 365680 699660 365686 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 504358 696940 504364 696992
rect 504416 696980 504422 696992
rect 580166 696980 580172 696992
rect 504416 696952 580172 696980
rect 504416 696940 504422 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 348694 695484 348700 695496
rect 348655 695456 348700 695484
rect 348694 695444 348700 695456
rect 348752 695444 348758 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 542538 692724 542544 692776
rect 542596 692764 542602 692776
rect 542722 692764 542728 692776
rect 542596 692736 542728 692764
rect 542596 692724 542602 692736
rect 542722 692724 542728 692736
rect 542780 692724 542786 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 348697 685899 348755 685905
rect 348697 685865 348709 685899
rect 348743 685896 348755 685899
rect 348786 685896 348792 685908
rect 348743 685868 348792 685896
rect 348743 685865 348755 685868
rect 348697 685859 348755 685865
rect 348786 685856 348792 685868
rect 348844 685856 348850 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 429194 684428 429200 684480
rect 429252 684468 429258 684480
rect 429838 684468 429844 684480
rect 429252 684440 429844 684468
rect 429252 684428 429258 684440
rect 429838 684428 429844 684440
rect 429896 684428 429902 684480
rect 558914 684428 558920 684480
rect 558972 684468 558978 684480
rect 559650 684468 559656 684480
rect 558972 684440 559656 684468
rect 558972 684428 558978 684440
rect 559650 684428 559656 684440
rect 559708 684428 559714 684480
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 429194 683068 429200 683120
rect 429252 683108 429258 683120
rect 429565 683111 429623 683117
rect 429565 683108 429577 683111
rect 429252 683080 429577 683108
rect 429252 683068 429258 683080
rect 429565 683077 429577 683080
rect 429611 683077 429623 683111
rect 429565 683071 429623 683077
rect 542354 683068 542360 683120
rect 542412 683108 542418 683120
rect 542725 683111 542783 683117
rect 542725 683108 542737 683111
rect 542412 683080 542737 683108
rect 542412 683068 542418 683080
rect 542725 683077 542737 683080
rect 542771 683077 542783 683111
rect 542725 683071 542783 683077
rect 558914 683068 558920 683120
rect 558972 683108 558978 683120
rect 559285 683111 559343 683117
rect 559285 683108 559297 683111
rect 558972 683080 559297 683108
rect 558972 683068 558978 683080
rect 559285 683077 559297 683080
rect 559331 683077 559343 683111
rect 559285 683071 559343 683077
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 8938 681748 8944 681760
rect 3568 681720 8944 681748
rect 3568 681708 3574 681720
rect 8938 681708 8944 681720
rect 8996 681708 9002 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 348694 676172 348700 676184
rect 348655 676144 348700 676172
rect 348694 676132 348700 676144
rect 348752 676132 348758 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 494054 673480 494060 673532
rect 494112 673520 494118 673532
rect 494238 673520 494244 673532
rect 494112 673492 494244 673520
rect 494112 673480 494118 673492
rect 494238 673480 494244 673492
rect 494296 673480 494302 673532
rect 514018 673480 514024 673532
rect 514076 673520 514082 673532
rect 580166 673520 580172 673532
rect 514076 673492 580172 673520
rect 514076 673480 514082 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 348697 666587 348755 666593
rect 348697 666553 348709 666587
rect 348743 666584 348755 666587
rect 348786 666584 348792 666596
rect 348743 666556 348792 666584
rect 348743 666553 348755 666556
rect 348697 666547 348755 666553
rect 348786 666544 348792 666556
rect 348844 666544 348850 666596
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 348878 659608 348884 659660
rect 348936 659648 348942 659660
rect 349062 659648 349068 659660
rect 348936 659620 349068 659648
rect 348936 659608 348942 659620
rect 349062 659608 349068 659620
rect 349120 659608 349126 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 348973 656863 349031 656869
rect 348973 656829 348985 656863
rect 349019 656860 349031 656863
rect 349062 656860 349068 656872
rect 349019 656832 349068 656860
rect 349019 656829 349031 656832
rect 348973 656823 349031 656829
rect 349062 656820 349068 656832
rect 349120 656820 349126 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 284018 654100 284024 654152
rect 284076 654140 284082 654152
rect 284202 654140 284208 654152
rect 284076 654112 284208 654140
rect 284076 654100 284082 654112
rect 284202 654100 284208 654112
rect 284260 654100 284266 654152
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 14458 652780 14464 652792
rect 3108 652752 14464 652780
rect 3108 652740 3114 652752
rect 14458 652740 14464 652752
rect 14516 652740 14522 652792
rect 525058 650020 525064 650072
rect 525116 650060 525122 650072
rect 580166 650060 580172 650072
rect 525116 650032 580172 650060
rect 525116 650020 525122 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 348970 647272 348976 647284
rect 348931 647244 348976 647272
rect 348970 647232 348976 647244
rect 349028 647232 349034 647284
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 348970 640404 348976 640416
rect 348804 640376 348976 640404
rect 348804 640280 348832 640376
rect 348970 640364 348976 640376
rect 349028 640364 349034 640416
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 348786 640228 348792 640280
rect 348844 640228 348850 640280
rect 72786 637548 72792 637560
rect 72747 637520 72792 637548
rect 72786 637508 72792 637520
rect 72844 637508 72850 637560
rect 219066 637548 219072 637560
rect 219027 637520 219072 637548
rect 219066 637508 219072 637520
rect 219124 637508 219130 637560
rect 348786 637548 348792 637560
rect 348747 637520 348792 637548
rect 348786 637508 348792 637520
rect 348844 637508 348850 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 284018 634788 284024 634840
rect 284076 634828 284082 634840
rect 284202 634828 284208 634840
rect 284076 634800 284208 634828
rect 284076 634788 284082 634800
rect 284202 634788 284208 634800
rect 284260 634788 284266 634840
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 72789 627963 72847 627969
rect 72789 627929 72801 627963
rect 72835 627960 72847 627963
rect 73062 627960 73068 627972
rect 72835 627932 73068 627960
rect 72835 627929 72847 627932
rect 72789 627923 72847 627929
rect 73062 627920 73068 627932
rect 73120 627920 73126 627972
rect 219069 627963 219127 627969
rect 219069 627929 219081 627963
rect 219115 627960 219127 627963
rect 219342 627960 219348 627972
rect 219115 627932 219348 627960
rect 219115 627929 219127 627932
rect 219069 627923 219127 627929
rect 219342 627920 219348 627932
rect 219400 627920 219406 627972
rect 348789 627963 348847 627969
rect 348789 627929 348801 627963
rect 348835 627960 348847 627963
rect 349062 627960 349068 627972
rect 348835 627932 349068 627960
rect 348835 627929 348847 627932
rect 348789 627923 348847 627929
rect 349062 627920 349068 627932
rect 349120 627920 349126 627972
rect 519538 626560 519544 626612
rect 519596 626600 519602 626612
rect 580166 626600 580172 626612
rect 519596 626572 580172 626600
rect 519596 626560 519602 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 10318 623812 10324 623824
rect 3292 623784 10324 623812
rect 3292 623772 3298 623784
rect 10318 623772 10324 623784
rect 10376 623772 10382 623824
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 284018 615476 284024 615528
rect 284076 615516 284082 615528
rect 284202 615516 284208 615528
rect 284076 615488 284208 615516
rect 284076 615476 284082 615488
rect 284202 615476 284208 615488
rect 284260 615476 284266 615528
rect 477494 615476 477500 615528
rect 477552 615516 477558 615528
rect 477678 615516 477684 615528
rect 477552 615488 477684 615516
rect 477552 615476 477558 615488
rect 477678 615476 477684 615488
rect 477736 615476 477742 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 137738 604120 137744 604172
rect 137796 604160 137802 604172
rect 224126 604160 224132 604172
rect 137796 604132 224132 604160
rect 137796 604120 137802 604132
rect 224126 604120 224132 604132
rect 224184 604120 224190 604172
rect 106182 604052 106188 604104
rect 106240 604092 106246 604104
rect 210602 604092 210608 604104
rect 106240 604064 210608 604092
rect 106240 604052 106246 604064
rect 210602 604052 210608 604064
rect 210660 604052 210666 604104
rect 89622 603984 89628 604036
rect 89680 604024 89686 604036
rect 197078 604024 197084 604036
rect 89680 603996 197084 604024
rect 89680 603984 89686 603996
rect 197078 603984 197084 603996
rect 197136 603984 197142 604036
rect 235902 603984 235908 604036
rect 235960 604024 235966 604036
rect 291838 604024 291844 604036
rect 235960 603996 291844 604024
rect 235960 603984 235966 603996
rect 291838 603984 291844 603996
rect 291896 603984 291902 604036
rect 73062 603916 73068 603968
rect 73120 603956 73126 603968
rect 183462 603956 183468 603968
rect 73120 603928 183468 603956
rect 73120 603916 73126 603928
rect 183462 603916 183468 603928
rect 183520 603916 183526 603968
rect 219342 603916 219348 603968
rect 219400 603956 219406 603968
rect 278314 603956 278320 603968
rect 219400 603928 278320 603956
rect 219400 603916 219406 603928
rect 278314 603916 278320 603928
rect 278372 603916 278378 603968
rect 41322 603848 41328 603900
rect 41380 603888 41386 603900
rect 169938 603888 169944 603900
rect 41380 603860 169944 603888
rect 41380 603848 41386 603860
rect 169938 603848 169944 603860
rect 169996 603848 170002 603900
rect 202782 603848 202788 603900
rect 202840 603888 202846 603900
rect 264790 603888 264796 603900
rect 202840 603860 264796 603888
rect 202840 603848 202846 603860
rect 264790 603848 264796 603860
rect 264848 603848 264854 603900
rect 300762 603848 300768 603900
rect 300820 603888 300826 603900
rect 332502 603888 332508 603900
rect 300820 603860 332508 603888
rect 300820 603848 300826 603860
rect 332502 603848 332508 603860
rect 332560 603848 332566 603900
rect 427354 603848 427360 603900
rect 427412 603888 427418 603900
rect 462314 603888 462320 603900
rect 427412 603860 462320 603888
rect 427412 603848 427418 603860
rect 462314 603848 462320 603860
rect 462372 603848 462378 603900
rect 468018 603848 468024 603900
rect 468076 603888 468082 603900
rect 527174 603888 527180 603900
rect 468076 603860 527180 603888
rect 468076 603848 468082 603860
rect 527174 603848 527180 603860
rect 527232 603848 527238 603900
rect 24762 603780 24768 603832
rect 24820 603820 24826 603832
rect 156414 603820 156420 603832
rect 24820 603792 156420 603820
rect 24820 603780 24826 603792
rect 156414 603780 156420 603792
rect 156472 603780 156478 603832
rect 171042 603780 171048 603832
rect 171100 603820 171106 603832
rect 251266 603820 251272 603832
rect 171100 603792 251272 603820
rect 171100 603780 171106 603792
rect 251266 603780 251272 603792
rect 251324 603780 251330 603832
rect 284018 603780 284024 603832
rect 284076 603820 284082 603832
rect 318978 603820 318984 603832
rect 284076 603792 318984 603820
rect 284076 603780 284082 603792
rect 318978 603780 318984 603792
rect 319036 603780 319042 603832
rect 440878 603780 440884 603832
rect 440936 603820 440942 603832
rect 477678 603820 477684 603832
rect 440936 603792 477684 603820
rect 440936 603780 440942 603792
rect 477678 603780 477684 603792
rect 477736 603780 477742 603832
rect 481542 603780 481548 603832
rect 481600 603820 481606 603832
rect 542446 603820 542452 603832
rect 481600 603792 542452 603820
rect 481600 603780 481606 603792
rect 542446 603780 542452 603792
rect 542504 603780 542510 603832
rect 8018 603712 8024 603764
rect 8076 603752 8082 603764
rect 142890 603752 142896 603764
rect 8076 603724 142896 603752
rect 8076 603712 8082 603724
rect 142890 603712 142896 603724
rect 142948 603712 142954 603764
rect 154298 603712 154304 603764
rect 154356 603752 154362 603764
rect 237650 603752 237656 603764
rect 154356 603724 237656 603752
rect 154356 603712 154362 603724
rect 237650 603712 237656 603724
rect 237708 603712 237714 603764
rect 267642 603712 267648 603764
rect 267700 603752 267706 603764
rect 305454 603752 305460 603764
rect 267700 603724 305460 603752
rect 267700 603712 267706 603724
rect 305454 603712 305460 603724
rect 305512 603712 305518 603764
rect 332318 603712 332324 603764
rect 332376 603752 332382 603764
rect 346026 603752 346032 603764
rect 332376 603724 346032 603752
rect 332376 603712 332382 603724
rect 346026 603712 346032 603724
rect 346084 603712 346090 603764
rect 349062 603712 349068 603764
rect 349120 603752 349126 603764
rect 359642 603752 359648 603764
rect 349120 603724 359648 603752
rect 349120 603712 349126 603724
rect 359642 603712 359648 603724
rect 359700 603712 359706 603764
rect 386690 603712 386696 603764
rect 386748 603752 386754 603764
rect 397454 603752 397460 603764
rect 386748 603724 397460 603752
rect 386748 603712 386754 603724
rect 397454 603712 397460 603724
rect 397512 603712 397518 603764
rect 400214 603712 400220 603764
rect 400272 603752 400278 603764
rect 412726 603752 412732 603764
rect 400272 603724 412732 603752
rect 400272 603712 400278 603724
rect 412726 603712 412732 603724
rect 412784 603712 412790 603764
rect 413830 603712 413836 603764
rect 413888 603752 413894 603764
rect 429286 603752 429292 603764
rect 413888 603724 429292 603752
rect 413888 603712 413894 603724
rect 429286 603712 429292 603724
rect 429344 603712 429350 603764
rect 454402 603712 454408 603764
rect 454460 603752 454466 603764
rect 494238 603752 494244 603764
rect 454460 603724 494244 603752
rect 454460 603712 454466 603724
rect 494238 603712 494244 603724
rect 494296 603712 494302 603764
rect 495066 603712 495072 603764
rect 495124 603752 495130 603764
rect 559006 603752 559012 603764
rect 495124 603724 559012 603752
rect 495124 603712 495130 603724
rect 559006 603712 559012 603724
rect 559064 603712 559070 603764
rect 365622 603236 365628 603288
rect 365680 603276 365686 603288
rect 373166 603276 373172 603288
rect 365680 603248 373172 603276
rect 365680 603236 365686 603248
rect 373166 603236 373172 603248
rect 373224 603236 373230 603288
rect 560938 603100 560944 603152
rect 560996 603140 561002 603152
rect 580166 603140 580172 603152
rect 560996 603112 580172 603140
rect 560996 603100 561002 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 8938 596096 8944 596148
rect 8996 596136 9002 596148
rect 78674 596136 78680 596148
rect 8996 596108 78680 596136
rect 8996 596096 9002 596108
rect 78674 596096 78680 596108
rect 78732 596096 78738 596148
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 9030 594844 9036 594856
rect 3384 594816 9036 594844
rect 3384 594804 3390 594816
rect 9030 594804 9036 594816
rect 9088 594804 9094 594856
rect 520918 592016 520924 592068
rect 520976 592056 520982 592068
rect 579890 592056 579896 592068
rect 520976 592028 579896 592056
rect 520976 592016 520982 592028
rect 579890 592016 579896 592028
rect 579948 592016 579954 592068
rect 3418 585080 3424 585132
rect 3476 585120 3482 585132
rect 78674 585120 78680 585132
rect 3476 585092 78680 585120
rect 3476 585080 3482 585092
rect 78674 585080 78680 585092
rect 78732 585080 78738 585132
rect 504358 581612 504364 581664
rect 504416 581652 504422 581664
rect 514018 581652 514024 581664
rect 504416 581624 514024 581652
rect 504416 581612 504422 581624
rect 514018 581612 514024 581624
rect 514076 581612 514082 581664
rect 514018 579640 514024 579692
rect 514076 579680 514082 579692
rect 580166 579680 580172 579692
rect 514076 579652 580172 579680
rect 514076 579640 514082 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 505002 575424 505008 575476
rect 505060 575464 505066 575476
rect 580258 575464 580264 575476
rect 505060 575436 580264 575464
rect 505060 575424 505066 575436
rect 580258 575424 580264 575436
rect 580316 575424 580322 575476
rect 14458 573996 14464 574048
rect 14516 574036 14522 574048
rect 78674 574036 78680 574048
rect 14516 574008 78680 574036
rect 14516 573996 14522 574008
rect 78674 573996 78680 574008
rect 78732 573996 78738 574048
rect 9030 567808 9036 567860
rect 9088 567848 9094 567860
rect 79318 567848 79324 567860
rect 9088 567820 79324 567848
rect 9088 567808 9094 567820
rect 79318 567808 79324 567820
rect 79376 567808 79382 567860
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 8938 567236 8944 567248
rect 3476 567208 8944 567236
rect 3476 567196 3482 567208
rect 8938 567196 8944 567208
rect 8996 567196 9002 567248
rect 10318 561620 10324 561672
rect 10376 561660 10382 561672
rect 78674 561660 78680 561672
rect 10376 561632 78680 561660
rect 10376 561620 10382 561632
rect 78674 561620 78680 561632
rect 78732 561620 78738 561672
rect 509878 556180 509884 556232
rect 509936 556220 509942 556232
rect 580166 556220 580172 556232
rect 509936 556192 580172 556220
rect 509936 556180 509942 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 503806 553324 503812 553376
rect 503864 553364 503870 553376
rect 525058 553364 525064 553376
rect 503864 553336 525064 553364
rect 503864 553324 503870 553336
rect 525058 553324 525064 553336
rect 525116 553324 525122 553376
rect 3510 550536 3516 550588
rect 3568 550576 3574 550588
rect 78674 550576 78680 550588
rect 3568 550548 78680 550576
rect 3568 550536 3574 550548
rect 78674 550536 78680 550548
rect 78732 550536 78738 550588
rect 505738 545096 505744 545148
rect 505796 545136 505802 545148
rect 580166 545136 580172 545148
rect 505796 545108 580172 545136
rect 505796 545096 505802 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 505002 542308 505008 542360
rect 505060 542348 505066 542360
rect 580350 542348 580356 542360
rect 505060 542320 580356 542348
rect 505060 542308 505066 542320
rect 580350 542308 580356 542320
rect 580408 542308 580414 542360
rect 504358 537480 504364 537532
rect 504416 537520 504422 537532
rect 519538 537520 519544 537532
rect 504416 537492 519544 537520
rect 504416 537480 504422 537492
rect 519538 537480 519544 537492
rect 519596 537480 519602 537532
rect 519538 532720 519544 532772
rect 519596 532760 519602 532772
rect 580166 532760 580172 532772
rect 519596 532732 580172 532760
rect 519596 532720 519602 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 8938 527076 8944 527128
rect 8996 527116 9002 527128
rect 78674 527116 78680 527128
rect 8996 527088 78680 527116
rect 8996 527076 9002 527088
rect 78674 527076 78680 527088
rect 78732 527076 78738 527128
rect 504634 521568 504640 521620
rect 504692 521608 504698 521620
rect 560938 521608 560944 521620
rect 504692 521580 560944 521608
rect 504692 521568 504698 521580
rect 560938 521568 560944 521580
rect 560996 521568 561002 521620
rect 3418 514700 3424 514752
rect 3476 514740 3482 514752
rect 78674 514740 78680 514752
rect 3476 514712 78680 514740
rect 3476 514700 3482 514712
rect 78674 514700 78680 514712
rect 78732 514700 78738 514752
rect 505002 510552 505008 510604
rect 505060 510592 505066 510604
rect 520918 510592 520924 510604
rect 505060 510564 520924 510592
rect 505060 510552 505066 510564
rect 520918 510552 520924 510564
rect 520976 510552 520982 510604
rect 578234 509600 578240 509652
rect 578292 509640 578298 509652
rect 579982 509640 579988 509652
rect 578292 509612 579988 509640
rect 578292 509600 578298 509612
rect 579982 509600 579988 509612
rect 580040 509600 580046 509652
rect 504358 508512 504364 508564
rect 504416 508552 504422 508564
rect 578234 508552 578240 508564
rect 504416 508524 578240 508552
rect 504416 508512 504422 508524
rect 578234 508512 578240 508524
rect 578292 508512 578298 508564
rect 3510 503616 3516 503668
rect 3568 503656 3574 503668
rect 78674 503656 78680 503668
rect 3568 503628 78680 503656
rect 3568 503616 3574 503628
rect 78674 503616 78680 503628
rect 78732 503616 78738 503668
rect 505002 499468 505008 499520
rect 505060 499508 505066 499520
rect 514018 499508 514024 499520
rect 505060 499480 514024 499508
rect 505060 499468 505066 499480
rect 514018 499468 514024 499480
rect 514076 499468 514082 499520
rect 3418 492600 3424 492652
rect 3476 492640 3482 492652
rect 78674 492640 78680 492652
rect 3476 492612 78680 492640
rect 3476 492600 3482 492612
rect 78674 492600 78680 492612
rect 78732 492600 78738 492652
rect 505002 487432 505008 487484
rect 505060 487472 505066 487484
rect 509878 487472 509884 487484
rect 505060 487444 509884 487472
rect 505060 487432 505066 487444
rect 509878 487432 509884 487444
rect 509936 487432 509942 487484
rect 514018 485800 514024 485852
rect 514076 485840 514082 485852
rect 579890 485840 579896 485852
rect 514076 485812 579896 485840
rect 514076 485800 514082 485812
rect 579890 485800 579896 485812
rect 579948 485800 579954 485852
rect 3510 480156 3516 480208
rect 3568 480196 3574 480208
rect 78674 480196 78680 480208
rect 3568 480168 78680 480196
rect 3568 480156 3574 480168
rect 78674 480156 78680 480168
rect 78732 480156 78738 480208
rect 503714 477232 503720 477284
rect 503772 477272 503778 477284
rect 505738 477272 505744 477284
rect 503772 477244 505744 477272
rect 503772 477232 503778 477244
rect 505738 477232 505744 477244
rect 505796 477232 505802 477284
rect 3418 469140 3424 469192
rect 3476 469180 3482 469192
rect 78674 469180 78680 469192
rect 3476 469152 78680 469180
rect 3476 469140 3482 469152
rect 78674 469140 78680 469152
rect 78732 469140 78738 469192
rect 505002 466352 505008 466404
rect 505060 466392 505066 466404
rect 519538 466392 519544 466404
rect 505060 466364 519544 466392
rect 505060 466352 505066 466364
rect 519538 466352 519544 466364
rect 519596 466352 519602 466404
rect 505738 462340 505744 462392
rect 505796 462380 505802 462392
rect 580166 462380 580172 462392
rect 505796 462352 580172 462380
rect 505796 462340 505802 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 3418 452548 3424 452600
rect 3476 452588 3482 452600
rect 78674 452588 78680 452600
rect 3476 452560 78680 452588
rect 3476 452548 3482 452560
rect 78674 452548 78680 452560
rect 78732 452548 78738 452600
rect 505002 444320 505008 444372
rect 505060 444360 505066 444372
rect 580258 444360 580264 444372
rect 505060 444332 580264 444360
rect 505060 444320 505066 444332
rect 580258 444320 580264 444332
rect 580316 444320 580322 444372
rect 504358 438880 504364 438932
rect 504416 438920 504422 438932
rect 580166 438920 580172 438932
rect 504416 438892 580172 438920
rect 504416 438880 504422 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 79318 438852 79324 438864
rect 3200 438824 79324 438852
rect 3200 438812 3206 438824
rect 79318 438812 79324 438824
rect 79376 438812 79382 438864
rect 504634 434664 504640 434716
rect 504692 434704 504698 434716
rect 514018 434704 514024 434716
rect 504692 434676 514024 434704
rect 504692 434664 504698 434676
rect 514018 434664 514024 434676
rect 514076 434664 514082 434716
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 79318 425048 79324 425060
rect 3292 425020 79324 425048
rect 3292 425008 3298 425020
rect 79318 425008 79324 425020
rect 79376 425008 79382 425060
rect 503714 423444 503720 423496
rect 503772 423484 503778 423496
rect 505738 423484 505744 423496
rect 503772 423456 505744 423484
rect 503772 423444 503778 423456
rect 505738 423444 505744 423456
rect 505796 423444 505802 423496
rect 505002 412564 505008 412616
rect 505060 412604 505066 412616
rect 580350 412604 580356 412616
rect 505060 412576 580356 412604
rect 505060 412564 505066 412576
rect 580350 412564 580356 412576
rect 580408 412564 580414 412616
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 79410 396012 79416 396024
rect 3200 395984 79416 396012
rect 3200 395972 3206 395984
rect 79410 395972 79416 395984
rect 79468 395972 79474 396024
rect 514018 391960 514024 392012
rect 514076 392000 514082 392012
rect 579890 392000 579896 392012
rect 514076 391972 579896 392000
rect 514076 391960 514082 391972
rect 579890 391960 579896 391972
rect 579948 391960 579954 392012
rect 505002 390464 505008 390516
rect 505060 390504 505066 390516
rect 580442 390504 580448 390516
rect 505060 390476 580448 390504
rect 505060 390464 505066 390476
rect 580442 390464 580448 390476
rect 580500 390464 580506 390516
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 79502 380848 79508 380860
rect 3292 380820 79508 380848
rect 3292 380808 3298 380820
rect 79502 380808 79508 380820
rect 79560 380808 79566 380860
rect 503898 379448 503904 379500
rect 503956 379488 503962 379500
rect 580258 379488 580264 379500
rect 503956 379460 580264 379488
rect 503956 379448 503962 379460
rect 580258 379448 580264 379460
rect 580316 379448 580322 379500
rect 505002 368432 505008 368484
rect 505060 368472 505066 368484
rect 514018 368472 514024 368484
rect 505060 368444 514024 368472
rect 505060 368432 505066 368444
rect 514018 368432 514024 368444
rect 514076 368432 514082 368484
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 79318 367044 79324 367056
rect 3200 367016 79324 367044
rect 3200 367004 3206 367016
rect 79318 367004 79324 367016
rect 79376 367004 79382 367056
rect 505002 357348 505008 357400
rect 505060 357388 505066 357400
rect 580258 357388 580264 357400
rect 505060 357360 580264 357388
rect 505060 357348 505066 357360
rect 580258 357348 580264 357360
rect 580316 357348 580322 357400
rect 505002 347692 505008 347744
rect 505060 347732 505066 347744
rect 580350 347732 580356 347744
rect 505060 347704 580356 347732
rect 505060 347692 505066 347704
rect 580350 347692 580356 347704
rect 580408 347692 580414 347744
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 79410 338076 79416 338088
rect 3476 338048 79416 338076
rect 3476 338036 3482 338048
rect 79410 338036 79416 338048
rect 79468 338036 79474 338088
rect 504542 336676 504548 336728
rect 504600 336716 504606 336728
rect 580258 336716 580264 336728
rect 504600 336688 580264 336716
rect 504600 336676 504606 336688
rect 580258 336676 580264 336688
rect 580316 336676 580322 336728
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 79686 324272 79692 324284
rect 3292 324244 79692 324272
rect 3292 324232 3298 324244
rect 79686 324232 79692 324244
rect 79744 324232 79750 324284
rect 505002 322872 505008 322924
rect 505060 322912 505066 322924
rect 580166 322912 580172 322924
rect 505060 322884 580172 322912
rect 505060 322872 505066 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 8938 316004 8944 316056
rect 8996 316044 9002 316056
rect 78674 316044 78680 316056
rect 8996 316016 78680 316044
rect 8996 316004 9002 316016
rect 78674 316004 78680 316016
rect 78732 316004 78738 316056
rect 504082 311788 504088 311840
rect 504140 311828 504146 311840
rect 580166 311828 580172 311840
rect 504140 311800 580172 311828
rect 504140 311788 504146 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 79318 309108 79324 309120
rect 3384 309080 79324 309108
rect 3384 309068 3390 309080
rect 79318 309068 79324 309080
rect 79376 309068 79382 309120
rect 504542 299412 504548 299464
rect 504600 299452 504606 299464
rect 579798 299452 579804 299464
rect 504600 299424 579804 299452
rect 504600 299412 504606 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 79594 295304 79600 295316
rect 3476 295276 79600 295304
rect 3476 295264 3482 295276
rect 79594 295264 79600 295276
rect 79652 295264 79658 295316
rect 17218 281528 17224 281580
rect 17276 281568 17282 281580
rect 78674 281568 78680 281580
rect 17276 281540 78680 281568
rect 17276 281528 17282 281540
rect 78674 281528 78680 281540
rect 78732 281528 78738 281580
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 79502 280140 79508 280152
rect 3476 280112 79508 280140
rect 3476 280100 3482 280112
rect 79502 280100 79508 280112
rect 79560 280100 79566 280152
rect 504358 275952 504364 276004
rect 504416 275992 504422 276004
rect 580166 275992 580172 276004
rect 504416 275964 580172 275992
rect 504416 275952 504422 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3142 266296 3148 266348
rect 3200 266336 3206 266348
rect 79410 266336 79416 266348
rect 3200 266308 79416 266336
rect 3200 266296 3206 266308
rect 79410 266296 79416 266308
rect 79468 266296 79474 266348
rect 504450 264868 504456 264920
rect 504508 264908 504514 264920
rect 580166 264908 580172 264920
rect 504508 264880 580172 264908
rect 504508 264868 504514 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 504358 252492 504364 252544
rect 504416 252532 504422 252544
rect 579798 252532 579804 252544
rect 504416 252504 579804 252532
rect 504416 252492 504422 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3234 252424 3240 252476
rect 3292 252464 3298 252476
rect 8938 252464 8944 252476
rect 3292 252436 8944 252464
rect 3292 252424 3298 252436
rect 8938 252424 8944 252436
rect 8996 252424 9002 252476
rect 28258 247052 28264 247104
rect 28316 247092 28322 247104
rect 78674 247092 78680 247104
rect 28316 247064 78680 247092
rect 28316 247052 28322 247064
rect 78674 247052 78680 247064
rect 78732 247052 78738 247104
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 79318 237368 79324 237380
rect 3476 237340 79324 237368
rect 3476 237328 3482 237340
rect 79318 237328 79324 237340
rect 79376 237328 79382 237380
rect 504542 229032 504548 229084
rect 504600 229072 504606 229084
rect 580166 229072 580172 229084
rect 504600 229044 580172 229072
rect 504600 229032 504606 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 14458 223592 14464 223644
rect 14516 223632 14522 223644
rect 78674 223632 78680 223644
rect 14516 223604 78680 223632
rect 14516 223592 14522 223604
rect 78674 223592 78680 223604
rect 78732 223592 78738 223644
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 79594 223564 79600 223576
rect 3200 223536 79600 223564
rect 3200 223524 3206 223536
rect 79594 223524 79600 223536
rect 79652 223524 79658 223576
rect 504450 217948 504456 218000
rect 504508 217988 504514 218000
rect 580166 217988 580172 218000
rect 504508 217960 580172 217988
rect 504508 217948 504514 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 8938 211148 8944 211200
rect 8996 211188 9002 211200
rect 78674 211188 78680 211200
rect 8996 211160 78680 211188
rect 8996 211148 9002 211160
rect 78674 211148 78680 211160
rect 78732 211148 78738 211200
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 17218 208332 17224 208344
rect 3476 208304 17224 208332
rect 3476 208292 3482 208304
rect 17218 208292 17224 208304
rect 17276 208292 17282 208344
rect 504358 205572 504364 205624
rect 504416 205612 504422 205624
rect 579798 205612 579804 205624
rect 504416 205584 579804 205612
rect 504416 205572 504422 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 79502 194528 79508 194540
rect 3200 194500 79508 194528
rect 3200 194488 3206 194500
rect 79502 194488 79508 194500
rect 79560 194488 79566 194540
rect 19978 189048 19984 189100
rect 20036 189088 20042 189100
rect 78674 189088 78680 189100
rect 20036 189060 78680 189088
rect 20036 189048 20042 189060
rect 78674 189048 78680 189060
rect 78732 189048 78738 189100
rect 504634 182112 504640 182164
rect 504692 182152 504698 182164
rect 580166 182152 580172 182164
rect 504692 182124 580172 182152
rect 504692 182112 504698 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 79410 180792 79416 180804
rect 3292 180764 79416 180792
rect 3292 180752 3298 180764
rect 79410 180752 79416 180764
rect 79468 180752 79474 180804
rect 17218 176672 17224 176724
rect 17276 176712 17282 176724
rect 78674 176712 78680 176724
rect 17276 176684 78680 176712
rect 17276 176672 17282 176684
rect 78674 176672 78680 176684
rect 78732 176672 78738 176724
rect 504542 171028 504548 171080
rect 504600 171068 504606 171080
rect 580166 171068 580172 171080
rect 504600 171040 580172 171068
rect 504600 171028 504606 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 28258 165560 28264 165572
rect 3568 165532 28264 165560
rect 3568 165520 3574 165532
rect 28258 165520 28264 165532
rect 28316 165520 28322 165572
rect 504450 158652 504456 158704
rect 504508 158692 504514 158704
rect 579798 158692 579804 158704
rect 504508 158664 579804 158692
rect 504508 158652 504514 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 79318 151756 79324 151768
rect 3200 151728 79324 151756
rect 3200 151716 3206 151728
rect 79318 151716 79324 151728
rect 79376 151716 79382 151768
rect 10318 142128 10324 142180
rect 10376 142168 10382 142180
rect 78674 142168 78680 142180
rect 10376 142140 78680 142168
rect 10376 142128 10382 142140
rect 78674 142128 78680 142140
rect 78732 142128 78738 142180
rect 505002 139408 505008 139460
rect 505060 139448 505066 139460
rect 519538 139448 519544 139460
rect 505060 139420 519544 139448
rect 505060 139408 505066 139420
rect 519538 139408 519544 139420
rect 519596 139408 519602 139460
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 14458 136592 14464 136604
rect 3292 136564 14464 136592
rect 3292 136552 3298 136564
rect 14458 136552 14464 136564
rect 14516 136552 14522 136604
rect 504358 135192 504364 135244
rect 504416 135232 504422 135244
rect 580166 135232 580172 135244
rect 504416 135204 580172 135232
rect 504416 135192 504422 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 504818 124108 504824 124160
rect 504876 124148 504882 124160
rect 580166 124148 580172 124160
rect 504876 124120 580172 124148
rect 504876 124108 504882 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 8938 122788 8944 122800
rect 3476 122760 8944 122788
rect 3476 122748 3482 122760
rect 8938 122748 8944 122760
rect 8996 122748 9002 122800
rect 504726 111732 504732 111784
rect 504784 111772 504790 111784
rect 579798 111772 579804 111784
rect 504784 111744 579804 111772
rect 504784 111732 504790 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 79686 108984 79692 108996
rect 3292 108956 79692 108984
rect 3292 108944 3298 108956
rect 79686 108944 79692 108956
rect 79744 108944 79750 108996
rect 157978 100648 157984 100700
rect 158036 100688 158042 100700
rect 165982 100688 165988 100700
rect 158036 100660 165988 100688
rect 158036 100648 158042 100660
rect 165982 100648 165988 100660
rect 166040 100648 166046 100700
rect 302510 100648 302516 100700
rect 302568 100688 302574 100700
rect 303522 100688 303528 100700
rect 302568 100660 303528 100688
rect 302568 100648 302574 100660
rect 303522 100648 303528 100660
rect 303580 100648 303586 100700
rect 309410 100648 309416 100700
rect 309468 100688 309474 100700
rect 310422 100688 310428 100700
rect 309468 100660 310428 100688
rect 309468 100648 309474 100660
rect 310422 100648 310428 100660
rect 310480 100648 310486 100700
rect 311894 100648 311900 100700
rect 311952 100688 311958 100700
rect 313090 100688 313096 100700
rect 311952 100660 313096 100688
rect 311952 100648 311958 100660
rect 313090 100648 313096 100660
rect 313148 100648 313154 100700
rect 313642 100648 313648 100700
rect 313700 100688 313706 100700
rect 314562 100688 314568 100700
rect 313700 100660 314568 100688
rect 313700 100648 313706 100660
rect 314562 100648 314568 100660
rect 314620 100648 314626 100700
rect 316218 100648 316224 100700
rect 316276 100688 316282 100700
rect 317230 100688 317236 100700
rect 316276 100660 317236 100688
rect 316276 100648 316282 100660
rect 317230 100648 317236 100660
rect 317288 100648 317294 100700
rect 317874 100648 317880 100700
rect 317932 100688 317938 100700
rect 318702 100688 318708 100700
rect 317932 100660 318708 100688
rect 317932 100648 317938 100660
rect 318702 100648 318708 100660
rect 318760 100648 318766 100700
rect 323026 100648 323032 100700
rect 323084 100688 323090 100700
rect 324222 100688 324228 100700
rect 323084 100660 324228 100688
rect 323084 100648 323090 100660
rect 324222 100648 324228 100660
rect 324280 100648 324286 100700
rect 324774 100648 324780 100700
rect 324832 100688 324838 100700
rect 325510 100688 325516 100700
rect 324832 100660 325516 100688
rect 324832 100648 324838 100660
rect 325510 100648 325516 100660
rect 325568 100648 325574 100700
rect 327258 100648 327264 100700
rect 327316 100688 327322 100700
rect 328362 100688 328368 100700
rect 327316 100660 328368 100688
rect 327316 100648 327322 100660
rect 328362 100648 328368 100660
rect 328420 100648 328426 100700
rect 329006 100648 329012 100700
rect 329064 100688 329070 100700
rect 329742 100688 329748 100700
rect 329064 100660 329748 100688
rect 329064 100648 329070 100660
rect 329742 100648 329748 100660
rect 329800 100648 329806 100700
rect 329834 100648 329840 100700
rect 329892 100688 329898 100700
rect 331030 100688 331036 100700
rect 329892 100660 331036 100688
rect 329892 100648 329898 100660
rect 331030 100648 331036 100660
rect 331088 100648 331094 100700
rect 331582 100648 331588 100700
rect 331640 100688 331646 100700
rect 333238 100688 333244 100700
rect 331640 100660 333244 100688
rect 331640 100648 331646 100660
rect 333238 100648 333244 100660
rect 333296 100648 333302 100700
rect 334158 100648 334164 100700
rect 334216 100688 334222 100700
rect 335262 100688 335268 100700
rect 334216 100660 335268 100688
rect 334216 100648 334222 100660
rect 335262 100648 335268 100660
rect 335320 100648 335326 100700
rect 335814 100648 335820 100700
rect 335872 100688 335878 100700
rect 336550 100688 336556 100700
rect 335872 100660 336556 100688
rect 335872 100648 335878 100660
rect 336550 100648 336556 100660
rect 336608 100648 336614 100700
rect 338390 100648 338396 100700
rect 338448 100688 338454 100700
rect 339402 100688 339408 100700
rect 338448 100660 339408 100688
rect 338448 100648 338454 100660
rect 339402 100648 339408 100660
rect 339460 100648 339466 100700
rect 345198 100648 345204 100700
rect 345256 100688 345262 100700
rect 346210 100688 346216 100700
rect 345256 100660 346216 100688
rect 345256 100648 345262 100660
rect 346210 100648 346216 100660
rect 346268 100648 346274 100700
rect 353754 100648 353760 100700
rect 353812 100688 353818 100700
rect 354582 100688 354588 100700
rect 353812 100660 354588 100688
rect 353812 100648 353818 100660
rect 354582 100648 354588 100660
rect 354640 100648 354646 100700
rect 356330 100648 356336 100700
rect 356388 100688 356394 100700
rect 357342 100688 357348 100700
rect 356388 100660 357348 100688
rect 356388 100648 356394 100660
rect 357342 100648 357348 100660
rect 357400 100648 357406 100700
rect 374270 100648 374276 100700
rect 374328 100688 374334 100700
rect 375190 100688 375196 100700
rect 374328 100660 375196 100688
rect 374328 100648 374334 100660
rect 375190 100648 375196 100660
rect 375248 100648 375254 100700
rect 383654 100648 383660 100700
rect 383712 100688 383718 100700
rect 384942 100688 384948 100700
rect 383712 100660 384948 100688
rect 383712 100648 383718 100660
rect 384942 100648 384948 100660
rect 385000 100648 385006 100700
rect 421190 100648 421196 100700
rect 421248 100688 421254 100700
rect 422202 100688 422208 100700
rect 421248 100660 422208 100688
rect 421248 100648 421254 100660
rect 422202 100648 422208 100660
rect 422260 100648 422266 100700
rect 425422 100648 425428 100700
rect 425480 100688 425486 100700
rect 426250 100688 426256 100700
rect 425480 100660 426256 100688
rect 425480 100648 425486 100660
rect 426250 100648 426256 100660
rect 426308 100648 426314 100700
rect 426342 100648 426348 100700
rect 426400 100688 426406 100700
rect 427078 100688 427084 100700
rect 426400 100660 427084 100688
rect 426400 100648 426406 100660
rect 427078 100648 427084 100660
rect 427136 100648 427142 100700
rect 430574 100648 430580 100700
rect 430632 100688 430638 100700
rect 431862 100688 431868 100700
rect 430632 100660 431868 100688
rect 430632 100648 430638 100660
rect 431862 100648 431868 100660
rect 431920 100648 431926 100700
rect 432322 100648 432328 100700
rect 432380 100688 432386 100700
rect 433978 100688 433984 100700
rect 432380 100660 433984 100688
rect 432380 100648 432386 100660
rect 433978 100648 433984 100660
rect 434036 100648 434042 100700
rect 434898 100648 434904 100700
rect 434956 100688 434962 100700
rect 436002 100688 436008 100700
rect 434956 100660 436008 100688
rect 434956 100648 434962 100660
rect 436002 100648 436008 100660
rect 436060 100648 436066 100700
rect 439130 100648 439136 100700
rect 439188 100688 439194 100700
rect 440142 100688 440148 100700
rect 439188 100660 440148 100688
rect 439188 100648 439194 100660
rect 440142 100648 440148 100660
rect 440200 100648 440206 100700
rect 444282 100648 444288 100700
rect 444340 100688 444346 100700
rect 445018 100688 445024 100700
rect 444340 100660 445024 100688
rect 444340 100648 444346 100660
rect 445018 100648 445024 100660
rect 445076 100648 445082 100700
rect 445938 100648 445944 100700
rect 445996 100688 446002 100700
rect 446950 100688 446956 100700
rect 445996 100660 446956 100688
rect 445996 100648 446002 100660
rect 446950 100648 446956 100660
rect 447008 100648 447014 100700
rect 448514 100648 448520 100700
rect 448572 100688 448578 100700
rect 449710 100688 449716 100700
rect 448572 100660 449716 100688
rect 448572 100648 448578 100660
rect 449710 100648 449716 100660
rect 449768 100648 449774 100700
rect 452746 100648 452752 100700
rect 452804 100688 452810 100700
rect 453850 100688 453856 100700
rect 452804 100660 453856 100688
rect 452804 100648 452810 100660
rect 453850 100648 453856 100660
rect 453908 100648 453914 100700
rect 466454 100648 466460 100700
rect 466512 100688 466518 100700
rect 467742 100688 467748 100700
rect 466512 100660 467748 100688
rect 466512 100648 466518 100660
rect 467742 100648 467748 100660
rect 467800 100648 467806 100700
rect 468110 100648 468116 100700
rect 468168 100688 468174 100700
rect 469858 100688 469864 100700
rect 468168 100660 469864 100688
rect 468168 100648 468174 100660
rect 469858 100648 469864 100660
rect 469916 100648 469922 100700
rect 475010 100648 475016 100700
rect 475068 100688 475074 100700
rect 475930 100688 475936 100700
rect 475068 100660 475936 100688
rect 475068 100648 475074 100660
rect 475930 100648 475936 100660
rect 475988 100648 475994 100700
rect 305086 100580 305092 100632
rect 305144 100620 305150 100632
rect 306282 100620 306288 100632
rect 305144 100592 306288 100620
rect 305144 100580 305150 100592
rect 306282 100580 306288 100592
rect 306340 100580 306346 100632
rect 340966 100580 340972 100632
rect 341024 100620 341030 100632
rect 342162 100620 342168 100632
rect 341024 100592 342168 100620
rect 341024 100580 341030 100592
rect 342162 100580 342168 100592
rect 342220 100580 342226 100632
rect 342622 100580 342628 100632
rect 342680 100620 342686 100632
rect 347038 100620 347044 100632
rect 342680 100592 347044 100620
rect 342680 100580 342686 100592
rect 347038 100580 347044 100592
rect 347096 100580 347102 100632
rect 347774 100580 347780 100632
rect 347832 100620 347838 100632
rect 348970 100620 348976 100632
rect 347832 100592 348976 100620
rect 347832 100580 347838 100592
rect 348970 100580 348976 100592
rect 349028 100580 349034 100632
rect 352006 100580 352012 100632
rect 352064 100620 352070 100632
rect 353202 100620 353208 100632
rect 352064 100592 353208 100620
rect 352064 100580 352070 100592
rect 353202 100580 353208 100592
rect 353260 100580 353266 100632
rect 371694 100580 371700 100632
rect 371752 100620 371758 100632
rect 372522 100620 372528 100632
rect 371752 100592 372528 100620
rect 371752 100580 371758 100592
rect 372522 100580 372528 100592
rect 372580 100580 372586 100632
rect 387886 100580 387892 100632
rect 387944 100620 387950 100632
rect 389082 100620 389088 100632
rect 387944 100592 389088 100620
rect 387944 100580 387950 100592
rect 389082 100580 389088 100592
rect 389140 100580 389146 100632
rect 423766 100580 423772 100632
rect 423824 100620 423830 100632
rect 424962 100620 424968 100632
rect 423824 100592 424968 100620
rect 423824 100580 423830 100592
rect 424962 100580 424968 100592
rect 425020 100580 425026 100632
rect 470686 100580 470692 100632
rect 470744 100620 470750 100632
rect 471882 100620 471888 100632
rect 470744 100592 471888 100620
rect 470744 100580 470750 100592
rect 471882 100580 471888 100592
rect 471940 100580 471946 100632
rect 369946 100512 369952 100564
rect 370004 100552 370010 100564
rect 376018 100552 376024 100564
rect 370004 100524 376024 100552
rect 370004 100512 370010 100524
rect 376018 100512 376024 100524
rect 376076 100512 376082 100564
rect 200758 100376 200764 100428
rect 200816 100416 200822 100428
rect 201770 100416 201776 100428
rect 200816 100388 201776 100416
rect 200816 100376 200822 100388
rect 201770 100376 201776 100388
rect 201828 100376 201834 100428
rect 337562 100104 337568 100156
rect 337620 100144 337626 100156
rect 338758 100144 338764 100156
rect 337620 100116 338764 100144
rect 337620 100104 337626 100116
rect 338758 100104 338764 100116
rect 338816 100104 338822 100156
rect 447686 100104 447692 100156
rect 447744 100144 447750 100156
rect 448422 100144 448428 100156
rect 447744 100116 448428 100144
rect 447744 100104 447750 100116
rect 448422 100104 448428 100116
rect 448480 100104 448486 100156
rect 485222 100104 485228 100156
rect 485280 100144 485286 100156
rect 502978 100144 502984 100156
rect 485280 100116 502984 100144
rect 485280 100104 485286 100116
rect 502978 100104 502984 100116
rect 503036 100104 503042 100156
rect 75178 100036 75184 100088
rect 75236 100076 75242 100088
rect 87414 100076 87420 100088
rect 75236 100048 87420 100076
rect 75236 100036 75242 100048
rect 87414 100036 87420 100048
rect 87472 100036 87478 100088
rect 124858 100036 124864 100088
rect 124916 100076 124922 100088
rect 153194 100076 153200 100088
rect 124916 100048 153200 100076
rect 124916 100036 124922 100048
rect 153194 100036 153200 100048
rect 153252 100036 153258 100088
rect 167638 100036 167644 100088
rect 167696 100076 167702 100088
rect 200942 100076 200948 100088
rect 167696 100048 200948 100076
rect 167696 100036 167702 100048
rect 200942 100036 200948 100048
rect 201000 100036 201006 100088
rect 360562 100036 360568 100088
rect 360620 100076 360626 100088
rect 370498 100076 370504 100088
rect 360620 100048 370504 100076
rect 360620 100036 360626 100048
rect 370498 100036 370504 100048
rect 370556 100036 370562 100088
rect 472434 100036 472440 100088
rect 472492 100076 472498 100088
rect 507118 100076 507124 100088
rect 472492 100048 507124 100076
rect 472492 100036 472498 100048
rect 507118 100036 507124 100048
rect 507176 100036 507182 100088
rect 8938 99968 8944 100020
rect 8996 100008 9002 100020
rect 83182 100008 83188 100020
rect 8996 99980 83188 100008
rect 8996 99968 9002 99980
rect 83182 99968 83188 99980
rect 83240 99968 83246 100020
rect 88242 99968 88248 100020
rect 88300 100008 88306 100020
rect 118970 100008 118976 100020
rect 88300 99980 118976 100008
rect 88300 99968 88306 99980
rect 118970 99968 118976 99980
rect 119028 99968 119034 100020
rect 120718 99968 120724 100020
rect 120776 100008 120782 100020
rect 129274 100008 129280 100020
rect 120776 99980 129280 100008
rect 120776 99968 120782 99980
rect 129274 99968 129280 99980
rect 129332 99968 129338 100020
rect 131758 99968 131764 100020
rect 131816 100008 131822 100020
rect 136910 100008 136916 100020
rect 131816 99980 136916 100008
rect 131816 99968 131822 99980
rect 136910 99968 136916 99980
rect 136968 99968 136974 100020
rect 142798 99968 142804 100020
rect 142856 100008 142862 100020
rect 177022 100008 177028 100020
rect 142856 99980 177028 100008
rect 142856 99968 142862 99980
rect 177022 99968 177028 99980
rect 177080 99968 177086 100020
rect 178678 99968 178684 100020
rect 178736 100008 178742 100020
rect 183922 100008 183928 100020
rect 178736 99980 183928 100008
rect 178736 99968 178742 99980
rect 183922 99968 183928 99980
rect 183980 99968 183986 100020
rect 207658 99968 207664 100020
rect 207716 100008 207722 100020
rect 224034 100008 224040 100020
rect 207716 99980 224040 100008
rect 207716 99968 207722 99980
rect 224034 99968 224040 99980
rect 224092 99968 224098 100020
rect 326430 99968 326436 100020
rect 326488 100008 326494 100020
rect 337378 100008 337384 100020
rect 326488 99980 337384 100008
rect 326488 99968 326494 99980
rect 337378 99968 337384 99980
rect 337436 99968 337442 100020
rect 346946 99968 346952 100020
rect 347004 100008 347010 100020
rect 368566 100008 368572 100020
rect 347004 99980 368572 100008
rect 347004 99968 347010 99980
rect 368566 99968 368572 99980
rect 368624 99968 368630 100020
rect 375926 99968 375932 100020
rect 375984 100008 375990 100020
rect 377398 100008 377404 100020
rect 375984 99980 377404 100008
rect 375984 99968 375990 99980
rect 377398 99968 377404 99980
rect 377456 99968 377462 100020
rect 377674 99968 377680 100020
rect 377732 100008 377738 100020
rect 411346 100008 411352 100020
rect 377732 99980 411352 100008
rect 377732 99968 377738 99980
rect 411346 99968 411352 99980
rect 411404 99968 411410 100020
rect 431402 99968 431408 100020
rect 431460 100008 431466 100020
rect 483658 100008 483664 100020
rect 431460 99980 483664 100008
rect 431460 99968 431466 99980
rect 483658 99968 483664 99980
rect 483716 99968 483722 100020
rect 498010 99968 498016 100020
rect 498068 100008 498074 100020
rect 545758 100008 545764 100020
rect 498068 99980 545764 100008
rect 498068 99968 498074 99980
rect 545758 99968 545764 99980
rect 545816 99968 545822 100020
rect 358906 99832 358912 99884
rect 358964 99872 358970 99884
rect 360102 99872 360108 99884
rect 358964 99844 360108 99872
rect 358964 99832 358970 99844
rect 360102 99832 360108 99844
rect 360160 99832 360166 99884
rect 381078 99832 381084 99884
rect 381136 99872 381142 99884
rect 382182 99872 382188 99884
rect 381136 99844 382188 99872
rect 381136 99832 381142 99844
rect 382182 99832 382188 99844
rect 382240 99832 382246 99884
rect 418614 99764 418620 99816
rect 418672 99804 418678 99816
rect 420178 99804 420184 99816
rect 418672 99776 420184 99804
rect 418672 99764 418678 99776
rect 420178 99764 420184 99776
rect 420236 99764 420242 99816
rect 450262 99764 450268 99816
rect 450320 99804 450326 99816
rect 451918 99804 451924 99816
rect 450320 99776 451924 99804
rect 450320 99764 450326 99776
rect 451918 99764 451924 99776
rect 451976 99764 451982 99816
rect 376846 99628 376852 99680
rect 376904 99668 376910 99680
rect 378042 99668 378048 99680
rect 376904 99640 378048 99668
rect 376904 99628 376910 99640
rect 378042 99628 378048 99640
rect 378100 99628 378106 99680
rect 339218 99492 339224 99544
rect 339276 99532 339282 99544
rect 344278 99532 344284 99544
rect 339276 99504 344284 99532
rect 339276 99492 339282 99504
rect 344278 99492 344284 99504
rect 344336 99492 344342 99544
rect 318794 99424 318800 99476
rect 318852 99464 318858 99476
rect 326338 99464 326344 99476
rect 318852 99436 326344 99464
rect 318852 99424 318858 99436
rect 326338 99424 326344 99436
rect 326396 99424 326402 99476
rect 397270 99424 397276 99476
rect 397328 99464 397334 99476
rect 399478 99464 399484 99476
rect 397328 99436 399484 99464
rect 397328 99424 397334 99436
rect 399478 99424 399484 99436
rect 399536 99424 399542 99476
rect 413554 99424 413560 99476
rect 413612 99464 413618 99476
rect 416038 99464 416044 99476
rect 413612 99436 416044 99464
rect 413612 99424 413618 99436
rect 416038 99424 416044 99436
rect 416096 99424 416102 99476
rect 427170 99424 427176 99476
rect 427228 99464 427234 99476
rect 431218 99464 431224 99476
rect 427228 99436 431224 99464
rect 427228 99424 427234 99436
rect 431218 99424 431224 99436
rect 431276 99424 431282 99476
rect 443362 99424 443368 99476
rect 443420 99464 443426 99476
rect 447778 99464 447784 99476
rect 443420 99436 447784 99464
rect 443420 99424 443426 99436
rect 447778 99424 447784 99436
rect 447836 99424 447842 99476
rect 77938 99356 77944 99408
rect 77996 99396 78002 99408
rect 84010 99396 84016 99408
rect 77996 99368 84016 99396
rect 77996 99356 78002 99368
rect 84010 99356 84016 99368
rect 84068 99356 84074 99408
rect 91738 99356 91744 99408
rect 91796 99396 91802 99408
rect 94222 99396 94228 99408
rect 91796 99368 94228 99396
rect 91796 99356 91802 99368
rect 94222 99356 94228 99368
rect 94280 99356 94286 99408
rect 106918 99356 106924 99408
rect 106976 99396 106982 99408
rect 112162 99396 112168 99408
rect 106976 99368 112168 99396
rect 106976 99356 106982 99368
rect 112162 99356 112168 99368
rect 112220 99356 112226 99408
rect 128998 99356 129004 99408
rect 129056 99396 129062 99408
rect 130102 99396 130108 99408
rect 129056 99368 130108 99396
rect 129056 99356 129062 99368
rect 130102 99356 130108 99368
rect 130160 99356 130166 99408
rect 156598 99356 156604 99408
rect 156656 99396 156662 99408
rect 157426 99396 157432 99408
rect 156656 99368 157432 99396
rect 156656 99356 156662 99368
rect 157426 99356 157432 99368
rect 157484 99356 157490 99408
rect 160094 99356 160100 99408
rect 160152 99396 160158 99408
rect 160830 99396 160836 99408
rect 160152 99368 160836 99396
rect 160152 99356 160158 99368
rect 160830 99356 160836 99368
rect 160888 99356 160894 99408
rect 185578 99356 185584 99408
rect 185636 99396 185642 99408
rect 188154 99396 188160 99408
rect 185636 99368 188160 99396
rect 185636 99356 185642 99368
rect 188154 99356 188160 99368
rect 188212 99356 188218 99408
rect 203518 99356 203524 99408
rect 203576 99396 203582 99408
rect 206094 99396 206100 99408
rect 203576 99368 206100 99396
rect 203576 99356 203582 99368
rect 206094 99356 206100 99368
rect 206152 99356 206158 99408
rect 214558 99356 214564 99408
rect 214616 99396 214622 99408
rect 219710 99396 219716 99408
rect 214616 99368 219716 99396
rect 214616 99356 214622 99368
rect 219710 99356 219716 99368
rect 219768 99356 219774 99408
rect 239398 99356 239404 99408
rect 239456 99396 239462 99408
rect 241974 99396 241980 99408
rect 239456 99368 241980 99396
rect 239456 99356 239462 99368
rect 241974 99356 241980 99368
rect 242032 99356 242038 99408
rect 293126 99356 293132 99408
rect 293184 99396 293190 99408
rect 293862 99396 293868 99408
rect 293184 99368 293868 99396
rect 293184 99356 293190 99368
rect 293862 99356 293868 99368
rect 293920 99356 293926 99408
rect 294046 99356 294052 99408
rect 294104 99396 294110 99408
rect 295150 99396 295156 99408
rect 294104 99368 295156 99396
rect 294104 99356 294110 99368
rect 295150 99356 295156 99368
rect 295208 99356 295214 99408
rect 295702 99356 295708 99408
rect 295760 99396 295766 99408
rect 296622 99396 296628 99408
rect 295760 99368 296628 99396
rect 295760 99356 295766 99368
rect 296622 99356 296628 99368
rect 296680 99356 296686 99408
rect 298278 99356 298284 99408
rect 298336 99396 298342 99408
rect 299382 99396 299388 99408
rect 298336 99368 299388 99396
rect 298336 99356 298342 99368
rect 299382 99356 299388 99368
rect 299440 99356 299446 99408
rect 300854 99356 300860 99408
rect 300912 99396 300918 99408
rect 302142 99396 302148 99408
rect 300912 99368 302148 99396
rect 300912 99356 300918 99368
rect 302142 99356 302148 99368
rect 302200 99356 302206 99408
rect 363138 99356 363144 99408
rect 363196 99396 363202 99408
rect 364150 99396 364156 99408
rect 363196 99368 364156 99396
rect 363196 99356 363202 99368
rect 364150 99356 364156 99368
rect 364208 99356 364214 99408
rect 364886 99356 364892 99408
rect 364944 99396 364950 99408
rect 365622 99396 365628 99408
rect 364944 99368 365628 99396
rect 364944 99356 364950 99368
rect 365622 99356 365628 99368
rect 365680 99356 365686 99408
rect 365714 99356 365720 99408
rect 365772 99396 365778 99408
rect 367002 99396 367008 99408
rect 365772 99368 367008 99396
rect 365772 99356 365778 99368
rect 367002 99356 367008 99368
rect 367060 99356 367066 99408
rect 389634 99356 389640 99408
rect 389692 99396 389698 99408
rect 389692 99368 390416 99396
rect 389692 99356 389698 99368
rect 386138 99288 386144 99340
rect 386196 99328 386202 99340
rect 386322 99328 386328 99340
rect 386196 99300 386328 99328
rect 386196 99288 386202 99300
rect 386322 99288 386328 99300
rect 386380 99288 386386 99340
rect 390388 99260 390416 99368
rect 390462 99356 390468 99408
rect 390520 99396 390526 99408
rect 391198 99396 391204 99408
rect 390520 99368 391204 99396
rect 390520 99356 390526 99368
rect 391198 99356 391204 99368
rect 391256 99356 391262 99408
rect 392210 99356 392216 99408
rect 392268 99396 392274 99408
rect 393130 99396 393136 99408
rect 392268 99368 393136 99396
rect 392268 99356 392274 99368
rect 393130 99356 393136 99368
rect 393188 99356 393194 99408
rect 394694 99356 394700 99408
rect 394752 99396 394758 99408
rect 395890 99396 395896 99408
rect 394752 99368 395896 99396
rect 394752 99356 394758 99368
rect 395890 99356 395896 99368
rect 395948 99356 395954 99408
rect 396442 99356 396448 99408
rect 396500 99396 396506 99408
rect 397362 99396 397368 99408
rect 396500 99368 397368 99396
rect 396500 99356 396506 99368
rect 397362 99356 397368 99368
rect 397420 99356 397426 99408
rect 399018 99356 399024 99408
rect 399076 99396 399082 99408
rect 400030 99396 400036 99408
rect 399076 99368 400036 99396
rect 399076 99356 399082 99368
rect 400030 99356 400036 99368
rect 400088 99356 400094 99408
rect 400674 99356 400680 99408
rect 400732 99396 400738 99408
rect 401502 99396 401508 99408
rect 400732 99368 401508 99396
rect 400732 99356 400738 99368
rect 401502 99356 401508 99368
rect 401560 99356 401566 99408
rect 401594 99356 401600 99408
rect 401652 99396 401658 99408
rect 402790 99396 402796 99408
rect 401652 99368 402796 99396
rect 401652 99356 401658 99368
rect 402790 99356 402796 99368
rect 402848 99356 402854 99408
rect 403250 99356 403256 99408
rect 403308 99396 403314 99408
rect 404170 99396 404176 99408
rect 403308 99368 404176 99396
rect 403308 99356 403314 99368
rect 404170 99356 404176 99368
rect 404228 99356 404234 99408
rect 405826 99356 405832 99408
rect 405884 99396 405890 99408
rect 407022 99396 407028 99408
rect 405884 99368 407028 99396
rect 405884 99356 405890 99368
rect 407022 99356 407028 99368
rect 407080 99356 407086 99408
rect 408402 99356 408408 99408
rect 408460 99396 408466 99408
rect 409138 99396 409144 99408
rect 408460 99368 409144 99396
rect 408460 99356 408466 99368
rect 409138 99356 409144 99368
rect 409196 99356 409202 99408
rect 410058 99356 410064 99408
rect 410116 99396 410122 99408
rect 411162 99396 411168 99408
rect 410116 99368 411168 99396
rect 410116 99356 410122 99368
rect 411162 99356 411168 99368
rect 411220 99356 411226 99408
rect 411806 99356 411812 99408
rect 411864 99396 411870 99408
rect 412542 99396 412548 99408
rect 411864 99368 412548 99396
rect 411864 99356 411870 99368
rect 412542 99356 412548 99368
rect 412600 99356 412606 99408
rect 412634 99356 412640 99408
rect 412692 99396 412698 99408
rect 413922 99396 413928 99408
rect 412692 99368 413928 99396
rect 412692 99356 412698 99368
rect 413922 99356 413928 99368
rect 413980 99356 413986 99408
rect 416958 99356 416964 99408
rect 417016 99396 417022 99408
rect 417970 99396 417976 99408
rect 417016 99368 417976 99396
rect 417016 99356 417022 99368
rect 417970 99356 417976 99368
rect 418028 99356 418034 99408
rect 436554 99356 436560 99408
rect 436612 99396 436618 99408
rect 438118 99396 438124 99408
rect 436612 99368 438124 99396
rect 436612 99356 436618 99368
rect 438118 99356 438124 99368
rect 438176 99356 438182 99408
rect 458726 99356 458732 99408
rect 458784 99396 458790 99408
rect 459462 99396 459468 99408
rect 458784 99368 459468 99396
rect 458784 99356 458790 99368
rect 459462 99356 459468 99368
rect 459520 99356 459526 99408
rect 459646 99356 459652 99408
rect 459704 99396 459710 99408
rect 460842 99396 460848 99408
rect 459704 99368 460848 99396
rect 459704 99356 459710 99368
rect 460842 99356 460848 99368
rect 460900 99356 460906 99408
rect 461302 99356 461308 99408
rect 461360 99396 461366 99408
rect 462222 99396 462228 99408
rect 461360 99368 462228 99396
rect 461360 99356 461366 99368
rect 462222 99356 462228 99368
rect 462280 99356 462286 99408
rect 463878 99356 463884 99408
rect 463936 99396 463942 99408
rect 464890 99396 464896 99408
rect 463936 99368 464896 99396
rect 463936 99356 463942 99368
rect 464890 99356 464896 99368
rect 464948 99356 464954 99408
rect 477494 99356 477500 99408
rect 477552 99396 477558 99408
rect 478782 99396 478788 99408
rect 477552 99368 478788 99396
rect 477552 99356 477558 99368
rect 478782 99356 478788 99368
rect 478840 99356 478846 99408
rect 479242 99356 479248 99408
rect 479300 99396 479306 99408
rect 480162 99396 480168 99408
rect 479300 99368 480168 99396
rect 479300 99356 479306 99368
rect 480162 99356 480168 99368
rect 480220 99356 480226 99408
rect 481818 99356 481824 99408
rect 481876 99396 481882 99408
rect 482922 99396 482928 99408
rect 481876 99368 482928 99396
rect 481876 99356 481882 99368
rect 482922 99356 482928 99368
rect 482980 99356 482986 99408
rect 483474 99356 483480 99408
rect 483532 99396 483538 99408
rect 484302 99396 484308 99408
rect 483532 99368 484308 99396
rect 483532 99356 483538 99368
rect 484302 99356 484308 99368
rect 484360 99356 484366 99408
rect 484394 99356 484400 99408
rect 484452 99396 484458 99408
rect 485682 99396 485688 99408
rect 484452 99368 485688 99396
rect 484452 99356 484458 99368
rect 485682 99356 485688 99368
rect 485740 99356 485746 99408
rect 486050 99356 486056 99408
rect 486108 99396 486114 99408
rect 486970 99396 486976 99408
rect 486108 99368 486976 99396
rect 486108 99356 486114 99368
rect 486970 99356 486976 99368
rect 487028 99356 487034 99408
rect 488626 99356 488632 99408
rect 488684 99396 488690 99408
rect 489730 99396 489736 99408
rect 488684 99368 489736 99396
rect 488684 99356 488690 99368
rect 489730 99356 489736 99368
rect 489788 99356 489794 99408
rect 490374 99356 490380 99408
rect 490432 99396 490438 99408
rect 491938 99396 491944 99408
rect 490432 99368 491944 99396
rect 490432 99356 490438 99368
rect 491938 99356 491944 99368
rect 491996 99356 492002 99408
rect 492858 99356 492864 99408
rect 492916 99396 492922 99408
rect 493870 99396 493876 99408
rect 492916 99368 493876 99396
rect 492916 99356 492922 99368
rect 493870 99356 493876 99368
rect 493928 99356 493934 99408
rect 494606 99356 494612 99408
rect 494664 99396 494670 99408
rect 495342 99396 495348 99408
rect 494664 99368 495348 99396
rect 494664 99356 494670 99368
rect 495342 99356 495348 99368
rect 495400 99356 495406 99408
rect 495434 99356 495440 99408
rect 495492 99396 495498 99408
rect 496630 99396 496636 99408
rect 495492 99368 496636 99396
rect 495492 99356 495498 99368
rect 496630 99356 496636 99368
rect 496688 99356 496694 99408
rect 497182 99356 497188 99408
rect 497240 99396 497246 99408
rect 498102 99396 498108 99408
rect 497240 99368 498108 99396
rect 497240 99356 497246 99368
rect 498102 99356 498108 99368
rect 498160 99356 498166 99408
rect 499758 99356 499764 99408
rect 499816 99396 499822 99408
rect 500862 99396 500868 99408
rect 499816 99368 500868 99396
rect 499816 99356 499822 99368
rect 500862 99356 500868 99368
rect 500920 99356 500926 99408
rect 390462 99260 390468 99272
rect 390388 99232 390468 99260
rect 390462 99220 390468 99232
rect 390520 99220 390526 99272
rect 399846 98676 399852 98728
rect 399904 98716 399910 98728
rect 442994 98716 443000 98728
rect 399904 98688 443000 98716
rect 399904 98676 399910 98688
rect 442994 98676 443000 98688
rect 443052 98676 443058 98728
rect 52362 98608 52368 98660
rect 52420 98648 52426 98660
rect 88242 98648 88248 98660
rect 52420 98620 88248 98648
rect 52420 98608 52426 98620
rect 88242 98608 88248 98620
rect 88300 98608 88306 98660
rect 336642 98608 336648 98660
rect 336700 98648 336706 98660
rect 354674 98648 354680 98660
rect 336700 98620 354680 98648
rect 336700 98608 336706 98620
rect 354674 98608 354680 98620
rect 354732 98608 354738 98660
rect 367462 98608 367468 98660
rect 367520 98648 367526 98660
rect 397454 98648 397460 98660
rect 367520 98620 397460 98648
rect 367520 98608 367526 98620
rect 397454 98608 397460 98620
rect 397512 98608 397518 98660
rect 427998 98608 428004 98660
rect 428056 98648 428062 98660
rect 429102 98648 429108 98660
rect 428056 98620 429108 98648
rect 428056 98608 428062 98620
rect 429102 98608 429108 98620
rect 429160 98608 429166 98660
rect 441706 98608 441712 98660
rect 441764 98648 441770 98660
rect 500954 98648 500960 98660
rect 441764 98620 500960 98648
rect 441764 98608 441770 98620
rect 500954 98608 500960 98620
rect 501012 98608 501018 98660
rect 194594 97928 194600 97980
rect 194652 97968 194658 97980
rect 195606 97968 195612 97980
rect 194652 97940 195612 97968
rect 194652 97928 194658 97940
rect 195606 97928 195612 97940
rect 195664 97928 195670 97980
rect 372614 97316 372620 97368
rect 372672 97316 372678 97368
rect 56502 97248 56508 97300
rect 56560 97288 56566 97300
rect 121546 97288 121552 97300
rect 56560 97260 121552 97288
rect 56560 97248 56566 97260
rect 121546 97248 121552 97260
rect 121604 97248 121610 97300
rect 349522 97248 349528 97300
rect 349580 97288 349586 97300
rect 372632 97288 372660 97316
rect 404354 97288 404360 97300
rect 349580 97260 366680 97288
rect 372632 97260 404360 97288
rect 349580 97248 349586 97260
rect 366652 97220 366680 97260
rect 404354 97248 404360 97260
rect 404412 97248 404418 97300
rect 454494 97248 454500 97300
rect 454552 97288 454558 97300
rect 518894 97288 518900 97300
rect 454552 97260 518900 97288
rect 454552 97248 454558 97260
rect 518894 97248 518900 97260
rect 518952 97248 518958 97300
rect 372614 97220 372620 97232
rect 366652 97192 372620 97220
rect 372614 97180 372620 97192
rect 372672 97180 372678 97232
rect 218330 96840 218336 96892
rect 218388 96880 218394 96892
rect 218882 96880 218888 96892
rect 218388 96852 218888 96880
rect 218388 96840 218394 96852
rect 218882 96840 218888 96852
rect 218940 96840 218946 96892
rect 211430 96704 211436 96756
rect 211488 96744 211494 96756
rect 212074 96744 212080 96756
rect 211488 96716 212080 96744
rect 211488 96704 211494 96716
rect 212074 96704 212080 96716
rect 212132 96704 212138 96756
rect 356882 96636 356888 96688
rect 356940 96676 356946 96688
rect 356974 96676 356980 96688
rect 356940 96648 356980 96676
rect 356940 96636 356946 96648
rect 356974 96636 356980 96648
rect 357032 96636 357038 96688
rect 468754 96636 468760 96688
rect 468812 96676 468818 96688
rect 468846 96676 468852 96688
rect 468812 96648 468852 96676
rect 468812 96636 468818 96648
rect 468846 96636 468852 96648
rect 468904 96636 468910 96688
rect 172885 96611 172943 96617
rect 172885 96577 172897 96611
rect 172931 96608 172943 96611
rect 173158 96608 173164 96620
rect 172931 96580 173164 96608
rect 172931 96577 172943 96580
rect 172885 96571 172943 96577
rect 173158 96568 173164 96580
rect 173216 96568 173222 96620
rect 178129 96611 178187 96617
rect 178129 96577 178141 96611
rect 178175 96608 178187 96611
rect 178402 96608 178408 96620
rect 178175 96580 178408 96608
rect 178175 96577 178187 96580
rect 178129 96571 178187 96577
rect 178402 96568 178408 96580
rect 178460 96568 178466 96620
rect 208670 96568 208676 96620
rect 208728 96608 208734 96620
rect 208854 96608 208860 96620
rect 208728 96580 208860 96608
rect 208728 96568 208734 96580
rect 208854 96568 208860 96580
rect 208912 96568 208918 96620
rect 328178 96568 328184 96620
rect 328236 96608 328242 96620
rect 328270 96608 328276 96620
rect 328236 96580 328276 96608
rect 328236 96568 328242 96580
rect 328270 96568 328276 96580
rect 328328 96568 328334 96620
rect 468846 96540 468852 96552
rect 468807 96512 468852 96540
rect 468846 96500 468852 96512
rect 468904 96500 468910 96552
rect 73062 95888 73068 95940
rect 73120 95928 73126 95940
rect 134334 95928 134340 95940
rect 73120 95900 134340 95928
rect 73120 95888 73126 95900
rect 134334 95888 134340 95900
rect 134392 95888 134398 95940
rect 354490 95888 354496 95940
rect 354548 95928 354554 95940
rect 379514 95928 379520 95940
rect 354548 95900 379520 95928
rect 354548 95888 354554 95900
rect 379514 95888 379520 95900
rect 379572 95888 379578 95940
rect 385310 95888 385316 95940
rect 385368 95928 385374 95940
rect 422294 95928 422300 95940
rect 385368 95900 422300 95928
rect 385368 95888 385374 95900
rect 422294 95888 422300 95900
rect 422352 95888 422358 95940
rect 457070 95888 457076 95940
rect 457128 95928 457134 95940
rect 521654 95928 521660 95940
rect 457128 95900 521660 95928
rect 457128 95888 457134 95900
rect 521654 95888 521660 95900
rect 521712 95888 521718 95940
rect 320450 95276 320456 95328
rect 320508 95316 320514 95328
rect 321462 95316 321468 95328
rect 320508 95288 321468 95316
rect 320508 95276 320514 95288
rect 321462 95276 321468 95288
rect 321520 95276 321526 95328
rect 164418 95208 164424 95260
rect 164476 95248 164482 95260
rect 165154 95248 165160 95260
rect 164476 95220 165160 95248
rect 164476 95208 164482 95220
rect 165154 95208 165160 95220
rect 165212 95208 165218 95260
rect 215570 95208 215576 95260
rect 215628 95248 215634 95260
rect 216306 95248 216312 95260
rect 215628 95220 216312 95248
rect 215628 95208 215634 95220
rect 216306 95208 216312 95220
rect 216364 95208 216370 95260
rect 230842 95208 230848 95260
rect 230900 95248 230906 95260
rect 231670 95248 231676 95260
rect 230900 95220 231676 95248
rect 230900 95208 230906 95220
rect 231670 95208 231676 95220
rect 231728 95208 231734 95260
rect 255866 95208 255872 95260
rect 255924 95248 255930 95260
rect 256418 95248 256424 95260
rect 255924 95220 256424 95248
rect 255924 95208 255930 95220
rect 256418 95208 256424 95220
rect 256476 95208 256482 95260
rect 258350 95208 258356 95260
rect 258408 95248 258414 95260
rect 258994 95248 259000 95260
rect 258408 95220 259000 95248
rect 258408 95208 258414 95220
rect 258994 95208 259000 95220
rect 259052 95208 259058 95260
rect 321186 95208 321192 95260
rect 321244 95248 321250 95260
rect 321370 95248 321376 95260
rect 321244 95220 321376 95248
rect 321244 95208 321250 95220
rect 321370 95208 321376 95220
rect 321428 95208 321434 95260
rect 407574 95208 407580 95260
rect 407632 95248 407638 95260
rect 408218 95248 408224 95260
rect 407632 95220 408224 95248
rect 407632 95208 407638 95220
rect 408218 95208 408224 95220
rect 408276 95208 408282 95260
rect 410886 95208 410892 95260
rect 410944 95248 410950 95260
rect 411070 95248 411076 95260
rect 410944 95220 411076 95248
rect 410944 95208 410950 95220
rect 411070 95208 411076 95220
rect 411128 95208 411134 95260
rect 428826 95208 428832 95260
rect 428884 95248 428890 95260
rect 429010 95248 429016 95260
rect 428884 95220 429016 95248
rect 428884 95208 428890 95220
rect 429010 95208 429016 95220
rect 429068 95208 429074 95260
rect 408218 95112 408224 95124
rect 408179 95084 408224 95112
rect 408218 95072 408224 95084
rect 408276 95072 408282 95124
rect 92474 94528 92480 94580
rect 92532 94568 92538 94580
rect 93118 94568 93124 94580
rect 92532 94540 93124 94568
rect 92532 94528 92538 94540
rect 93118 94528 93124 94540
rect 93176 94528 93182 94580
rect 99374 94528 99380 94580
rect 99432 94568 99438 94580
rect 99926 94568 99932 94580
rect 99432 94540 99932 94568
rect 99432 94528 99438 94540
rect 99926 94528 99932 94540
rect 99984 94528 99990 94580
rect 114554 94528 114560 94580
rect 114612 94568 114618 94580
rect 115198 94568 115204 94580
rect 114612 94540 115204 94568
rect 114612 94528 114618 94540
rect 115198 94528 115204 94540
rect 115256 94528 115262 94580
rect 117314 94528 117320 94580
rect 117372 94568 117378 94580
rect 117774 94568 117780 94580
rect 117372 94540 117780 94568
rect 117372 94528 117378 94540
rect 117774 94528 117780 94540
rect 117832 94528 117838 94580
rect 122834 94528 122840 94580
rect 122892 94568 122898 94580
rect 123846 94568 123852 94580
rect 122892 94540 123852 94568
rect 122892 94528 122898 94540
rect 123846 94528 123852 94540
rect 123904 94528 123910 94580
rect 125594 94528 125600 94580
rect 125652 94568 125658 94580
rect 126422 94568 126428 94580
rect 125652 94540 126428 94568
rect 125652 94528 125658 94540
rect 126422 94528 126428 94540
rect 126480 94528 126486 94580
rect 132494 94528 132500 94580
rect 132552 94568 132558 94580
rect 133230 94568 133236 94580
rect 132552 94540 133236 94568
rect 132552 94528 132558 94540
rect 133230 94528 133236 94540
rect 133288 94528 133294 94580
rect 135254 94528 135260 94580
rect 135312 94568 135318 94580
rect 135806 94568 135812 94580
rect 135312 94540 135812 94568
rect 135312 94528 135318 94540
rect 135806 94528 135812 94540
rect 135864 94528 135870 94580
rect 139394 94528 139400 94580
rect 139452 94568 139458 94580
rect 140038 94568 140044 94580
rect 139452 94540 140044 94568
rect 139452 94528 139458 94540
rect 140038 94528 140044 94540
rect 140096 94528 140102 94580
rect 140774 94528 140780 94580
rect 140832 94568 140838 94580
rect 141694 94568 141700 94580
rect 140832 94540 141700 94568
rect 140832 94528 140838 94540
rect 141694 94528 141700 94540
rect 141752 94528 141758 94580
rect 146294 94528 146300 94580
rect 146352 94568 146358 94580
rect 146846 94568 146852 94580
rect 146352 94540 146852 94568
rect 146352 94528 146358 94540
rect 146846 94528 146852 94540
rect 146904 94528 146910 94580
rect 150434 94528 150440 94580
rect 150492 94568 150498 94580
rect 151078 94568 151084 94580
rect 150492 94540 151084 94568
rect 150492 94528 150498 94540
rect 151078 94528 151084 94540
rect 151136 94528 151142 94580
rect 168374 94528 168380 94580
rect 168432 94568 168438 94580
rect 169110 94568 169116 94580
rect 168432 94540 169116 94568
rect 168432 94528 168438 94540
rect 169110 94528 169116 94540
rect 169168 94528 169174 94580
rect 182174 94528 182180 94580
rect 182232 94568 182238 94580
rect 182726 94568 182732 94580
rect 182232 94540 182732 94568
rect 182232 94528 182238 94540
rect 182726 94528 182732 94540
rect 182784 94528 182790 94580
rect 197354 94528 197360 94580
rect 197412 94568 197418 94580
rect 197998 94568 198004 94580
rect 197412 94540 198004 94568
rect 197412 94528 197418 94540
rect 197998 94528 198004 94540
rect 198056 94528 198062 94580
rect 222194 94528 222200 94580
rect 222252 94568 222258 94580
rect 222838 94568 222844 94580
rect 222252 94540 222844 94568
rect 222252 94528 222258 94540
rect 222838 94528 222844 94540
rect 222896 94528 222902 94580
rect 233326 94528 233332 94580
rect 233384 94568 233390 94580
rect 233878 94568 233884 94580
rect 233384 94540 233884 94568
rect 233384 94528 233390 94540
rect 233878 94528 233884 94540
rect 233936 94528 233942 94580
rect 236086 94528 236092 94580
rect 236144 94568 236150 94580
rect 236454 94568 236460 94580
rect 236144 94540 236460 94568
rect 236144 94528 236150 94540
rect 236454 94528 236460 94540
rect 236512 94528 236518 94580
rect 237374 94528 237380 94580
rect 237432 94568 237438 94580
rect 238110 94568 238116 94580
rect 237432 94540 238116 94568
rect 237432 94528 237438 94540
rect 238110 94528 238116 94540
rect 238168 94528 238174 94580
rect 240134 94528 240140 94580
rect 240192 94568 240198 94580
rect 240686 94568 240692 94580
rect 240192 94540 240692 94568
rect 240192 94528 240198 94540
rect 240686 94528 240692 94540
rect 240744 94528 240750 94580
rect 247034 94528 247040 94580
rect 247092 94568 247098 94580
rect 247678 94568 247684 94580
rect 247092 94540 247684 94568
rect 247092 94528 247098 94540
rect 247678 94528 247684 94540
rect 247736 94528 247742 94580
rect 264974 94528 264980 94580
rect 265032 94568 265038 94580
rect 265526 94568 265532 94580
rect 265032 94540 265532 94568
rect 265032 94528 265038 94540
rect 265526 94528 265532 94540
rect 265584 94528 265590 94580
rect 276014 94528 276020 94580
rect 276072 94568 276078 94580
rect 276566 94568 276572 94580
rect 276072 94540 276572 94568
rect 276072 94528 276078 94540
rect 276566 94528 276572 94540
rect 276624 94528 276630 94580
rect 13722 94460 13728 94512
rect 13780 94500 13786 94512
rect 90818 94500 90824 94512
rect 13780 94472 90824 94500
rect 13780 94460 13786 94472
rect 90818 94460 90824 94472
rect 90876 94460 90882 94512
rect 378502 94460 378508 94512
rect 378560 94500 378566 94512
rect 412634 94500 412640 94512
rect 378560 94472 412640 94500
rect 378560 94460 378566 94472
rect 412634 94460 412640 94472
rect 412692 94460 412698 94512
rect 414382 94460 414388 94512
rect 414440 94500 414446 94512
rect 462314 94500 462320 94512
rect 414440 94472 462320 94500
rect 414440 94460 414446 94472
rect 462314 94460 462320 94472
rect 462372 94460 462378 94512
rect 462406 94460 462412 94512
rect 462464 94500 462470 94512
rect 528554 94500 528560 94512
rect 462464 94472 528560 94500
rect 462464 94460 462470 94472
rect 528554 94460 528560 94472
rect 528612 94460 528618 94512
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 19978 93820 19984 93832
rect 3476 93792 19984 93820
rect 3476 93780 3482 93792
rect 19978 93780 19984 93792
rect 20036 93780 20042 93832
rect 251453 93823 251511 93829
rect 251453 93789 251465 93823
rect 251499 93820 251511 93823
rect 251542 93820 251548 93832
rect 251499 93792 251548 93820
rect 251499 93789 251511 93792
rect 251453 93783 251511 93789
rect 251542 93780 251548 93792
rect 251600 93780 251606 93832
rect 258261 93823 258319 93829
rect 258261 93789 258273 93823
rect 258307 93820 258319 93823
rect 258350 93820 258356 93832
rect 258307 93792 258356 93820
rect 258307 93789 258319 93792
rect 258261 93783 258319 93789
rect 258350 93780 258356 93792
rect 258408 93780 258414 93832
rect 22002 93100 22008 93152
rect 22060 93140 22066 93152
rect 97166 93140 97172 93152
rect 22060 93112 97172 93140
rect 22060 93100 22066 93112
rect 97166 93100 97172 93112
rect 97224 93100 97230 93152
rect 467650 93100 467656 93152
rect 467708 93140 467714 93152
rect 536834 93140 536840 93152
rect 467708 93112 536840 93140
rect 467708 93100 467714 93112
rect 536834 93100 536840 93112
rect 536892 93100 536898 93152
rect 415026 92460 415032 92472
rect 414987 92432 415032 92460
rect 415026 92420 415032 92432
rect 415084 92420 415090 92472
rect 422110 92460 422116 92472
rect 422071 92432 422116 92460
rect 422110 92420 422116 92432
rect 422168 92420 422174 92472
rect 179414 92352 179420 92404
rect 179472 92392 179478 92404
rect 180150 92392 180156 92404
rect 179472 92364 180156 92392
rect 179472 92352 179478 92364
rect 180150 92352 180156 92364
rect 180208 92352 180214 92404
rect 244274 92352 244280 92404
rect 244332 92392 244338 92404
rect 245102 92392 245108 92404
rect 244332 92364 245108 92392
rect 244332 92352 244338 92364
rect 245102 92352 245108 92364
rect 245160 92352 245166 92404
rect 262214 92352 262220 92404
rect 262272 92392 262278 92404
rect 262950 92392 262956 92404
rect 262272 92364 262956 92392
rect 262272 92352 262278 92364
rect 262950 92352 262956 92364
rect 263008 92352 263014 92404
rect 273254 92352 273260 92404
rect 273312 92392 273318 92404
rect 273990 92392 273996 92404
rect 273312 92364 273996 92392
rect 273312 92352 273318 92364
rect 273990 92352 273996 92364
rect 274048 92352 274054 92404
rect 88242 91740 88248 91792
rect 88300 91780 88306 91792
rect 144086 91780 144092 91792
rect 88300 91752 144092 91780
rect 88300 91740 88306 91752
rect 144086 91740 144092 91752
rect 144144 91740 144150 91792
rect 475930 91740 475936 91792
rect 475988 91780 475994 91792
rect 546586 91780 546592 91792
rect 475988 91752 546592 91780
rect 475988 91740 475994 91752
rect 546586 91740 546592 91752
rect 546644 91740 546650 91792
rect 270494 91536 270500 91588
rect 270552 91576 270558 91588
rect 271414 91576 271420 91588
rect 270552 91548 271420 91576
rect 270552 91536 270558 91548
rect 271414 91536 271420 91548
rect 271472 91536 271478 91588
rect 259454 91264 259460 91316
rect 259512 91304 259518 91316
rect 260374 91304 260380 91316
rect 259512 91276 260380 91304
rect 259512 91264 259518 91276
rect 260374 91264 260380 91276
rect 260432 91264 260438 91316
rect 27522 90312 27528 90364
rect 27580 90352 27586 90364
rect 100846 90352 100852 90364
rect 27580 90324 100852 90352
rect 27580 90312 27586 90324
rect 100846 90312 100852 90324
rect 100904 90312 100910 90364
rect 139302 90312 139308 90364
rect 139360 90352 139366 90364
rect 180794 90352 180800 90364
rect 139360 90324 180800 90352
rect 139360 90312 139366 90324
rect 180794 90312 180800 90324
rect 180852 90312 180858 90364
rect 400030 90312 400036 90364
rect 400088 90352 400094 90364
rect 441614 90352 441620 90364
rect 400088 90324 441620 90352
rect 400088 90312 400094 90324
rect 441614 90312 441620 90324
rect 441672 90312 441678 90364
rect 480070 90312 480076 90364
rect 480128 90352 480134 90364
rect 554774 90352 554780 90364
rect 480128 90324 554780 90352
rect 480128 90312 480134 90324
rect 554774 90312 554780 90324
rect 554832 90312 554838 90364
rect 175550 89808 175556 89820
rect 175476 89780 175556 89808
rect 175476 89752 175504 89780
rect 175550 89768 175556 89780
rect 175608 89768 175614 89820
rect 118786 89700 118792 89752
rect 118844 89740 118850 89752
rect 119522 89740 119528 89752
rect 118844 89712 119528 89740
rect 118844 89700 118850 89712
rect 119522 89700 119528 89712
rect 119580 89700 119586 89752
rect 129734 89700 129740 89752
rect 129792 89740 129798 89752
rect 130378 89740 130384 89752
rect 129792 89712 130384 89740
rect 129792 89700 129798 89712
rect 130378 89700 130384 89712
rect 130436 89700 130442 89752
rect 158898 89700 158904 89752
rect 158956 89740 158962 89752
rect 159634 89740 159640 89752
rect 158956 89712 159640 89740
rect 158956 89700 158962 89712
rect 159634 89700 159640 89712
rect 159692 89700 159698 89752
rect 160094 89700 160100 89752
rect 160152 89700 160158 89752
rect 165706 89700 165712 89752
rect 165764 89740 165770 89752
rect 166350 89740 166356 89752
rect 165764 89712 166356 89740
rect 165764 89700 165770 89712
rect 166350 89700 166356 89712
rect 166408 89700 166414 89752
rect 169938 89700 169944 89752
rect 169996 89740 170002 89752
rect 170398 89740 170404 89752
rect 169996 89712 170404 89740
rect 169996 89700 170002 89712
rect 170398 89700 170404 89712
rect 170456 89700 170462 89752
rect 175458 89700 175464 89752
rect 175516 89700 175522 89752
rect 332318 89700 332324 89752
rect 332376 89740 332382 89752
rect 332502 89740 332508 89752
rect 332376 89712 332508 89740
rect 332376 89700 332382 89712
rect 332502 89700 332508 89712
rect 332560 89700 332566 89752
rect 379238 89700 379244 89752
rect 379296 89740 379302 89752
rect 379422 89740 379428 89752
rect 379296 89712 379428 89740
rect 379296 89700 379302 89712
rect 379422 89700 379428 89712
rect 379480 89700 379486 89752
rect 450998 89700 451004 89752
rect 451056 89740 451062 89752
rect 451182 89740 451188 89752
rect 451056 89712 451188 89740
rect 451056 89700 451062 89712
rect 451182 89700 451188 89712
rect 451240 89700 451246 89752
rect 160112 89604 160140 89700
rect 172882 89672 172888 89684
rect 172843 89644 172888 89672
rect 172882 89632 172888 89644
rect 172940 89632 172946 89684
rect 468849 89675 468907 89681
rect 468849 89641 468861 89675
rect 468895 89672 468907 89675
rect 469030 89672 469036 89684
rect 468895 89644 469036 89672
rect 468895 89641 468907 89644
rect 468849 89635 468907 89641
rect 469030 89632 469036 89644
rect 469088 89632 469094 89684
rect 160186 89604 160192 89616
rect 160112 89576 160192 89604
rect 160186 89564 160192 89576
rect 160244 89564 160250 89616
rect 34422 88952 34428 89004
rect 34480 88992 34486 89004
rect 105538 88992 105544 89004
rect 34480 88964 105544 88992
rect 34480 88952 34486 88964
rect 105538 88952 105544 88964
rect 105596 88952 105602 89004
rect 397362 88952 397368 89004
rect 397420 88992 397426 89004
rect 437474 88992 437480 89004
rect 397420 88964 437480 88992
rect 397420 88952 397426 88964
rect 437474 88952 437480 88964
rect 437532 88952 437538 89004
rect 482830 88952 482836 89004
rect 482888 88992 482894 89004
rect 557534 88992 557540 89004
rect 482888 88964 557540 88992
rect 482888 88952 482894 88964
rect 557534 88952 557540 88964
rect 557592 88952 557598 89004
rect 504634 88272 504640 88324
rect 504692 88312 504698 88324
rect 580166 88312 580172 88324
rect 504692 88284 580172 88312
rect 504692 88272 504698 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 38562 87592 38568 87644
rect 38620 87632 38626 87644
rect 108298 87632 108304 87644
rect 38620 87604 108304 87632
rect 38620 87592 38626 87604
rect 108298 87592 108304 87604
rect 108356 87592 108362 87644
rect 218330 87156 218336 87168
rect 218256 87128 218336 87156
rect 178126 87088 178132 87100
rect 178087 87060 178132 87088
rect 178126 87048 178132 87060
rect 178184 87048 178190 87100
rect 218256 87032 218284 87128
rect 218330 87116 218336 87128
rect 218388 87116 218394 87168
rect 95602 86980 95608 87032
rect 95660 86980 95666 87032
rect 218238 86980 218244 87032
rect 218296 86980 218302 87032
rect 224862 86980 224868 87032
rect 224920 87020 224926 87032
rect 225322 87020 225328 87032
rect 224920 86992 225328 87020
rect 224920 86980 224926 86992
rect 225322 86980 225328 86992
rect 225380 86980 225386 87032
rect 230842 87020 230848 87032
rect 230803 86992 230848 87020
rect 230842 86980 230848 86992
rect 230900 86980 230906 87032
rect 248874 86980 248880 87032
rect 248932 87020 248938 87032
rect 248966 87020 248972 87032
rect 248932 86992 248972 87020
rect 248932 86980 248938 86992
rect 248966 86980 248972 86992
rect 249024 86980 249030 87032
rect 86126 86952 86132 86964
rect 86087 86924 86132 86952
rect 86126 86912 86132 86924
rect 86184 86912 86190 86964
rect 88518 86952 88524 86964
rect 88479 86924 88524 86952
rect 88518 86912 88524 86924
rect 88576 86912 88582 86964
rect 95620 86884 95648 86980
rect 110509 86955 110567 86961
rect 110509 86921 110521 86955
rect 110555 86952 110567 86955
rect 110598 86952 110604 86964
rect 110555 86924 110604 86952
rect 110555 86921 110567 86924
rect 110509 86915 110567 86921
rect 110598 86912 110604 86924
rect 110656 86912 110662 86964
rect 124217 86955 124275 86961
rect 124217 86921 124229 86955
rect 124263 86952 124275 86955
rect 124306 86952 124312 86964
rect 124263 86924 124312 86952
rect 124263 86921 124275 86924
rect 124217 86915 124275 86921
rect 124306 86912 124312 86924
rect 124364 86912 124370 86964
rect 129829 86955 129887 86961
rect 129829 86921 129841 86955
rect 129875 86952 129887 86955
rect 129918 86952 129924 86964
rect 129875 86924 129924 86952
rect 129875 86921 129887 86924
rect 129829 86915 129887 86921
rect 129918 86912 129924 86924
rect 129976 86912 129982 86964
rect 142157 86955 142215 86961
rect 142157 86921 142169 86955
rect 142203 86952 142215 86955
rect 142246 86952 142252 86964
rect 142203 86924 142252 86952
rect 142203 86921 142215 86924
rect 142157 86915 142215 86921
rect 142246 86912 142252 86924
rect 142304 86912 142310 86964
rect 184014 86952 184020 86964
rect 183975 86924 184020 86952
rect 184014 86912 184020 86924
rect 184072 86912 184078 86964
rect 195977 86955 196035 86961
rect 195977 86921 195989 86955
rect 196023 86952 196035 86955
rect 196066 86952 196072 86964
rect 196023 86924 196072 86952
rect 196023 86921 196035 86924
rect 195977 86915 196035 86921
rect 196066 86912 196072 86924
rect 196124 86912 196130 86964
rect 200298 86952 200304 86964
rect 200259 86924 200304 86952
rect 200298 86912 200304 86924
rect 200356 86912 200362 86964
rect 252649 86955 252707 86961
rect 252649 86921 252661 86955
rect 252695 86952 252707 86955
rect 252738 86952 252744 86964
rect 252695 86924 252744 86952
rect 252695 86921 252707 86924
rect 252649 86915 252707 86921
rect 252738 86912 252744 86924
rect 252796 86912 252802 86964
rect 290001 86955 290059 86961
rect 290001 86921 290013 86955
rect 290047 86952 290059 86955
rect 290090 86952 290096 86964
rect 290047 86924 290096 86952
rect 290047 86921 290059 86924
rect 290001 86915 290059 86921
rect 290090 86912 290096 86924
rect 290148 86912 290154 86964
rect 310146 86952 310152 86964
rect 310107 86924 310152 86952
rect 310146 86912 310152 86924
rect 310204 86912 310210 86964
rect 95694 86884 95700 86896
rect 95620 86856 95700 86884
rect 95694 86844 95700 86856
rect 95752 86844 95758 86896
rect 49602 86232 49608 86284
rect 49660 86272 49666 86284
rect 117406 86272 117412 86284
rect 49660 86244 117412 86272
rect 49660 86232 49666 86244
rect 117406 86232 117412 86244
rect 117464 86232 117470 86284
rect 491938 86232 491944 86284
rect 491996 86272 492002 86284
rect 568574 86272 568580 86284
rect 491996 86244 568580 86272
rect 491996 86232 492002 86244
rect 568574 86232 568580 86244
rect 568632 86232 568638 86284
rect 229278 85552 229284 85604
rect 229336 85592 229342 85604
rect 229646 85592 229652 85604
rect 229336 85564 229652 85592
rect 229336 85552 229342 85564
rect 229646 85552 229652 85564
rect 229704 85552 229710 85604
rect 230842 85592 230848 85604
rect 230803 85564 230848 85592
rect 230842 85552 230848 85564
rect 230900 85552 230906 85604
rect 284570 85552 284576 85604
rect 284628 85592 284634 85604
rect 284754 85592 284760 85604
rect 284628 85564 284760 85592
rect 284628 85552 284634 85564
rect 284754 85552 284760 85564
rect 284812 85552 284818 85604
rect 321186 85552 321192 85604
rect 321244 85592 321250 85604
rect 321278 85592 321284 85604
rect 321244 85564 321284 85592
rect 321244 85552 321250 85564
rect 321278 85552 321284 85564
rect 321336 85552 321342 85604
rect 408218 85592 408224 85604
rect 408179 85564 408224 85592
rect 408218 85552 408224 85564
rect 408276 85552 408282 85604
rect 428826 85552 428832 85604
rect 428884 85592 428890 85604
rect 428918 85592 428924 85604
rect 428884 85564 428924 85592
rect 428884 85552 428890 85564
rect 428918 85552 428924 85564
rect 428976 85552 428982 85604
rect 160186 85524 160192 85536
rect 160147 85496 160192 85524
rect 160186 85484 160192 85496
rect 160244 85484 160250 85536
rect 164418 85524 164424 85536
rect 164379 85496 164424 85524
rect 164418 85484 164424 85496
rect 164476 85484 164482 85536
rect 169938 85524 169944 85536
rect 169899 85496 169944 85524
rect 169938 85484 169944 85496
rect 169996 85484 170002 85536
rect 178126 85524 178132 85536
rect 178087 85496 178132 85524
rect 178126 85484 178132 85496
rect 178184 85484 178190 85536
rect 215389 85527 215447 85533
rect 215389 85493 215401 85527
rect 215435 85524 215447 85527
rect 215478 85524 215484 85536
rect 215435 85496 215484 85524
rect 215435 85493 215447 85496
rect 215389 85487 215447 85493
rect 215478 85484 215484 85496
rect 215536 85484 215542 85536
rect 218149 85527 218207 85533
rect 218149 85493 218161 85527
rect 218195 85524 218207 85527
rect 218238 85524 218244 85536
rect 218195 85496 218244 85524
rect 218195 85493 218207 85496
rect 218149 85487 218207 85493
rect 218238 85484 218244 85496
rect 218296 85484 218302 85536
rect 224862 85524 224868 85536
rect 224823 85496 224868 85524
rect 224862 85484 224868 85496
rect 224920 85484 224926 85536
rect 226518 85524 226524 85536
rect 226479 85496 226524 85524
rect 226518 85484 226524 85496
rect 226576 85484 226582 85536
rect 426066 85484 426072 85536
rect 426124 85524 426130 85536
rect 426158 85524 426164 85536
rect 426124 85496 426164 85524
rect 426124 85484 426130 85496
rect 426158 85484 426164 85496
rect 426216 85484 426222 85536
rect 468941 85527 468999 85533
rect 468941 85493 468953 85527
rect 468987 85524 468999 85527
rect 469030 85524 469036 85536
rect 468987 85496 469036 85524
rect 468987 85493 468999 85496
rect 468941 85487 468999 85493
rect 469030 85484 469036 85496
rect 469088 85484 469094 85536
rect 53742 84804 53748 84856
rect 53800 84844 53806 84856
rect 118786 84844 118792 84856
rect 53800 84816 118792 84844
rect 53800 84804 53806 84816
rect 118786 84804 118792 84816
rect 118844 84804 118850 84856
rect 493870 84804 493876 84856
rect 493928 84844 493934 84856
rect 571426 84844 571432 84856
rect 493928 84816 571432 84844
rect 493928 84804 493934 84816
rect 571426 84804 571432 84816
rect 571484 84804 571490 84856
rect 241606 84192 241612 84244
rect 241664 84232 241670 84244
rect 241790 84232 241796 84244
rect 241664 84204 241796 84232
rect 241664 84192 241670 84204
rect 241790 84192 241796 84204
rect 241848 84192 241854 84244
rect 251450 84232 251456 84244
rect 251411 84204 251456 84232
rect 251450 84192 251456 84204
rect 251508 84192 251514 84244
rect 258258 84232 258264 84244
rect 258219 84204 258264 84232
rect 258258 84192 258264 84204
rect 258316 84192 258322 84244
rect 64782 83444 64788 83496
rect 64840 83484 64846 83496
rect 126974 83484 126980 83496
rect 64840 83456 126980 83484
rect 64840 83444 64846 83456
rect 126974 83444 126980 83456
rect 127032 83444 127038 83496
rect 438762 83444 438768 83496
rect 438820 83484 438826 83496
rect 495434 83484 495440 83496
rect 438820 83456 495440 83484
rect 438820 83444 438826 83456
rect 495434 83444 495440 83456
rect 495492 83444 495498 83496
rect 496630 83444 496636 83496
rect 496688 83484 496694 83496
rect 574738 83484 574744 83496
rect 496688 83456 574744 83484
rect 496688 83444 496694 83456
rect 574738 83444 574744 83456
rect 574796 83444 574802 83496
rect 421926 82900 421932 82952
rect 421984 82940 421990 82952
rect 422113 82943 422171 82949
rect 422113 82940 422125 82943
rect 421984 82912 422125 82940
rect 421984 82900 421990 82912
rect 422113 82909 422125 82912
rect 422159 82909 422171 82943
rect 422113 82903 422171 82909
rect 415026 82872 415032 82884
rect 414987 82844 415032 82872
rect 415026 82832 415032 82844
rect 415084 82832 415090 82884
rect 67542 82084 67548 82136
rect 67600 82124 67606 82136
rect 128998 82124 129004 82136
rect 67600 82096 129004 82124
rect 67600 82084 67606 82096
rect 128998 82084 129004 82096
rect 129056 82084 129062 82136
rect 212718 82084 212724 82136
rect 212776 82124 212782 82136
rect 213086 82124 213092 82136
rect 212776 82096 213092 82124
rect 212776 82084 212782 82096
rect 213086 82084 213092 82096
rect 213144 82084 213150 82136
rect 390186 82084 390192 82136
rect 390244 82124 390250 82136
rect 390370 82124 390376 82136
rect 390244 82096 390376 82124
rect 390244 82084 390250 82096
rect 390370 82084 390376 82096
rect 390428 82084 390434 82136
rect 453850 82084 453856 82136
rect 453908 82124 453914 82136
rect 516134 82124 516140 82136
rect 453908 82096 516140 82124
rect 453908 82084 453914 82096
rect 516134 82084 516140 82096
rect 516192 82084 516198 82136
rect 422018 81376 422024 81388
rect 421979 81348 422024 81376
rect 422018 81336 422024 81348
rect 422076 81336 422082 81388
rect 154761 80767 154819 80773
rect 154761 80733 154773 80767
rect 154807 80764 154819 80767
rect 154942 80764 154948 80776
rect 154807 80736 154948 80764
rect 154807 80733 154819 80736
rect 154761 80727 154819 80733
rect 154942 80724 154948 80736
rect 155000 80724 155006 80776
rect 172609 80767 172667 80773
rect 172609 80733 172621 80767
rect 172655 80764 172667 80767
rect 172882 80764 172888 80776
rect 172655 80736 172888 80764
rect 172655 80733 172667 80736
rect 172609 80727 172667 80733
rect 172882 80724 172888 80736
rect 172940 80724 172946 80776
rect 428642 80724 428648 80776
rect 428700 80764 428706 80776
rect 428829 80767 428887 80773
rect 428829 80764 428841 80767
rect 428700 80736 428841 80764
rect 428700 80724 428706 80736
rect 428829 80733 428841 80736
rect 428875 80733 428887 80767
rect 428829 80727 428887 80733
rect 71682 80656 71688 80708
rect 71740 80696 71746 80708
rect 132586 80696 132592 80708
rect 71740 80668 132592 80696
rect 71740 80656 71746 80668
rect 132586 80656 132592 80668
rect 132644 80656 132650 80708
rect 455322 80656 455328 80708
rect 455380 80696 455386 80708
rect 520274 80696 520280 80708
rect 455380 80668 520280 80696
rect 455380 80656 455386 80668
rect 520274 80656 520280 80668
rect 520332 80656 520338 80708
rect 205726 80180 205732 80232
rect 205784 80220 205790 80232
rect 206462 80220 206468 80232
rect 205784 80192 206468 80220
rect 205784 80180 205790 80192
rect 206462 80180 206468 80192
rect 206520 80180 206526 80232
rect 272061 80223 272119 80229
rect 272061 80189 272073 80223
rect 272107 80220 272119 80223
rect 272150 80220 272156 80232
rect 272107 80192 272156 80220
rect 272107 80189 272119 80192
rect 272061 80183 272119 80189
rect 272150 80180 272156 80192
rect 272208 80180 272214 80232
rect 287333 80223 287391 80229
rect 287333 80189 287345 80223
rect 287379 80220 287391 80223
rect 287422 80220 287428 80232
rect 287379 80192 287428 80220
rect 287379 80189 287391 80192
rect 287333 80183 287391 80189
rect 287422 80180 287428 80192
rect 287480 80180 287486 80232
rect 357066 80180 357072 80232
rect 357124 80180 357130 80232
rect 161750 80152 161756 80164
rect 161676 80124 161756 80152
rect 161676 80096 161704 80124
rect 161750 80112 161756 80124
rect 161808 80112 161814 80164
rect 248874 80152 248880 80164
rect 248835 80124 248880 80152
rect 248874 80112 248880 80124
rect 248932 80112 248938 80164
rect 350169 80155 350227 80161
rect 350169 80121 350181 80155
rect 350215 80152 350227 80155
rect 350258 80152 350264 80164
rect 350215 80124 350264 80152
rect 350215 80121 350227 80124
rect 350169 80115 350227 80121
rect 350258 80112 350264 80124
rect 350316 80112 350322 80164
rect 100754 80044 100760 80096
rect 100812 80084 100818 80096
rect 101490 80084 101496 80096
rect 100812 80056 101496 80084
rect 100812 80044 100818 80056
rect 101490 80044 101496 80056
rect 101548 80044 101554 80096
rect 147674 80044 147680 80096
rect 147732 80084 147738 80096
rect 147858 80084 147864 80096
rect 147732 80056 147864 80084
rect 147732 80044 147738 80056
rect 147858 80044 147864 80056
rect 147916 80044 147922 80096
rect 161658 80044 161664 80096
rect 161716 80044 161722 80096
rect 176654 80044 176660 80096
rect 176712 80084 176718 80096
rect 177114 80084 177120 80096
rect 176712 80056 177120 80084
rect 176712 80044 176718 80056
rect 177114 80044 177120 80056
rect 177172 80044 177178 80096
rect 327994 80044 328000 80096
rect 328052 80044 328058 80096
rect 332502 80084 332508 80096
rect 332428 80056 332508 80084
rect 3418 79976 3424 80028
rect 3476 80016 3482 80028
rect 17218 80016 17224 80028
rect 3476 79988 17224 80016
rect 3476 79976 3482 79988
rect 17218 79976 17224 79988
rect 17276 79976 17282 80028
rect 183738 79976 183744 80028
rect 183796 80016 183802 80028
rect 184017 80019 184075 80025
rect 184017 80016 184029 80019
rect 183796 79988 184029 80016
rect 183796 79976 183802 79988
rect 184017 79985 184029 79988
rect 184063 79985 184075 80019
rect 184017 79979 184075 79985
rect 310149 80019 310207 80025
rect 310149 79985 310161 80019
rect 310195 80016 310207 80019
rect 310238 80016 310244 80028
rect 310195 79988 310244 80016
rect 310195 79985 310207 79988
rect 310149 79979 310207 79985
rect 310238 79976 310244 79988
rect 310296 79976 310302 80028
rect 328012 79948 328040 80044
rect 332428 80028 332456 80056
rect 332502 80044 332508 80056
rect 332560 80044 332566 80096
rect 357084 80028 357112 80180
rect 379330 80112 379336 80164
rect 379388 80112 379394 80164
rect 379348 80028 379376 80112
rect 415026 80044 415032 80096
rect 415084 80044 415090 80096
rect 433058 80044 433064 80096
rect 433116 80084 433122 80096
rect 433242 80084 433248 80096
rect 433116 80056 433248 80084
rect 433116 80044 433122 80056
rect 433242 80044 433248 80056
rect 433300 80044 433306 80096
rect 439866 80044 439872 80096
rect 439924 80044 439930 80096
rect 332410 79976 332416 80028
rect 332468 79976 332474 80028
rect 357066 79976 357072 80028
rect 357124 79976 357130 80028
rect 379330 79976 379336 80028
rect 379388 79976 379394 80028
rect 328086 79948 328092 79960
rect 328012 79920 328092 79948
rect 328086 79908 328092 79920
rect 328144 79908 328150 79960
rect 415044 79948 415072 80044
rect 415118 79948 415124 79960
rect 415044 79920 415124 79948
rect 415118 79908 415124 79920
rect 415176 79908 415182 79960
rect 439884 79948 439912 80044
rect 439958 79948 439964 79960
rect 439884 79920 439964 79948
rect 439958 79908 439964 79920
rect 440016 79908 440022 79960
rect 17862 79296 17868 79348
rect 17920 79336 17926 79348
rect 91738 79336 91744 79348
rect 17920 79308 91744 79336
rect 17920 79296 17926 79308
rect 91738 79296 91744 79308
rect 91796 79296 91802 79348
rect 92382 79296 92388 79348
rect 92440 79336 92446 79348
rect 147766 79336 147772 79348
rect 92440 79308 147772 79336
rect 92440 79296 92446 79308
rect 147766 79296 147772 79308
rect 147824 79296 147830 79348
rect 460750 79296 460756 79348
rect 460808 79336 460814 79348
rect 527174 79336 527180 79348
rect 460808 79308 527180 79336
rect 460808 79296 460814 79308
rect 527174 79296 527180 79308
rect 527232 79296 527238 79348
rect 223666 78548 223672 78600
rect 223724 78588 223730 78600
rect 224126 78588 224132 78600
rect 223724 78560 224132 78588
rect 223724 78548 223730 78560
rect 224126 78548 224132 78560
rect 224184 78548 224190 78600
rect 74442 77936 74448 77988
rect 74500 77976 74506 77988
rect 135346 77976 135352 77988
rect 74500 77948 135352 77976
rect 74500 77936 74506 77948
rect 135346 77936 135352 77948
rect 135404 77936 135410 77988
rect 478690 77936 478696 77988
rect 478748 77976 478754 77988
rect 552014 77976 552020 77988
rect 478748 77948 552020 77976
rect 478748 77936 478754 77948
rect 552014 77936 552020 77948
rect 552072 77936 552078 77988
rect 258258 77324 258264 77376
rect 258316 77324 258322 77376
rect 284570 77364 284576 77376
rect 284404 77336 284576 77364
rect 85850 77256 85856 77308
rect 85908 77296 85914 77308
rect 86129 77299 86187 77305
rect 86129 77296 86141 77299
rect 85908 77268 86141 77296
rect 85908 77256 85914 77268
rect 86129 77265 86141 77268
rect 86175 77265 86187 77299
rect 86129 77259 86187 77265
rect 87230 77256 87236 77308
rect 87288 77296 87294 77308
rect 87598 77296 87604 77308
rect 87288 77268 87604 77296
rect 87288 77256 87294 77268
rect 87598 77256 87604 77268
rect 87656 77256 87662 77308
rect 88518 77296 88524 77308
rect 88479 77268 88524 77296
rect 88518 77256 88524 77268
rect 88576 77256 88582 77308
rect 103606 77256 103612 77308
rect 103664 77296 103670 77308
rect 104066 77296 104072 77308
rect 103664 77268 104072 77296
rect 103664 77256 103670 77268
rect 104066 77256 104072 77268
rect 104124 77256 104130 77308
rect 106274 77256 106280 77308
rect 106332 77296 106338 77308
rect 106642 77296 106648 77308
rect 106332 77268 106648 77296
rect 106332 77256 106338 77268
rect 106642 77256 106648 77268
rect 106700 77256 106706 77308
rect 110506 77296 110512 77308
rect 110467 77268 110512 77296
rect 110506 77256 110512 77268
rect 110564 77256 110570 77308
rect 111794 77256 111800 77308
rect 111852 77296 111858 77308
rect 112070 77296 112076 77308
rect 111852 77268 112076 77296
rect 111852 77256 111858 77268
rect 112070 77256 112076 77268
rect 112128 77256 112134 77308
rect 124214 77296 124220 77308
rect 124175 77268 124220 77296
rect 124214 77256 124220 77268
rect 124272 77256 124278 77308
rect 129826 77296 129832 77308
rect 129787 77268 129832 77296
rect 129826 77256 129832 77268
rect 129884 77256 129890 77308
rect 142154 77296 142160 77308
rect 142115 77268 142160 77296
rect 142154 77256 142160 77268
rect 142212 77256 142218 77308
rect 195974 77296 195980 77308
rect 195935 77268 195980 77296
rect 195974 77256 195980 77268
rect 196032 77256 196038 77308
rect 200298 77296 200304 77308
rect 200259 77268 200304 77296
rect 200298 77256 200304 77268
rect 200356 77256 200362 77308
rect 248598 77256 248604 77308
rect 248656 77296 248662 77308
rect 248877 77299 248935 77305
rect 248877 77296 248889 77299
rect 248656 77268 248889 77296
rect 248656 77256 248662 77268
rect 248877 77265 248889 77268
rect 248923 77265 248935 77299
rect 252646 77296 252652 77308
rect 252607 77268 252652 77296
rect 248877 77259 248935 77265
rect 252646 77256 252652 77268
rect 252704 77256 252710 77308
rect 258276 77240 258304 77324
rect 272058 77296 272064 77308
rect 272019 77268 272064 77296
rect 272058 77256 272064 77268
rect 272116 77256 272122 77308
rect 277578 77256 277584 77308
rect 277636 77296 277642 77308
rect 277670 77296 277676 77308
rect 277636 77268 277676 77296
rect 277636 77256 277642 77268
rect 277670 77256 277676 77268
rect 277728 77256 277734 77308
rect 278866 77256 278872 77308
rect 278924 77296 278930 77308
rect 278958 77296 278964 77308
rect 278924 77268 278964 77296
rect 278924 77256 278930 77268
rect 278958 77256 278964 77268
rect 279016 77256 279022 77308
rect 284404 77240 284432 77336
rect 284570 77324 284576 77336
rect 284628 77324 284634 77376
rect 287330 77296 287336 77308
rect 287291 77268 287336 77296
rect 287330 77256 287336 77268
rect 287388 77256 287394 77308
rect 289998 77296 290004 77308
rect 289959 77268 290004 77296
rect 289998 77256 290004 77268
rect 290056 77256 290062 77308
rect 136726 77228 136732 77240
rect 136687 77200 136732 77228
rect 136726 77188 136732 77200
rect 136784 77188 136790 77240
rect 183738 77228 183744 77240
rect 183699 77200 183744 77228
rect 183738 77188 183744 77200
rect 183796 77188 183802 77240
rect 258258 77188 258264 77240
rect 258316 77188 258322 77240
rect 284386 77188 284392 77240
rect 284444 77188 284450 77240
rect 439958 77228 439964 77240
rect 439919 77200 439964 77228
rect 439958 77188 439964 77200
rect 440016 77188 440022 77240
rect 504542 77188 504548 77240
rect 504600 77228 504606 77240
rect 580166 77228 580172 77240
rect 504600 77200 580172 77228
rect 504600 77188 504606 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 142154 77160 142160 77172
rect 142115 77132 142160 77160
rect 142154 77120 142160 77132
rect 142212 77120 142218 77172
rect 230842 76644 230848 76696
rect 230900 76644 230906 76696
rect 230860 76560 230888 76644
rect 28902 76508 28908 76560
rect 28960 76548 28966 76560
rect 100754 76548 100760 76560
rect 28960 76520 100760 76548
rect 28960 76508 28966 76520
rect 100754 76508 100760 76520
rect 100812 76508 100818 76560
rect 230842 76508 230848 76560
rect 230900 76508 230906 76560
rect 408126 75964 408132 76016
rect 408184 76004 408190 76016
rect 408218 76004 408224 76016
rect 408184 75976 408224 76004
rect 408184 75964 408190 75976
rect 408218 75964 408224 75976
rect 408276 75964 408282 76016
rect 160186 75936 160192 75948
rect 160147 75908 160192 75936
rect 160186 75896 160192 75908
rect 160244 75896 160250 75948
rect 164418 75936 164424 75948
rect 164379 75908 164424 75936
rect 164418 75896 164424 75908
rect 164476 75896 164482 75948
rect 169938 75936 169944 75948
rect 169899 75908 169944 75936
rect 169938 75896 169944 75908
rect 169996 75896 170002 75948
rect 172606 75936 172612 75948
rect 172567 75908 172612 75936
rect 172606 75896 172612 75908
rect 172664 75896 172670 75948
rect 178129 75939 178187 75945
rect 178129 75905 178141 75939
rect 178175 75936 178187 75939
rect 178402 75936 178408 75948
rect 178175 75908 178408 75936
rect 178175 75905 178187 75908
rect 178129 75899 178187 75905
rect 178402 75896 178408 75908
rect 178460 75896 178466 75948
rect 215386 75936 215392 75948
rect 215347 75908 215392 75936
rect 215386 75896 215392 75908
rect 215444 75896 215450 75948
rect 218146 75936 218152 75948
rect 218107 75908 218152 75936
rect 218146 75896 218152 75908
rect 218204 75896 218210 75948
rect 224865 75939 224923 75945
rect 224865 75905 224877 75939
rect 224911 75936 224923 75939
rect 224954 75936 224960 75948
rect 224911 75908 224960 75936
rect 224911 75905 224923 75908
rect 224865 75899 224923 75905
rect 224954 75896 224960 75908
rect 225012 75896 225018 75948
rect 226521 75939 226579 75945
rect 226521 75905 226533 75939
rect 226567 75936 226579 75939
rect 226610 75936 226616 75948
rect 226567 75908 226616 75936
rect 226567 75905 226579 75908
rect 226521 75899 226579 75905
rect 226610 75896 226616 75908
rect 226668 75896 226674 75948
rect 350166 75936 350172 75948
rect 350127 75908 350172 75936
rect 350166 75896 350172 75908
rect 350224 75896 350230 75948
rect 386138 75896 386144 75948
rect 386196 75936 386202 75948
rect 386322 75936 386328 75948
rect 386196 75908 386328 75936
rect 386196 75896 386202 75908
rect 386322 75896 386328 75908
rect 386380 75896 386386 75948
rect 327997 75871 328055 75877
rect 327997 75837 328009 75871
rect 328043 75868 328055 75871
rect 328086 75868 328092 75880
rect 328043 75840 328092 75868
rect 328043 75837 328055 75840
rect 327997 75831 328055 75837
rect 328086 75828 328092 75840
rect 328144 75828 328150 75880
rect 408126 75868 408132 75880
rect 408087 75840 408132 75868
rect 408126 75828 408132 75840
rect 408184 75828 408190 75880
rect 31665 75191 31723 75197
rect 31665 75157 31677 75191
rect 31711 75188 31723 75191
rect 103606 75188 103612 75200
rect 31711 75160 103612 75188
rect 31711 75157 31723 75160
rect 31665 75151 31723 75157
rect 103606 75148 103612 75160
rect 103664 75148 103670 75200
rect 486970 75148 486976 75200
rect 487028 75188 487034 75200
rect 563146 75188 563152 75200
rect 487028 75160 563152 75188
rect 487028 75148 487034 75160
rect 563146 75148 563152 75160
rect 563204 75148 563210 75200
rect 95513 74511 95571 74517
rect 95513 74477 95525 74511
rect 95559 74508 95571 74511
rect 95786 74508 95792 74520
rect 95559 74480 95792 74508
rect 95559 74477 95571 74480
rect 95513 74471 95571 74477
rect 95786 74468 95792 74480
rect 95844 74468 95850 74520
rect 410886 74508 410892 74520
rect 410847 74480 410892 74508
rect 410886 74468 410892 74480
rect 410944 74468 410950 74520
rect 42702 73788 42708 73840
rect 42760 73828 42766 73840
rect 106918 73828 106924 73840
rect 42760 73800 106924 73828
rect 42760 73788 42766 73800
rect 106918 73788 106924 73800
rect 106976 73788 106982 73840
rect 342070 73788 342076 73840
rect 342128 73828 342134 73840
rect 361574 73828 361580 73840
rect 342128 73800 361580 73828
rect 342128 73788 342134 73800
rect 361574 73788 361580 73800
rect 361632 73788 361638 73840
rect 491202 73788 491208 73840
rect 491260 73828 491266 73840
rect 569954 73828 569960 73840
rect 491260 73800 569960 73828
rect 491260 73788 491266 73800
rect 569954 73788 569960 73800
rect 570012 73788 570018 73840
rect 415118 73108 415124 73160
rect 415176 73148 415182 73160
rect 415394 73148 415400 73160
rect 415176 73120 415400 73148
rect 415176 73108 415182 73120
rect 415394 73108 415400 73120
rect 415452 73108 415458 73160
rect 46842 72428 46848 72480
rect 46900 72468 46906 72480
rect 114646 72468 114652 72480
rect 46900 72440 114652 72468
rect 46900 72428 46906 72440
rect 114646 72428 114652 72440
rect 114704 72428 114710 72480
rect 164329 72471 164387 72477
rect 164329 72437 164341 72471
rect 164375 72468 164387 72471
rect 164418 72468 164424 72480
rect 164375 72440 164424 72468
rect 164375 72437 164387 72440
rect 164329 72431 164387 72437
rect 164418 72428 164424 72440
rect 164476 72428 164482 72480
rect 332410 72428 332416 72480
rect 332468 72468 332474 72480
rect 332594 72468 332600 72480
rect 332468 72440 332600 72468
rect 332468 72428 332474 72440
rect 332594 72428 332600 72440
rect 332652 72428 332658 72480
rect 449710 72428 449716 72480
rect 449768 72468 449774 72480
rect 510614 72468 510620 72480
rect 449768 72440 510620 72468
rect 449768 72428 449774 72440
rect 510614 72428 510620 72440
rect 510672 72428 510678 72480
rect 252462 71544 252468 71596
rect 252520 71584 252526 71596
rect 252646 71584 252652 71596
rect 252520 71556 252652 71584
rect 252520 71544 252526 71556
rect 252646 71544 252652 71556
rect 252704 71544 252710 71596
rect 321186 71068 321192 71120
rect 321244 71108 321250 71120
rect 321370 71108 321376 71120
rect 321244 71080 321376 71108
rect 321244 71068 321250 71080
rect 321370 71068 321376 71080
rect 321428 71068 321434 71120
rect 57882 71000 57888 71052
rect 57940 71040 57946 71052
rect 122926 71040 122932 71052
rect 57940 71012 122932 71040
rect 57940 71000 57946 71012
rect 122926 71000 122932 71012
rect 122984 71000 122990 71052
rect 450998 71000 451004 71052
rect 451056 71040 451062 71052
rect 513374 71040 513380 71052
rect 451056 71012 513380 71040
rect 451056 71000 451062 71012
rect 513374 71000 513380 71012
rect 513432 71000 513438 71052
rect 161658 70456 161664 70508
rect 161716 70456 161722 70508
rect 212718 70496 212724 70508
rect 212679 70468 212724 70496
rect 212718 70456 212724 70468
rect 212776 70456 212782 70508
rect 158806 70388 158812 70440
rect 158864 70388 158870 70440
rect 124214 70320 124220 70372
rect 124272 70360 124278 70372
rect 124398 70360 124404 70372
rect 124272 70332 124404 70360
rect 124272 70320 124278 70332
rect 124398 70320 124404 70332
rect 124456 70320 124462 70372
rect 142157 70363 142215 70369
rect 142157 70329 142169 70363
rect 142203 70360 142215 70363
rect 142246 70360 142252 70372
rect 142203 70332 142252 70360
rect 142203 70329 142215 70332
rect 142157 70323 142215 70329
rect 142246 70320 142252 70332
rect 142304 70320 142310 70372
rect 158824 70292 158852 70388
rect 158898 70292 158904 70304
rect 158824 70264 158904 70292
rect 158898 70252 158904 70264
rect 158956 70252 158962 70304
rect 161676 70236 161704 70456
rect 169938 70388 169944 70440
rect 169996 70388 170002 70440
rect 175458 70388 175464 70440
rect 175516 70388 175522 70440
rect 208486 70388 208492 70440
rect 208544 70388 208550 70440
rect 248598 70428 248604 70440
rect 248559 70400 248604 70428
rect 248598 70388 248604 70400
rect 248656 70388 248662 70440
rect 277578 70428 277584 70440
rect 277504 70400 277584 70428
rect 169956 70292 169984 70388
rect 170030 70292 170036 70304
rect 169956 70264 170036 70292
rect 170030 70252 170036 70264
rect 170088 70252 170094 70304
rect 175476 70292 175504 70388
rect 175550 70292 175556 70304
rect 175476 70264 175556 70292
rect 175550 70252 175556 70264
rect 175608 70252 175614 70304
rect 208504 70292 208532 70388
rect 277504 70372 277532 70400
rect 277578 70388 277584 70400
rect 277636 70388 277642 70440
rect 277486 70320 277492 70372
rect 277544 70320 277550 70372
rect 208578 70292 208584 70304
rect 208504 70264 208584 70292
rect 208578 70252 208584 70264
rect 208636 70252 208642 70304
rect 161658 70184 161664 70236
rect 161716 70184 161722 70236
rect 410889 70023 410947 70029
rect 410889 69989 410901 70023
rect 410935 70020 410947 70023
rect 410978 70020 410984 70032
rect 410935 69992 410984 70020
rect 410935 69989 410947 69992
rect 410889 69983 410947 69989
rect 410978 69980 410984 69992
rect 411036 69980 411042 70032
rect 176838 69844 176844 69896
rect 176896 69844 176902 69896
rect 176856 69760 176884 69844
rect 176838 69708 176844 69760
rect 176896 69708 176902 69760
rect 62022 69640 62028 69692
rect 62080 69680 62086 69692
rect 125686 69680 125692 69692
rect 62080 69652 125692 69680
rect 62080 69640 62086 69652
rect 125686 69640 125692 69652
rect 125744 69640 125750 69692
rect 459462 69640 459468 69692
rect 459520 69680 459526 69692
rect 524414 69680 524420 69692
rect 459520 69652 524420 69680
rect 459520 69640 459526 69652
rect 524414 69640 524420 69652
rect 524472 69640 524478 69692
rect 68922 68280 68928 68332
rect 68980 68320 68986 68332
rect 130010 68320 130016 68332
rect 68980 68292 130016 68320
rect 68980 68280 68986 68292
rect 130010 68280 130016 68292
rect 130068 68280 130074 68332
rect 464890 68280 464896 68332
rect 464948 68320 464954 68332
rect 531314 68320 531320 68332
rect 464948 68292 531320 68320
rect 464948 68280 464954 68292
rect 531314 68280 531320 68292
rect 531372 68280 531378 68332
rect 85758 67776 85764 67788
rect 85719 67748 85764 67776
rect 85758 67736 85764 67748
rect 85816 67736 85822 67788
rect 178126 67668 178132 67720
rect 178184 67708 178190 67720
rect 178402 67708 178408 67720
rect 178184 67680 178408 67708
rect 178184 67668 178190 67680
rect 178402 67668 178408 67680
rect 178460 67668 178466 67720
rect 226610 67708 226616 67720
rect 226536 67680 226616 67708
rect 31662 67640 31668 67652
rect 31623 67612 31668 67640
rect 31662 67600 31668 67612
rect 31720 67600 31726 67652
rect 110506 67600 110512 67652
rect 110564 67640 110570 67652
rect 110598 67640 110604 67652
rect 110564 67612 110604 67640
rect 110564 67600 110570 67612
rect 110598 67600 110604 67612
rect 110656 67600 110662 67652
rect 136729 67643 136787 67649
rect 136729 67609 136741 67643
rect 136775 67640 136787 67643
rect 136818 67640 136824 67652
rect 136775 67612 136824 67640
rect 136775 67609 136787 67612
rect 136729 67603 136787 67609
rect 136818 67600 136824 67612
rect 136876 67600 136882 67652
rect 154758 67640 154764 67652
rect 154719 67612 154764 67640
rect 154758 67600 154764 67612
rect 154816 67600 154822 67652
rect 164326 67640 164332 67652
rect 164287 67612 164332 67640
rect 164326 67600 164332 67612
rect 164384 67600 164390 67652
rect 212718 67640 212724 67652
rect 212679 67612 212724 67640
rect 212718 67600 212724 67612
rect 212776 67600 212782 67652
rect 226536 67584 226564 67680
rect 226610 67668 226616 67680
rect 226668 67668 226674 67720
rect 248598 67640 248604 67652
rect 248559 67612 248604 67640
rect 248598 67600 248604 67612
rect 248656 67600 248662 67652
rect 255406 67600 255412 67652
rect 255464 67640 255470 67652
rect 255498 67640 255504 67652
rect 255464 67612 255504 67640
rect 255464 67600 255470 67612
rect 255498 67600 255504 67612
rect 255556 67600 255562 67652
rect 280338 67600 280344 67652
rect 280396 67640 280402 67652
rect 280430 67640 280436 67652
rect 280396 67612 280436 67640
rect 280396 67600 280402 67612
rect 280430 67600 280436 67612
rect 280488 67600 280494 67652
rect 284386 67600 284392 67652
rect 284444 67640 284450 67652
rect 284478 67640 284484 67652
rect 284444 67612 284484 67640
rect 284444 67600 284450 67612
rect 284478 67600 284484 67612
rect 284536 67600 284542 67652
rect 350166 67600 350172 67652
rect 350224 67640 350230 67652
rect 350350 67640 350356 67652
rect 350224 67612 350356 67640
rect 350224 67600 350230 67612
rect 350350 67600 350356 67612
rect 350408 67600 350414 67652
rect 428829 67643 428887 67649
rect 428829 67609 428841 67643
rect 428875 67640 428887 67643
rect 428918 67640 428924 67652
rect 428875 67612 428924 67640
rect 428875 67609 428887 67612
rect 428829 67603 428887 67609
rect 428918 67600 428924 67612
rect 428976 67600 428982 67652
rect 439961 67643 440019 67649
rect 439961 67609 439973 67643
rect 440007 67640 440019 67643
rect 440050 67640 440056 67652
rect 440007 67612 440056 67640
rect 440007 67609 440019 67612
rect 439961 67603 440019 67609
rect 440050 67600 440056 67612
rect 440108 67600 440114 67652
rect 468938 67640 468944 67652
rect 468899 67612 468944 67640
rect 468938 67600 468944 67612
rect 468996 67600 469002 67652
rect 160186 67572 160192 67584
rect 160147 67544 160192 67572
rect 160186 67532 160192 67544
rect 160244 67532 160250 67584
rect 169846 67532 169852 67584
rect 169904 67572 169910 67584
rect 170030 67572 170036 67584
rect 169904 67544 170036 67572
rect 169904 67532 169910 67544
rect 170030 67532 170036 67544
rect 170088 67532 170094 67584
rect 226518 67532 226524 67584
rect 226576 67532 226582 67584
rect 251358 67532 251364 67584
rect 251416 67532 251422 67584
rect 283098 67572 283104 67584
rect 283059 67544 283104 67572
rect 283098 67532 283104 67544
rect 283156 67532 283162 67584
rect 251376 67504 251404 67532
rect 251450 67504 251456 67516
rect 251376 67476 251456 67504
rect 251450 67464 251456 67476
rect 251508 67464 251514 67516
rect 15102 66852 15108 66904
rect 15160 66892 15166 66904
rect 92566 66892 92572 66904
rect 15160 66864 92572 66892
rect 15160 66852 15166 66864
rect 92566 66852 92572 66864
rect 92624 66852 92630 66904
rect 462222 66852 462228 66904
rect 462280 66892 462286 66904
rect 528646 66892 528652 66904
rect 462280 66864 528652 66892
rect 462280 66852 462286 66864
rect 528646 66852 528652 66864
rect 528704 66852 528710 66904
rect 310054 66376 310060 66428
rect 310112 66416 310118 66428
rect 310238 66416 310244 66428
rect 310112 66388 310244 66416
rect 310112 66376 310118 66388
rect 310238 66376 310244 66388
rect 310296 66376 310302 66428
rect 85758 66280 85764 66292
rect 85719 66252 85764 66280
rect 85758 66240 85764 66252
rect 85816 66240 85822 66292
rect 183738 66280 183744 66292
rect 183699 66252 183744 66280
rect 183738 66240 183744 66252
rect 183796 66240 183802 66292
rect 258166 66240 258172 66292
rect 258224 66280 258230 66292
rect 258258 66280 258264 66292
rect 258224 66252 258264 66280
rect 258224 66240 258230 66252
rect 258258 66240 258264 66252
rect 258316 66240 258322 66292
rect 327994 66280 328000 66292
rect 327955 66252 328000 66280
rect 327994 66240 328000 66252
rect 328052 66240 328058 66292
rect 408129 66283 408187 66289
rect 408129 66249 408141 66283
rect 408175 66280 408187 66283
rect 408218 66280 408224 66292
rect 408175 66252 408224 66280
rect 408175 66249 408187 66252
rect 408129 66243 408187 66249
rect 408218 66240 408224 66252
rect 408276 66240 408282 66292
rect 87138 66212 87144 66224
rect 87099 66184 87144 66212
rect 87138 66172 87144 66184
rect 87196 66172 87202 66224
rect 88337 66215 88395 66221
rect 88337 66181 88349 66215
rect 88383 66212 88395 66215
rect 88426 66212 88432 66224
rect 88383 66184 88432 66212
rect 88383 66181 88395 66184
rect 88337 66175 88395 66181
rect 88426 66172 88432 66184
rect 88484 66172 88490 66224
rect 111794 66172 111800 66224
rect 111852 66212 111858 66224
rect 111889 66215 111947 66221
rect 111889 66212 111901 66215
rect 111852 66184 111901 66212
rect 111852 66172 111858 66184
rect 111889 66181 111901 66184
rect 111935 66181 111947 66215
rect 111889 66175 111947 66181
rect 178126 66172 178132 66224
rect 178184 66212 178190 66224
rect 178405 66215 178463 66221
rect 178405 66212 178417 66215
rect 178184 66184 178417 66212
rect 178184 66172 178190 66184
rect 178405 66181 178417 66184
rect 178451 66181 178463 66215
rect 212718 66212 212724 66224
rect 212679 66184 212724 66212
rect 178405 66175 178463 66181
rect 212718 66172 212724 66184
rect 212776 66172 212782 66224
rect 229278 66172 229284 66224
rect 229336 66212 229342 66224
rect 229373 66215 229431 66221
rect 229373 66212 229385 66215
rect 229336 66184 229385 66212
rect 229336 66172 229342 66184
rect 229373 66181 229385 66184
rect 229419 66181 229431 66215
rect 229373 66175 229431 66181
rect 230658 66172 230664 66224
rect 230716 66212 230722 66224
rect 230750 66212 230756 66224
rect 230716 66184 230756 66212
rect 230716 66172 230722 66184
rect 230750 66172 230756 66184
rect 230808 66172 230814 66224
rect 287241 66215 287299 66221
rect 287241 66181 287253 66215
rect 287287 66212 287299 66215
rect 287330 66212 287336 66224
rect 287287 66184 287336 66212
rect 287287 66181 287299 66184
rect 287241 66175 287299 66181
rect 287330 66172 287336 66184
rect 287388 66172 287394 66224
rect 332318 66212 332324 66224
rect 332279 66184 332324 66212
rect 332318 66172 332324 66184
rect 332376 66172 332382 66224
rect 350169 66215 350227 66221
rect 350169 66181 350181 66215
rect 350215 66212 350227 66215
rect 350350 66212 350356 66224
rect 350215 66184 350356 66212
rect 350215 66181 350227 66184
rect 350169 66175 350227 66181
rect 350350 66172 350356 66184
rect 350408 66172 350414 66224
rect 356974 66212 356980 66224
rect 356935 66184 356980 66212
rect 356974 66172 356980 66184
rect 357032 66172 357038 66224
rect 327994 66144 328000 66156
rect 327955 66116 328000 66144
rect 327994 66104 328000 66116
rect 328052 66104 328058 66156
rect 24762 65492 24768 65544
rect 24820 65532 24826 65544
rect 99466 65532 99472 65544
rect 24820 65504 99472 65532
rect 24820 65492 24826 65504
rect 99466 65492 99472 65504
rect 99524 65492 99530 65544
rect 456702 65492 456708 65544
rect 456760 65532 456766 65544
rect 520366 65532 520372 65544
rect 456760 65504 520372 65532
rect 456760 65492 456766 65504
rect 520366 65492 520372 65504
rect 520424 65492 520430 65544
rect 95510 64920 95516 64932
rect 95471 64892 95516 64920
rect 95510 64880 95516 64892
rect 95568 64880 95574 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 79594 64852 79600 64864
rect 3384 64824 79600 64852
rect 3384 64812 3390 64824
rect 79594 64812 79600 64824
rect 79652 64812 79658 64864
rect 321094 64852 321100 64864
rect 321055 64824 321100 64852
rect 321094 64812 321100 64824
rect 321152 64812 321158 64864
rect 519538 64812 519544 64864
rect 519596 64852 519602 64864
rect 579798 64852 579804 64864
rect 519596 64824 579804 64852
rect 519596 64812 519602 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 226518 63928 226524 63980
rect 226576 63968 226582 63980
rect 226613 63971 226671 63977
rect 226613 63968 226625 63971
rect 226576 63940 226625 63968
rect 226576 63928 226582 63940
rect 226613 63937 226625 63940
rect 226659 63937 226671 63971
rect 226613 63931 226671 63937
rect 350169 63903 350227 63909
rect 350169 63869 350181 63903
rect 350215 63900 350227 63903
rect 350350 63900 350356 63912
rect 350215 63872 350356 63900
rect 350215 63869 350227 63872
rect 350169 63863 350227 63869
rect 350350 63860 350356 63872
rect 350408 63860 350414 63912
rect 422018 63560 422024 63572
rect 421979 63532 422024 63560
rect 422018 63520 422024 63532
rect 422076 63520 422082 63572
rect 310054 63452 310060 63504
rect 310112 63492 310118 63504
rect 310241 63495 310299 63501
rect 310241 63492 310253 63495
rect 310112 63464 310253 63492
rect 310112 63452 310118 63464
rect 310241 63461 310253 63464
rect 310287 63461 310299 63495
rect 310241 63455 310299 63461
rect 410978 63452 410984 63504
rect 411036 63492 411042 63504
rect 411070 63492 411076 63504
rect 411036 63464 411076 63492
rect 411036 63452 411042 63464
rect 411070 63452 411076 63464
rect 411128 63452 411134 63504
rect 215386 62772 215392 62824
rect 215444 62812 215450 62824
rect 215570 62812 215576 62824
rect 215444 62784 215576 62812
rect 215444 62772 215450 62784
rect 215570 62772 215576 62784
rect 215628 62772 215634 62824
rect 218146 62772 218152 62824
rect 218204 62812 218210 62824
rect 218330 62812 218336 62824
rect 218204 62784 218336 62812
rect 218204 62772 218210 62784
rect 218330 62772 218336 62784
rect 218388 62772 218394 62824
rect 453942 62772 453948 62824
rect 454000 62812 454006 62824
rect 517514 62812 517520 62824
rect 454000 62784 517520 62812
rect 454000 62772 454006 62784
rect 517514 62772 517520 62784
rect 517572 62772 517578 62824
rect 390002 62092 390008 62144
rect 390060 62132 390066 62144
rect 390094 62132 390100 62144
rect 390060 62104 390100 62132
rect 390060 62092 390066 62104
rect 390094 62092 390100 62104
rect 390152 62092 390158 62144
rect 446950 61344 446956 61396
rect 447008 61384 447014 61396
rect 506474 61384 506480 61396
rect 447008 61356 506480 61384
rect 447008 61344 447014 61356
rect 506474 61344 506480 61356
rect 506532 61344 506538 61396
rect 277486 60868 277492 60920
rect 277544 60908 277550 60920
rect 277544 60880 277624 60908
rect 277544 60868 277550 60880
rect 124398 60840 124404 60852
rect 124359 60812 124404 60840
rect 124398 60800 124404 60812
rect 124456 60800 124462 60852
rect 176838 60840 176844 60852
rect 176764 60812 176844 60840
rect 176764 60784 176792 60812
rect 176838 60800 176844 60812
rect 176896 60800 176902 60852
rect 266630 60840 266636 60852
rect 266556 60812 266636 60840
rect 266556 60784 266584 60812
rect 266630 60800 266636 60812
rect 266688 60800 266694 60852
rect 157518 60772 157524 60784
rect 157352 60744 157524 60772
rect 157352 60716 157380 60744
rect 157518 60732 157524 60744
rect 157576 60732 157582 60784
rect 172790 60732 172796 60784
rect 172848 60772 172854 60784
rect 172848 60744 172928 60772
rect 172848 60732 172854 60744
rect 172900 60716 172928 60744
rect 176746 60732 176752 60784
rect 176804 60732 176810 60784
rect 248690 60732 248696 60784
rect 248748 60732 248754 60784
rect 266538 60732 266544 60784
rect 266596 60732 266602 60784
rect 147858 60664 147864 60716
rect 147916 60664 147922 60716
rect 157334 60664 157340 60716
rect 157392 60664 157398 60716
rect 172882 60664 172888 60716
rect 172940 60664 172946 60716
rect 175366 60664 175372 60716
rect 175424 60704 175430 60716
rect 175550 60704 175556 60716
rect 175424 60676 175556 60704
rect 175424 60664 175430 60676
rect 175550 60664 175556 60676
rect 175608 60664 175614 60716
rect 147876 60636 147904 60664
rect 248708 60648 248736 60732
rect 277596 60716 277624 60880
rect 277578 60664 277584 60716
rect 277636 60664 277642 60716
rect 147950 60636 147956 60648
rect 147876 60608 147956 60636
rect 147950 60596 147956 60608
rect 148008 60596 148014 60648
rect 248690 60596 248696 60648
rect 248748 60596 248754 60648
rect 91002 59984 91008 60036
rect 91060 60024 91066 60036
rect 146386 60024 146392 60036
rect 91060 59996 146392 60024
rect 91060 59984 91066 59996
rect 146386 59984 146392 59996
rect 146444 59984 146450 60036
rect 441522 59984 441528 60036
rect 441580 60024 441586 60036
rect 499574 60024 499580 60036
rect 441580 59996 499580 60024
rect 441580 59984 441586 59996
rect 499574 59984 499580 59996
rect 499632 59984 499638 60036
rect 224862 59848 224868 59900
rect 224920 59888 224926 59900
rect 225046 59888 225052 59900
rect 224920 59860 225052 59888
rect 224920 59848 224926 59860
rect 225046 59848 225052 59860
rect 225104 59848 225110 59900
rect 310238 59208 310244 59220
rect 310199 59180 310244 59208
rect 310238 59168 310244 59180
rect 310296 59168 310302 59220
rect 82722 58624 82728 58676
rect 82780 58664 82786 58676
rect 140866 58664 140872 58676
rect 82780 58636 140872 58664
rect 82780 58624 82786 58636
rect 140866 58624 140872 58636
rect 140924 58624 140930 58676
rect 395890 58624 395896 58676
rect 395948 58664 395954 58676
rect 434714 58664 434720 58676
rect 395948 58636 434720 58664
rect 395948 58624 395954 58636
rect 434714 58624 434720 58636
rect 434772 58624 434778 58676
rect 435910 58624 435916 58676
rect 435968 58664 435974 58676
rect 492674 58664 492680 58676
rect 435968 58636 492680 58664
rect 435968 58624 435974 58636
rect 492674 58624 492680 58636
rect 492732 58624 492738 58676
rect 124306 57944 124312 57996
rect 124364 57984 124370 57996
rect 124401 57987 124459 57993
rect 124401 57984 124413 57987
rect 124364 57956 124413 57984
rect 124364 57944 124370 57956
rect 124401 57953 124413 57956
rect 124447 57953 124459 57987
rect 160186 57984 160192 57996
rect 160147 57956 160192 57984
rect 124401 57947 124459 57953
rect 160186 57944 160192 57956
rect 160244 57944 160250 57996
rect 183738 57944 183744 57996
rect 183796 57944 183802 57996
rect 252462 57944 252468 57996
rect 252520 57984 252526 57996
rect 252646 57984 252652 57996
rect 252520 57956 252652 57984
rect 252520 57944 252526 57956
rect 252646 57944 252652 57956
rect 252704 57944 252710 57996
rect 271966 57944 271972 57996
rect 272024 57984 272030 57996
rect 272058 57984 272064 57996
rect 272024 57956 272064 57984
rect 272024 57944 272030 57956
rect 272058 57944 272064 57956
rect 272116 57944 272122 57996
rect 283098 57984 283104 57996
rect 283059 57956 283104 57984
rect 283098 57944 283104 57956
rect 283156 57944 283162 57996
rect 439866 57944 439872 57996
rect 439924 57984 439930 57996
rect 439958 57984 439964 57996
rect 439924 57956 439964 57984
rect 439924 57944 439930 57956
rect 439958 57944 439964 57956
rect 440016 57944 440022 57996
rect 31662 57916 31668 57928
rect 31623 57888 31668 57916
rect 31662 57876 31668 57888
rect 31720 57876 31726 57928
rect 110690 57916 110696 57928
rect 110651 57888 110696 57916
rect 110690 57876 110696 57888
rect 110748 57876 110754 57928
rect 136821 57919 136879 57925
rect 136821 57885 136833 57919
rect 136867 57916 136879 57919
rect 136910 57916 136916 57928
rect 136867 57888 136916 57916
rect 136867 57885 136879 57888
rect 136821 57879 136879 57885
rect 136910 57876 136916 57888
rect 136968 57876 136974 57928
rect 172882 57916 172888 57928
rect 172843 57888 172888 57916
rect 172882 57876 172888 57888
rect 172940 57876 172946 57928
rect 183756 57860 183784 57944
rect 260834 57876 260840 57928
rect 260892 57916 260898 57928
rect 266449 57919 266507 57925
rect 260892 57888 260937 57916
rect 260892 57876 260898 57888
rect 266449 57885 266461 57919
rect 266495 57916 266507 57919
rect 266538 57916 266544 57928
rect 266495 57888 266544 57916
rect 266495 57885 266507 57888
rect 266449 57879 266507 57885
rect 266538 57876 266544 57888
rect 266596 57876 266602 57928
rect 422294 57876 422300 57928
rect 422352 57916 422358 57928
rect 422386 57916 422392 57928
rect 422352 57888 422392 57916
rect 422352 57876 422358 57888
rect 422386 57876 422392 57888
rect 422444 57876 422450 57928
rect 426250 57916 426256 57928
rect 426211 57888 426256 57916
rect 426250 57876 426256 57888
rect 426308 57876 426314 57928
rect 183738 57808 183744 57860
rect 183796 57808 183802 57860
rect 439866 57848 439872 57860
rect 439827 57820 439872 57848
rect 439866 57808 439872 57820
rect 439924 57808 439930 57860
rect 75822 57196 75828 57248
rect 75880 57236 75886 57248
rect 135254 57236 135260 57248
rect 75880 57208 135260 57236
rect 75880 57196 75886 57208
rect 135254 57196 135260 57208
rect 135312 57196 135318 57248
rect 161382 57196 161388 57248
rect 161440 57236 161446 57248
rect 197446 57236 197452 57248
rect 161440 57208 197452 57236
rect 161440 57196 161446 57208
rect 197446 57196 197452 57208
rect 197504 57196 197510 57248
rect 393130 57196 393136 57248
rect 393188 57236 393194 57248
rect 427817 57239 427875 57245
rect 427817 57236 427829 57239
rect 393188 57208 427829 57236
rect 393188 57196 393194 57208
rect 427817 57205 427829 57208
rect 427863 57205 427875 57239
rect 427817 57199 427875 57205
rect 433242 57196 433248 57248
rect 433300 57236 433306 57248
rect 488534 57236 488540 57248
rect 433300 57208 488540 57236
rect 433300 57196 433306 57208
rect 488534 57196 488540 57208
rect 488592 57196 488598 57248
rect 87138 56624 87144 56636
rect 87099 56596 87144 56624
rect 87138 56584 87144 56596
rect 87196 56584 87202 56636
rect 88334 56624 88340 56636
rect 88295 56596 88340 56624
rect 88334 56584 88340 56596
rect 88392 56584 88398 56636
rect 111886 56624 111892 56636
rect 111847 56596 111892 56624
rect 111886 56584 111892 56596
rect 111944 56584 111950 56636
rect 178402 56584 178408 56636
rect 178460 56624 178466 56636
rect 178460 56596 178505 56624
rect 178460 56584 178466 56596
rect 208486 56584 208492 56636
rect 208544 56624 208550 56636
rect 208670 56624 208676 56636
rect 208544 56596 208676 56624
rect 208544 56584 208550 56596
rect 208670 56584 208676 56596
rect 208728 56584 208734 56636
rect 287238 56624 287244 56636
rect 287199 56596 287244 56624
rect 287238 56584 287244 56596
rect 287296 56584 287302 56636
rect 327994 56624 328000 56636
rect 327955 56596 328000 56624
rect 327994 56584 328000 56596
rect 328052 56584 328058 56636
rect 332321 56627 332379 56633
rect 332321 56593 332333 56627
rect 332367 56624 332379 56627
rect 332410 56624 332416 56636
rect 332367 56596 332416 56624
rect 332367 56593 332379 56596
rect 332321 56587 332379 56593
rect 332410 56584 332416 56596
rect 332468 56584 332474 56636
rect 356977 56627 357035 56633
rect 356977 56593 356989 56627
rect 357023 56624 357035 56627
rect 357066 56624 357072 56636
rect 357023 56596 357072 56624
rect 357023 56593 357035 56596
rect 356977 56587 357035 56593
rect 357066 56584 357072 56596
rect 357124 56584 357130 56636
rect 427817 56627 427875 56633
rect 427817 56593 427829 56627
rect 427863 56624 427875 56627
rect 431954 56624 431960 56636
rect 427863 56596 431960 56624
rect 427863 56593 427875 56596
rect 427817 56587 427875 56593
rect 431954 56584 431960 56596
rect 432012 56584 432018 56636
rect 85758 56556 85764 56568
rect 85719 56528 85764 56556
rect 85758 56516 85764 56528
rect 85816 56516 85822 56568
rect 258166 56488 258172 56500
rect 258127 56460 258172 56488
rect 258166 56448 258172 56460
rect 258224 56448 258230 56500
rect 386138 56012 386144 56024
rect 386099 55984 386144 56012
rect 386138 55972 386144 55984
rect 386196 55972 386202 56024
rect 125502 55836 125508 55888
rect 125560 55876 125566 55888
rect 169846 55876 169852 55888
rect 125560 55848 169852 55876
rect 125560 55836 125566 55848
rect 169846 55836 169852 55848
rect 169904 55836 169910 55888
rect 431862 55836 431868 55888
rect 431920 55876 431926 55888
rect 485774 55876 485780 55888
rect 431920 55848 485780 55876
rect 431920 55836 431926 55848
rect 485774 55836 485780 55848
rect 485832 55836 485838 55888
rect 95326 55224 95332 55276
rect 95384 55264 95390 55276
rect 95418 55264 95424 55276
rect 95384 55236 95424 55264
rect 95384 55224 95390 55236
rect 95418 55224 95424 55236
rect 95476 55224 95482 55276
rect 321097 55267 321155 55273
rect 321097 55233 321109 55267
rect 321143 55264 321155 55267
rect 321186 55264 321192 55276
rect 321143 55236 321192 55264
rect 321143 55233 321155 55236
rect 321097 55227 321155 55233
rect 321186 55224 321192 55236
rect 321244 55224 321250 55276
rect 55122 54476 55128 54528
rect 55180 54516 55186 54528
rect 120074 54516 120080 54528
rect 55180 54488 120080 54516
rect 55180 54476 55186 54488
rect 120074 54476 120080 54488
rect 120132 54476 120138 54528
rect 121362 54476 121368 54528
rect 121420 54516 121426 54528
rect 168466 54516 168472 54528
rect 121420 54488 168472 54516
rect 121420 54476 121426 54488
rect 168466 54476 168472 54488
rect 168524 54476 168530 54528
rect 391198 54476 391204 54528
rect 391256 54516 391262 54528
rect 429194 54516 429200 54528
rect 391256 54488 429200 54516
rect 391256 54476 391262 54488
rect 429194 54476 429200 54488
rect 429252 54476 429258 54528
rect 431218 54476 431224 54528
rect 431276 54516 431282 54528
rect 480254 54516 480260 54528
rect 431276 54488 480260 54516
rect 431276 54476 431282 54488
rect 480254 54476 480260 54488
rect 480312 54476 480318 54528
rect 212721 53839 212779 53845
rect 212721 53805 212733 53839
rect 212767 53836 212779 53839
rect 212810 53836 212816 53848
rect 212767 53808 212816 53836
rect 212767 53805 212779 53808
rect 212721 53799 212779 53805
rect 212810 53796 212816 53808
rect 212868 53796 212874 53848
rect 421926 53796 421932 53848
rect 421984 53836 421990 53848
rect 422018 53836 422024 53848
rect 421984 53808 422024 53836
rect 421984 53796 421990 53808
rect 422018 53796 422024 53808
rect 422076 53796 422082 53848
rect 424870 53116 424876 53168
rect 424928 53156 424934 53168
rect 477586 53156 477592 53168
rect 424928 53128 477592 53156
rect 424928 53116 424934 53128
rect 477586 53116 477592 53128
rect 477644 53116 477650 53168
rect 38470 53048 38476 53100
rect 38528 53088 38534 53100
rect 109034 53088 109040 53100
rect 38528 53060 109040 53088
rect 38528 53048 38534 53060
rect 109034 53048 109040 53060
rect 109092 53048 109098 53100
rect 114462 53048 114468 53100
rect 114520 53088 114526 53100
rect 162854 53088 162860 53100
rect 114520 53060 162860 53088
rect 114520 53048 114526 53060
rect 162854 53048 162860 53060
rect 162912 53048 162918 53100
rect 471790 53048 471796 53100
rect 471848 53088 471854 53100
rect 542354 53088 542360 53100
rect 471848 53060 542360 53088
rect 471848 53048 471854 53060
rect 542354 53048 542360 53060
rect 542412 53048 542418 53100
rect 390186 52436 390192 52488
rect 390244 52476 390250 52488
rect 390278 52476 390284 52488
rect 390244 52448 390284 52476
rect 390244 52436 390250 52448
rect 390278 52436 390284 52448
rect 390336 52436 390342 52488
rect 428829 51867 428887 51873
rect 428829 51833 428841 51867
rect 428875 51864 428887 51867
rect 429010 51864 429016 51876
rect 428875 51836 429016 51864
rect 428875 51833 428887 51836
rect 428829 51827 428887 51833
rect 429010 51824 429016 51836
rect 429068 51824 429074 51876
rect 421926 51756 421932 51808
rect 421984 51796 421990 51808
rect 473354 51796 473360 51808
rect 421984 51768 473360 51796
rect 421984 51756 421990 51768
rect 473354 51756 473360 51768
rect 473412 51756 473418 51808
rect 35802 51688 35808 51740
rect 35860 51728 35866 51740
rect 106458 51728 106464 51740
rect 35860 51700 106464 51728
rect 35860 51688 35866 51700
rect 106458 51688 106464 51700
rect 106516 51688 106522 51740
rect 110322 51688 110328 51740
rect 110380 51728 110386 51740
rect 160186 51728 160192 51740
rect 110380 51700 160192 51728
rect 110380 51688 110386 51700
rect 160186 51688 160192 51700
rect 160244 51688 160250 51740
rect 384850 51688 384856 51740
rect 384908 51728 384914 51740
rect 420914 51728 420920 51740
rect 384908 51700 420920 51728
rect 384908 51688 384914 51700
rect 420914 51688 420920 51700
rect 420972 51688 420978 51740
rect 469122 51688 469128 51740
rect 469180 51728 469186 51740
rect 538214 51728 538220 51740
rect 469180 51700 538220 51728
rect 469180 51688 469186 51700
rect 538214 51688 538220 51700
rect 538272 51688 538278 51740
rect 223666 51144 223672 51196
rect 223724 51144 223730 51196
rect 124306 51116 124312 51128
rect 124267 51088 124312 51116
rect 124306 51076 124312 51088
rect 124364 51076 124370 51128
rect 175550 51116 175556 51128
rect 175384 51088 175556 51116
rect 175384 51060 175412 51088
rect 175550 51076 175556 51088
rect 175608 51076 175614 51128
rect 183738 51076 183744 51128
rect 183796 51076 183802 51128
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 79502 51048 79508 51060
rect 3476 51020 79508 51048
rect 3476 51008 3482 51020
rect 79502 51008 79508 51020
rect 79560 51008 79566 51060
rect 113174 51008 113180 51060
rect 113232 51048 113238 51060
rect 113358 51048 113364 51060
rect 113232 51020 113364 51048
rect 113232 51008 113238 51020
rect 113358 51008 113364 51020
rect 113416 51008 113422 51060
rect 121454 51008 121460 51060
rect 121512 51048 121518 51060
rect 121638 51048 121644 51060
rect 121512 51020 121644 51048
rect 121512 51008 121518 51020
rect 121638 51008 121644 51020
rect 121696 51008 121702 51060
rect 175366 51008 175372 51060
rect 175424 51008 175430 51060
rect 183756 50992 183784 51076
rect 223684 51060 223712 51144
rect 321186 51116 321192 51128
rect 321112 51088 321192 51116
rect 321112 51060 321140 51088
rect 321186 51076 321192 51088
rect 321244 51076 321250 51128
rect 223666 51008 223672 51060
rect 223724 51008 223730 51060
rect 321094 51008 321100 51060
rect 321152 51008 321158 51060
rect 183738 50940 183744 50992
rect 183796 50940 183802 50992
rect 419442 50396 419448 50448
rect 419500 50436 419506 50448
rect 469214 50436 469220 50448
rect 419500 50408 469220 50436
rect 419500 50396 419506 50408
rect 469214 50396 469220 50408
rect 469272 50396 469278 50448
rect 107562 50328 107568 50380
rect 107620 50368 107626 50380
rect 157334 50368 157340 50380
rect 107620 50340 157340 50368
rect 107620 50328 107626 50340
rect 157334 50328 157340 50340
rect 157392 50328 157398 50380
rect 467742 50328 467748 50380
rect 467800 50368 467806 50380
rect 535454 50368 535460 50380
rect 467800 50340 535460 50368
rect 467800 50328 467806 50340
rect 535454 50328 535460 50340
rect 535512 50328 535518 50380
rect 10410 48968 10416 49020
rect 10468 49008 10474 49020
rect 87138 49008 87144 49020
rect 10468 48980 87144 49008
rect 10468 48968 10474 48980
rect 87138 48968 87144 48980
rect 87196 48968 87202 49020
rect 124122 48968 124128 49020
rect 124180 49008 124186 49020
rect 169754 49008 169760 49020
rect 124180 48980 169760 49008
rect 124180 48968 124186 48980
rect 169754 48968 169760 48980
rect 169812 48968 169818 49020
rect 382090 48968 382096 49020
rect 382148 49008 382154 49020
rect 416774 49008 416780 49020
rect 382148 48980 416780 49008
rect 382148 48968 382154 48980
rect 416774 48968 416780 48980
rect 416832 48968 416838 49020
rect 417970 48968 417976 49020
rect 418028 49008 418034 49020
rect 466454 49008 466460 49020
rect 418028 48980 466460 49008
rect 418028 48968 418034 48980
rect 466454 48968 466460 48980
rect 466512 48968 466518 49020
rect 484302 48968 484308 49020
rect 484360 49008 484366 49020
rect 558914 49008 558920 49020
rect 484360 48980 558920 49008
rect 484360 48968 484366 48980
rect 558914 48968 558920 48980
rect 558972 48968 558978 49020
rect 415305 48943 415363 48949
rect 415305 48909 415317 48943
rect 415351 48940 415363 48943
rect 415394 48940 415400 48952
rect 415351 48912 415400 48940
rect 415351 48909 415363 48912
rect 415305 48903 415363 48909
rect 415394 48900 415400 48912
rect 415452 48900 415458 48952
rect 252465 48467 252523 48473
rect 252465 48433 252477 48467
rect 252511 48464 252523 48467
rect 252646 48464 252652 48476
rect 252511 48436 252652 48464
rect 252511 48433 252523 48436
rect 252465 48427 252523 48433
rect 252646 48424 252652 48436
rect 252704 48424 252710 48476
rect 252554 48356 252560 48408
rect 252612 48356 252618 48408
rect 332321 48399 332379 48405
rect 332321 48365 332333 48399
rect 332367 48396 332379 48399
rect 332410 48396 332416 48408
rect 332367 48368 332416 48396
rect 332367 48365 332379 48368
rect 332321 48359 332379 48365
rect 332410 48356 332416 48368
rect 332468 48356 332474 48408
rect 31662 48328 31668 48340
rect 31623 48300 31668 48328
rect 31662 48288 31668 48300
rect 31720 48288 31726 48340
rect 88334 48288 88340 48340
rect 88392 48328 88398 48340
rect 88426 48328 88432 48340
rect 88392 48300 88432 48328
rect 88392 48288 88398 48300
rect 88426 48288 88432 48300
rect 88484 48288 88490 48340
rect 93946 48288 93952 48340
rect 94004 48328 94010 48340
rect 94038 48328 94044 48340
rect 94004 48300 94044 48328
rect 94004 48288 94010 48300
rect 94038 48288 94044 48300
rect 94096 48288 94102 48340
rect 110693 48331 110751 48337
rect 110693 48297 110705 48331
rect 110739 48328 110751 48331
rect 110782 48328 110788 48340
rect 110739 48300 110788 48328
rect 110739 48297 110751 48300
rect 110693 48291 110751 48297
rect 110782 48288 110788 48300
rect 110840 48288 110846 48340
rect 124306 48328 124312 48340
rect 124267 48300 124312 48328
rect 124306 48288 124312 48300
rect 124364 48288 124370 48340
rect 136818 48328 136824 48340
rect 136779 48300 136824 48328
rect 136818 48288 136824 48300
rect 136876 48288 136882 48340
rect 176654 48288 176660 48340
rect 176712 48328 176718 48340
rect 176930 48328 176936 48340
rect 176712 48300 176936 48328
rect 176712 48288 176718 48300
rect 176930 48288 176936 48300
rect 176988 48288 176994 48340
rect 178126 48288 178132 48340
rect 178184 48328 178190 48340
rect 178402 48328 178408 48340
rect 178184 48300 178408 48328
rect 178184 48288 178190 48300
rect 178402 48288 178408 48300
rect 178460 48288 178466 48340
rect 215478 48288 215484 48340
rect 215536 48328 215542 48340
rect 215570 48328 215576 48340
rect 215536 48300 215576 48328
rect 215536 48288 215542 48300
rect 215570 48288 215576 48300
rect 215628 48288 215634 48340
rect 218238 48288 218244 48340
rect 218296 48328 218302 48340
rect 218330 48328 218336 48340
rect 218296 48300 218336 48328
rect 218296 48288 218302 48300
rect 218330 48288 218336 48300
rect 218388 48288 218394 48340
rect 226610 48328 226616 48340
rect 226571 48300 226616 48328
rect 226610 48288 226616 48300
rect 226668 48288 226674 48340
rect 229370 48328 229376 48340
rect 229331 48300 229376 48328
rect 229370 48288 229376 48300
rect 229428 48288 229434 48340
rect 241698 48288 241704 48340
rect 241756 48328 241762 48340
rect 241790 48328 241796 48340
rect 241756 48300 241796 48328
rect 241756 48288 241762 48300
rect 241790 48288 241796 48300
rect 241848 48288 241854 48340
rect 121638 48260 121644 48272
rect 121599 48232 121644 48260
rect 121638 48220 121644 48232
rect 121696 48220 121702 48272
rect 205726 48220 205732 48272
rect 205784 48260 205790 48272
rect 205818 48260 205824 48272
rect 205784 48232 205824 48260
rect 205784 48220 205790 48232
rect 205818 48220 205824 48232
rect 205876 48220 205882 48272
rect 206922 48220 206928 48272
rect 206980 48260 206986 48272
rect 207106 48260 207112 48272
rect 206980 48232 207112 48260
rect 206980 48220 206986 48232
rect 207106 48220 207112 48232
rect 207164 48220 207170 48272
rect 208489 48263 208547 48269
rect 208489 48229 208501 48263
rect 208535 48260 208547 48263
rect 208578 48260 208584 48272
rect 208535 48232 208584 48260
rect 208535 48229 208547 48232
rect 208489 48223 208547 48229
rect 208578 48220 208584 48232
rect 208636 48220 208642 48272
rect 224954 48220 224960 48272
rect 225012 48260 225018 48272
rect 225046 48260 225052 48272
rect 225012 48232 225052 48260
rect 225012 48220 225018 48232
rect 225046 48220 225052 48232
rect 225104 48220 225110 48272
rect 252572 48204 252600 48356
rect 260834 48288 260840 48340
rect 260892 48328 260898 48340
rect 266446 48328 266452 48340
rect 260892 48300 260937 48328
rect 266407 48300 266452 48328
rect 260892 48288 260898 48300
rect 266446 48288 266452 48300
rect 266504 48288 266510 48340
rect 271966 48288 271972 48340
rect 272024 48328 272030 48340
rect 272058 48328 272064 48340
rect 272024 48300 272064 48328
rect 272024 48288 272030 48300
rect 272058 48288 272064 48300
rect 272116 48288 272122 48340
rect 386141 48331 386199 48337
rect 386141 48297 386153 48331
rect 386187 48328 386199 48331
rect 386322 48328 386328 48340
rect 386187 48300 386328 48328
rect 386187 48297 386199 48300
rect 386141 48291 386199 48297
rect 386322 48288 386328 48300
rect 386380 48288 386386 48340
rect 426253 48331 426311 48337
rect 426253 48297 426265 48331
rect 426299 48328 426311 48331
rect 426342 48328 426348 48340
rect 426299 48300 426348 48328
rect 426299 48297 426311 48300
rect 426253 48291 426311 48297
rect 426342 48288 426348 48300
rect 426400 48288 426406 48340
rect 428826 48328 428832 48340
rect 428787 48300 428832 48328
rect 428826 48288 428832 48300
rect 428884 48288 428890 48340
rect 439869 48331 439927 48337
rect 439869 48297 439881 48331
rect 439915 48328 439927 48331
rect 439958 48328 439964 48340
rect 439915 48300 439964 48328
rect 439915 48297 439927 48300
rect 439869 48291 439927 48297
rect 439958 48288 439964 48300
rect 440016 48288 440022 48340
rect 287238 48260 287244 48272
rect 287199 48232 287244 48260
rect 287238 48220 287244 48232
rect 287296 48220 287302 48272
rect 390189 48263 390247 48269
rect 390189 48229 390201 48263
rect 390235 48260 390247 48263
rect 390278 48260 390284 48272
rect 390235 48232 390284 48260
rect 390235 48229 390247 48232
rect 390189 48223 390247 48229
rect 390278 48220 390284 48232
rect 390336 48220 390342 48272
rect 252554 48152 252560 48204
rect 252612 48152 252618 48204
rect 260834 48152 260840 48204
rect 260892 48192 260898 48204
rect 260892 48164 260937 48192
rect 260892 48152 260898 48164
rect 30282 47540 30288 47592
rect 30340 47580 30346 47592
rect 102134 47580 102140 47592
rect 30340 47552 102140 47580
rect 30340 47540 30346 47552
rect 102134 47540 102140 47552
rect 102192 47540 102198 47592
rect 103422 47540 103428 47592
rect 103480 47580 103486 47592
rect 154758 47580 154764 47592
rect 103480 47552 154764 47580
rect 103480 47540 103486 47552
rect 154758 47540 154764 47552
rect 154816 47540 154822 47592
rect 158622 47540 158628 47592
rect 158680 47580 158686 47592
rect 194686 47580 194692 47592
rect 158680 47552 194692 47580
rect 158680 47540 158686 47552
rect 194686 47540 194692 47552
rect 194744 47540 194750 47592
rect 379238 47540 379244 47592
rect 379296 47580 379302 47592
rect 414014 47580 414020 47592
rect 379296 47552 414020 47580
rect 379296 47540 379302 47552
rect 414014 47540 414020 47552
rect 414072 47540 414078 47592
rect 433978 47540 433984 47592
rect 434036 47580 434042 47592
rect 487154 47580 487160 47592
rect 434036 47552 487160 47580
rect 434036 47540 434042 47552
rect 487154 47540 487160 47552
rect 487212 47540 487218 47592
rect 85758 47036 85764 47048
rect 85719 47008 85764 47036
rect 85758 46996 85764 47008
rect 85816 46996 85822 47048
rect 327902 46996 327908 47048
rect 327960 47036 327966 47048
rect 327994 47036 328000 47048
rect 327960 47008 328000 47036
rect 327960 46996 327966 47008
rect 327994 46996 328000 47008
rect 328052 46996 328058 47048
rect 172606 46928 172612 46980
rect 172664 46968 172670 46980
rect 172885 46971 172943 46977
rect 172885 46968 172897 46971
rect 172664 46940 172897 46968
rect 172664 46928 172670 46940
rect 172885 46937 172897 46940
rect 172931 46937 172943 46971
rect 252462 46968 252468 46980
rect 252423 46940 252468 46968
rect 172885 46931 172943 46937
rect 252462 46928 252468 46940
rect 252520 46928 252526 46980
rect 258166 46968 258172 46980
rect 258127 46940 258172 46968
rect 258166 46928 258172 46940
rect 258224 46928 258230 46980
rect 332318 46968 332324 46980
rect 332279 46940 332324 46968
rect 332318 46928 332324 46940
rect 332376 46928 332382 46980
rect 85758 46860 85764 46912
rect 85816 46900 85822 46912
rect 86034 46900 86040 46912
rect 85816 46872 86040 46900
rect 85816 46860 85822 46872
rect 86034 46860 86040 46872
rect 86092 46860 86098 46912
rect 224954 46900 224960 46912
rect 224915 46872 224960 46900
rect 224954 46860 224960 46872
rect 225012 46860 225018 46912
rect 248966 46900 248972 46912
rect 248927 46872 248972 46900
rect 248966 46860 248972 46872
rect 249024 46860 249030 46912
rect 431954 46900 431960 46912
rect 431915 46872 431960 46900
rect 431954 46860 431960 46872
rect 432012 46860 432018 46912
rect 332318 46792 332324 46844
rect 332376 46832 332382 46844
rect 332410 46832 332416 46844
rect 332376 46804 332416 46832
rect 332376 46792 332382 46804
rect 332410 46792 332416 46804
rect 332468 46792 332474 46844
rect 20622 46180 20628 46232
rect 20680 46220 20686 46232
rect 95418 46220 95424 46232
rect 20680 46192 95424 46220
rect 20680 46180 20686 46192
rect 95418 46180 95424 46192
rect 95476 46180 95482 46232
rect 96522 46180 96528 46232
rect 96580 46220 96586 46232
rect 150526 46220 150532 46232
rect 96580 46192 150532 46220
rect 96580 46180 96586 46192
rect 150526 46180 150532 46192
rect 150584 46180 150590 46232
rect 154482 46180 154488 46232
rect 154540 46220 154546 46232
rect 191834 46220 191840 46232
rect 154540 46192 191840 46220
rect 154540 46180 154546 46192
rect 191834 46180 191840 46192
rect 191892 46180 191898 46232
rect 412542 46180 412548 46232
rect 412600 46220 412606 46232
rect 459646 46220 459652 46232
rect 412600 46192 459652 46220
rect 412600 46180 412606 46192
rect 459646 46180 459652 46192
rect 459704 46180 459710 46232
rect 473262 46180 473268 46232
rect 473320 46220 473326 46232
rect 545114 46220 545120 46232
rect 473320 46192 545120 46220
rect 473320 46180 473326 46192
rect 545114 46180 545120 46192
rect 545172 46180 545178 46232
rect 408126 45568 408132 45620
rect 408184 45608 408190 45620
rect 408310 45608 408316 45620
rect 408184 45580 408316 45608
rect 408184 45568 408190 45580
rect 408310 45568 408316 45580
rect 408368 45568 408374 45620
rect 310054 45500 310060 45552
rect 310112 45540 310118 45552
rect 310241 45543 310299 45549
rect 310241 45540 310253 45543
rect 310112 45512 310253 45540
rect 310112 45500 310118 45512
rect 310241 45509 310253 45512
rect 310287 45509 310299 45543
rect 310241 45503 310299 45509
rect 327994 45500 328000 45552
rect 328052 45540 328058 45552
rect 328086 45540 328092 45552
rect 328052 45512 328092 45540
rect 328052 45500 328058 45512
rect 328086 45500 328092 45512
rect 328144 45500 328150 45552
rect 410978 45500 410984 45552
rect 411036 45500 411042 45552
rect 410996 45416 411024 45500
rect 410978 45364 410984 45416
rect 411036 45364 411042 45416
rect 89622 44820 89628 44872
rect 89680 44860 89686 44872
rect 144914 44860 144920 44872
rect 89680 44832 144920 44860
rect 89680 44820 89686 44832
rect 144914 44820 144920 44832
rect 144972 44820 144978 44872
rect 151722 44820 151728 44872
rect 151780 44860 151786 44872
rect 189074 44860 189080 44872
rect 151780 44832 189080 44860
rect 151780 44820 151786 44832
rect 189074 44820 189080 44832
rect 189132 44820 189138 44872
rect 378042 44820 378048 44872
rect 378100 44860 378106 44872
rect 409874 44860 409880 44872
rect 378100 44832 409880 44860
rect 378100 44820 378106 44832
rect 409874 44820 409880 44832
rect 409932 44820 409938 44872
rect 451918 44820 451924 44872
rect 451976 44860 451982 44872
rect 511994 44860 512000 44872
rect 451976 44832 512000 44860
rect 451976 44820 451982 44832
rect 511994 44820 512000 44832
rect 512052 44820 512058 44872
rect 350350 44208 350356 44260
rect 350408 44248 350414 44260
rect 350534 44248 350540 44260
rect 350408 44220 350540 44248
rect 350408 44208 350414 44220
rect 350534 44208 350540 44220
rect 350592 44208 350598 44260
rect 212810 44112 212816 44124
rect 212771 44084 212816 44112
rect 212810 44072 212816 44084
rect 212868 44072 212874 44124
rect 350350 44112 350356 44124
rect 350311 44084 350356 44112
rect 350350 44072 350356 44084
rect 350408 44072 350414 44124
rect 271966 43460 271972 43512
rect 272024 43500 272030 43512
rect 272242 43500 272248 43512
rect 272024 43472 272248 43500
rect 272024 43460 272030 43472
rect 272242 43460 272248 43472
rect 272300 43460 272306 43512
rect 90910 43392 90916 43444
rect 90968 43432 90974 43444
rect 146294 43432 146300 43444
rect 90968 43404 146300 43432
rect 90968 43392 90974 43404
rect 146294 43392 146300 43404
rect 146352 43392 146358 43444
rect 147582 43392 147588 43444
rect 147640 43432 147646 43444
rect 186406 43432 186412 43444
rect 147640 43404 186412 43432
rect 147640 43392 147646 43404
rect 186406 43392 186412 43404
rect 186464 43392 186470 43444
rect 409782 43392 409788 43444
rect 409840 43432 409846 43444
rect 455414 43432 455420 43444
rect 409840 43404 455420 43432
rect 409840 43392 409846 43404
rect 455414 43392 455420 43404
rect 455472 43392 455478 43444
rect 466362 43392 466368 43444
rect 466420 43432 466426 43444
rect 534074 43432 534080 43444
rect 466420 43404 534080 43432
rect 466420 43392 466426 43404
rect 534074 43392 534080 43404
rect 534132 43392 534138 43444
rect 85482 42032 85488 42084
rect 85540 42072 85546 42084
rect 142338 42072 142344 42084
rect 85540 42044 142344 42072
rect 85540 42032 85546 42044
rect 142338 42032 142344 42044
rect 142396 42032 142402 42084
rect 143442 42032 143448 42084
rect 143500 42072 143506 42084
rect 183738 42072 183744 42084
rect 143500 42044 183744 42072
rect 143500 42032 143506 42044
rect 183738 42032 183744 42044
rect 183796 42032 183802 42084
rect 375190 42032 375196 42084
rect 375248 42072 375254 42084
rect 407114 42072 407120 42084
rect 375248 42044 407120 42072
rect 375248 42032 375254 42044
rect 407114 42032 407120 42044
rect 407172 42032 407178 42084
rect 448422 42032 448428 42084
rect 448480 42072 448486 42084
rect 509234 42072 509240 42084
rect 448480 42044 509240 42072
rect 448480 42032 448486 42044
rect 509234 42032 509240 42044
rect 509292 42032 509298 42084
rect 88426 41460 88432 41472
rect 88352 41432 88432 41460
rect 88352 41404 88380 41432
rect 88426 41420 88432 41432
rect 88484 41420 88490 41472
rect 113358 41420 113364 41472
rect 113416 41420 113422 41472
rect 147950 41460 147956 41472
rect 147911 41432 147956 41460
rect 147950 41420 147956 41432
rect 148008 41420 148014 41472
rect 172606 41420 172612 41472
rect 172664 41420 172670 41472
rect 356974 41420 356980 41472
rect 357032 41420 357038 41472
rect 386322 41460 386328 41472
rect 386248 41432 386328 41460
rect 88334 41352 88340 41404
rect 88392 41352 88398 41404
rect 113376 41336 113404 41420
rect 113358 41284 113364 41336
rect 113416 41284 113422 41336
rect 172624 41324 172652 41420
rect 172698 41324 172704 41336
rect 172624 41296 172704 41324
rect 172698 41284 172704 41296
rect 172756 41284 172762 41336
rect 356992 41324 357020 41420
rect 386248 41404 386276 41432
rect 386322 41420 386328 41432
rect 386380 41420 386386 41472
rect 439869 41463 439927 41469
rect 439869 41429 439881 41463
rect 439915 41460 439927 41463
rect 439958 41460 439964 41472
rect 439915 41432 439964 41460
rect 439915 41429 439927 41432
rect 439869 41423 439927 41429
rect 439958 41420 439964 41432
rect 440016 41420 440022 41472
rect 386230 41352 386236 41404
rect 386288 41352 386294 41404
rect 426158 41352 426164 41404
rect 426216 41392 426222 41404
rect 426342 41392 426348 41404
rect 426216 41364 426348 41392
rect 426216 41352 426222 41364
rect 426342 41352 426348 41364
rect 426400 41352 426406 41404
rect 504450 41352 504456 41404
rect 504508 41392 504514 41404
rect 580166 41392 580172 41404
rect 504508 41364 580172 41392
rect 504508 41352 504514 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 357066 41324 357072 41336
rect 356992 41296 357072 41324
rect 357066 41284 357072 41296
rect 357124 41284 357130 41336
rect 81342 40672 81348 40724
rect 81400 40712 81406 40724
rect 139486 40712 139492 40724
rect 81400 40684 139492 40712
rect 81400 40672 81406 40684
rect 139486 40672 139492 40684
rect 139544 40672 139550 40724
rect 140682 40672 140688 40724
rect 140740 40712 140746 40724
rect 182266 40712 182272 40724
rect 140740 40684 182272 40712
rect 140740 40672 140746 40684
rect 182266 40672 182272 40684
rect 182324 40672 182330 40724
rect 310238 40712 310244 40724
rect 310199 40684 310244 40712
rect 310238 40672 310244 40684
rect 310296 40672 310302 40724
rect 406930 40672 406936 40724
rect 406988 40712 406994 40724
rect 451274 40712 451280 40724
rect 406988 40684 451280 40712
rect 406988 40672 406994 40684
rect 451274 40672 451280 40684
rect 451332 40672 451338 40724
rect 287238 39828 287244 39840
rect 287199 39800 287244 39828
rect 287238 39788 287244 39800
rect 287296 39788 287302 39840
rect 64690 39312 64696 39364
rect 64748 39352 64754 39364
rect 128446 39352 128452 39364
rect 64748 39324 128452 39352
rect 64748 39312 64754 39324
rect 128446 39312 128452 39324
rect 128504 39312 128510 39364
rect 136542 39312 136548 39364
rect 136600 39352 136606 39364
rect 179506 39352 179512 39364
rect 136600 39324 179512 39352
rect 136600 39312 136606 39324
rect 179506 39312 179512 39324
rect 179564 39312 179570 39364
rect 402790 39312 402796 39364
rect 402848 39352 402854 39364
rect 444374 39352 444380 39364
rect 402848 39324 444380 39352
rect 402848 39312 402854 39324
rect 444374 39312 444380 39324
rect 444432 39312 444438 39364
rect 445662 39312 445668 39364
rect 445720 39352 445726 39364
rect 505094 39352 505100 39364
rect 445720 39324 505100 39352
rect 445720 39312 445726 39324
rect 505094 39312 505100 39324
rect 505152 39312 505158 39364
rect 178218 38768 178224 38820
rect 178276 38768 178282 38820
rect 219618 38768 219624 38820
rect 219676 38768 219682 38820
rect 153378 38700 153384 38752
rect 153436 38740 153442 38752
rect 153470 38740 153476 38752
rect 153436 38712 153476 38740
rect 153436 38700 153442 38712
rect 153470 38700 153476 38712
rect 153528 38700 153534 38752
rect 176930 38740 176936 38752
rect 176856 38712 176936 38740
rect 176856 38684 176884 38712
rect 176930 38700 176936 38712
rect 176988 38700 176994 38752
rect 178236 38684 178264 38768
rect 219636 38684 219664 38768
rect 223577 38743 223635 38749
rect 223577 38709 223589 38743
rect 223623 38740 223635 38743
rect 223666 38740 223672 38752
rect 223623 38712 223672 38740
rect 223623 38709 223635 38712
rect 223577 38703 223635 38709
rect 223666 38700 223672 38712
rect 223724 38700 223730 38752
rect 260834 38700 260840 38752
rect 260892 38740 260898 38752
rect 260892 38712 260937 38740
rect 260892 38700 260898 38712
rect 110690 38632 110696 38684
rect 110748 38672 110754 38684
rect 110782 38672 110788 38684
rect 110748 38644 110788 38672
rect 110748 38632 110754 38644
rect 110782 38632 110788 38644
rect 110840 38632 110846 38684
rect 121641 38675 121699 38681
rect 121641 38641 121653 38675
rect 121687 38672 121699 38675
rect 121730 38672 121736 38684
rect 121687 38644 121736 38672
rect 121687 38641 121699 38644
rect 121641 38635 121699 38641
rect 121730 38632 121736 38644
rect 121788 38632 121794 38684
rect 147950 38672 147956 38684
rect 147911 38644 147956 38672
rect 147950 38632 147956 38644
rect 148008 38632 148014 38684
rect 176838 38632 176844 38684
rect 176896 38632 176902 38684
rect 178218 38632 178224 38684
rect 178276 38632 178282 38684
rect 208486 38672 208492 38684
rect 208447 38644 208492 38672
rect 208486 38632 208492 38644
rect 208544 38632 208550 38684
rect 211338 38632 211344 38684
rect 211396 38672 211402 38684
rect 211522 38672 211528 38684
rect 211396 38644 211528 38672
rect 211396 38632 211402 38644
rect 211522 38632 211528 38644
rect 211580 38632 211586 38684
rect 219618 38632 219624 38684
rect 219676 38632 219682 38684
rect 230750 38632 230756 38684
rect 230808 38672 230814 38684
rect 230842 38672 230848 38684
rect 230808 38644 230848 38672
rect 230808 38632 230814 38644
rect 230842 38632 230848 38644
rect 230900 38632 230906 38684
rect 252462 38632 252468 38684
rect 252520 38672 252526 38684
rect 252646 38672 252652 38684
rect 252520 38644 252652 38672
rect 252520 38632 252526 38644
rect 252646 38632 252652 38644
rect 252704 38632 252710 38684
rect 266446 38632 266452 38684
rect 266504 38672 266510 38684
rect 266538 38672 266544 38684
rect 266504 38644 266544 38672
rect 266504 38632 266510 38644
rect 266538 38632 266544 38644
rect 266596 38632 266602 38684
rect 390186 38672 390192 38684
rect 390147 38644 390192 38672
rect 390186 38632 390192 38644
rect 390244 38632 390250 38684
rect 439866 38672 439872 38684
rect 439827 38644 439872 38672
rect 439866 38632 439872 38644
rect 439924 38632 439930 38684
rect 31662 38604 31668 38616
rect 31623 38576 31668 38604
rect 31662 38564 31668 38576
rect 31720 38564 31726 38616
rect 158806 38604 158812 38616
rect 158767 38576 158812 38604
rect 158806 38564 158812 38576
rect 158864 38564 158870 38616
rect 207014 38604 207020 38616
rect 206975 38576 207020 38604
rect 207014 38564 207020 38576
rect 207072 38564 207078 38616
rect 226610 38604 226616 38616
rect 226571 38576 226616 38604
rect 226610 38564 226616 38576
rect 226668 38564 226674 38616
rect 229370 38604 229376 38616
rect 229331 38576 229376 38604
rect 229370 38564 229376 38576
rect 229428 38564 229434 38616
rect 258166 38564 258172 38616
rect 258224 38604 258230 38616
rect 258258 38604 258264 38616
rect 258224 38576 258264 38604
rect 258224 38564 258230 38576
rect 258258 38564 258264 38576
rect 258316 38564 258322 38616
rect 271782 38564 271788 38616
rect 271840 38604 271846 38616
rect 271966 38604 271972 38616
rect 271840 38576 271972 38604
rect 271840 38564 271846 38576
rect 271966 38564 271972 38576
rect 272024 38564 272030 38616
rect 284478 38604 284484 38616
rect 284439 38576 284484 38604
rect 284478 38564 284484 38576
rect 284536 38564 284542 38616
rect 386230 38604 386236 38616
rect 386191 38576 386236 38604
rect 386230 38564 386236 38576
rect 386288 38564 386294 38616
rect 422294 38564 422300 38616
rect 422352 38604 422358 38616
rect 422386 38604 422392 38616
rect 422352 38576 422392 38604
rect 422352 38564 422358 38576
rect 422386 38564 422392 38576
rect 422444 38564 422450 38616
rect 50982 37884 50988 37936
rect 51040 37924 51046 37936
rect 117314 37924 117320 37936
rect 51040 37896 117320 37924
rect 51040 37884 51046 37896
rect 117314 37884 117320 37896
rect 117372 37884 117378 37936
rect 119982 37884 119988 37936
rect 120040 37924 120046 37936
rect 166994 37924 167000 37936
rect 120040 37896 167000 37924
rect 120040 37884 120046 37896
rect 166994 37884 167000 37896
rect 167052 37884 167058 37936
rect 168282 37884 168288 37936
rect 168340 37924 168346 37936
rect 201586 37924 201592 37936
rect 168340 37896 201592 37924
rect 168340 37884 168346 37896
rect 201586 37884 201592 37896
rect 201644 37884 201650 37936
rect 372522 37884 372528 37936
rect 372580 37924 372586 37936
rect 402974 37924 402980 37936
rect 372580 37896 402980 37924
rect 372580 37884 372586 37896
rect 402974 37884 402980 37896
rect 403032 37884 403038 37936
rect 442810 37884 442816 37936
rect 442868 37924 442874 37936
rect 502334 37924 502340 37936
rect 442868 37896 502340 37924
rect 442868 37884 442874 37896
rect 502334 37884 502340 37896
rect 502392 37884 502398 37936
rect 223574 37312 223580 37324
rect 223535 37284 223580 37312
rect 223574 37272 223580 37284
rect 223632 37272 223638 37324
rect 224954 37312 224960 37324
rect 224915 37284 224960 37312
rect 224954 37272 224960 37284
rect 225012 37272 225018 37324
rect 248966 37312 248972 37324
rect 248927 37284 248972 37312
rect 248966 37272 248972 37284
rect 249024 37272 249030 37324
rect 431954 37312 431960 37324
rect 431915 37284 431960 37312
rect 431954 37272 431960 37284
rect 432012 37272 432018 37324
rect 321097 37247 321155 37253
rect 321097 37213 321109 37247
rect 321143 37244 321155 37247
rect 321186 37244 321192 37256
rect 321143 37216 321192 37244
rect 321143 37213 321155 37216
rect 321097 37207 321155 37213
rect 321186 37204 321192 37216
rect 321244 37204 321250 37256
rect 357066 37244 357072 37256
rect 357027 37216 357072 37244
rect 357066 37204 357072 37216
rect 357124 37204 357130 37256
rect 369762 36592 369768 36644
rect 369820 36632 369826 36644
rect 400214 36632 400220 36644
rect 369820 36604 400220 36632
rect 369820 36592 369826 36604
rect 400214 36592 400220 36604
rect 400272 36592 400278 36644
rect 10962 36524 10968 36576
rect 11020 36564 11026 36576
rect 88334 36564 88340 36576
rect 11020 36536 88340 36564
rect 11020 36524 11026 36536
rect 88334 36524 88340 36536
rect 88392 36524 88398 36576
rect 117222 36524 117228 36576
rect 117280 36564 117286 36576
rect 164326 36564 164332 36576
rect 117280 36536 164332 36564
rect 117280 36524 117286 36536
rect 164326 36524 164332 36536
rect 164384 36524 164390 36576
rect 165522 36524 165528 36576
rect 165580 36564 165586 36576
rect 200298 36564 200304 36576
rect 165580 36536 200304 36564
rect 165580 36524 165586 36536
rect 200298 36524 200304 36536
rect 200356 36524 200362 36576
rect 399478 36524 399484 36576
rect 399536 36564 399542 36576
rect 438854 36564 438860 36576
rect 399536 36536 438860 36564
rect 399536 36524 399542 36536
rect 438854 36524 438860 36536
rect 438912 36524 438918 36576
rect 439866 36524 439872 36576
rect 439924 36564 439930 36576
rect 498194 36564 498200 36576
rect 439924 36536 498200 36564
rect 439924 36524 439930 36536
rect 498194 36524 498200 36536
rect 498252 36524 498258 36576
rect 415302 35952 415308 35964
rect 415263 35924 415308 35952
rect 415302 35912 415308 35924
rect 415360 35912 415366 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 10318 35884 10324 35896
rect 3476 35856 10324 35884
rect 3476 35844 3482 35856
rect 10318 35844 10324 35856
rect 10376 35844 10382 35896
rect 82630 35164 82636 35216
rect 82688 35204 82694 35216
rect 139394 35204 139400 35216
rect 82688 35176 139400 35204
rect 82688 35164 82694 35176
rect 139394 35164 139400 35176
rect 139452 35164 139458 35216
rect 160002 35164 160008 35216
rect 160060 35204 160066 35216
rect 195974 35204 195980 35216
rect 160060 35176 195980 35204
rect 160060 35164 160066 35176
rect 195974 35164 195980 35176
rect 196032 35164 196038 35216
rect 394602 35164 394608 35216
rect 394660 35204 394666 35216
rect 433334 35204 433340 35216
rect 394660 35176 433340 35204
rect 394660 35164 394666 35176
rect 433334 35164 433340 35176
rect 433392 35164 433398 35216
rect 437382 35164 437388 35216
rect 437440 35204 437446 35216
rect 494054 35204 494060 35216
rect 437440 35176 494060 35204
rect 437440 35164 437446 35176
rect 494054 35164 494060 35176
rect 494112 35164 494118 35216
rect 176746 34660 176752 34672
rect 176707 34632 176752 34660
rect 176746 34620 176752 34632
rect 176804 34620 176810 34672
rect 78582 33736 78588 33788
rect 78640 33776 78646 33788
rect 136910 33776 136916 33788
rect 78640 33748 136916 33776
rect 78640 33736 78646 33748
rect 136910 33736 136916 33748
rect 136968 33736 136974 33788
rect 157242 33736 157248 33788
rect 157300 33776 157306 33788
rect 193306 33776 193312 33788
rect 157300 33748 193312 33776
rect 157300 33736 157306 33748
rect 193306 33736 193312 33748
rect 193364 33736 193370 33788
rect 391842 33736 391848 33788
rect 391900 33776 391906 33788
rect 430574 33776 430580 33788
rect 391900 33748 430580 33776
rect 391900 33736 391906 33748
rect 430574 33736 430580 33748
rect 430632 33736 430638 33788
rect 436002 33736 436008 33788
rect 436060 33776 436066 33788
rect 491294 33776 491300 33788
rect 436060 33748 491300 33776
rect 436060 33736 436066 33748
rect 491294 33736 491300 33748
rect 491352 33736 491358 33788
rect 493962 33736 493968 33788
rect 494020 33776 494026 33788
rect 572714 33776 572720 33788
rect 494020 33748 572720 33776
rect 494020 33736 494026 33748
rect 572714 33736 572720 33748
rect 572772 33736 572778 33788
rect 366910 32444 366916 32496
rect 366968 32484 366974 32496
rect 396074 32484 396080 32496
rect 366968 32456 396080 32484
rect 366968 32444 366974 32456
rect 396074 32444 396080 32456
rect 396132 32444 396138 32496
rect 60642 32376 60648 32428
rect 60700 32416 60706 32428
rect 124214 32416 124220 32428
rect 60700 32388 124220 32416
rect 60700 32376 60706 32388
rect 124214 32376 124220 32388
rect 124272 32376 124278 32428
rect 153102 32376 153108 32428
rect 153160 32416 153166 32428
rect 190546 32416 190552 32428
rect 153160 32388 190552 32416
rect 153160 32376 153166 32388
rect 190546 32376 190552 32388
rect 190604 32376 190610 32428
rect 390186 32376 390192 32428
rect 390244 32416 390250 32428
rect 427814 32416 427820 32428
rect 390244 32388 427820 32416
rect 390244 32376 390250 32388
rect 427814 32376 427820 32388
rect 427872 32376 427878 32428
rect 430482 32376 430488 32428
rect 430540 32416 430546 32428
rect 484394 32416 484400 32428
rect 430540 32388 484400 32416
rect 430540 32376 430546 32388
rect 484394 32376 484400 32388
rect 484452 32376 484458 32428
rect 489730 32376 489736 32428
rect 489788 32416 489794 32428
rect 565814 32416 565820 32428
rect 489788 32388 565820 32416
rect 489788 32376 489794 32388
rect 565814 32376 565820 32388
rect 565872 32376 565878 32428
rect 429010 31872 429016 31884
rect 428971 31844 429016 31872
rect 429010 31832 429016 31844
rect 429068 31832 429074 31884
rect 153470 31804 153476 31816
rect 153431 31776 153476 31804
rect 153470 31764 153476 31776
rect 153528 31764 153534 31816
rect 219618 31764 219624 31816
rect 219676 31764 219682 31816
rect 224954 31764 224960 31816
rect 225012 31764 225018 31816
rect 310238 31804 310244 31816
rect 310164 31776 310244 31804
rect 219636 31668 219664 31764
rect 224972 31680 225000 31764
rect 310164 31748 310192 31776
rect 310238 31764 310244 31776
rect 310296 31764 310302 31816
rect 332410 31804 332416 31816
rect 332336 31776 332416 31804
rect 332336 31748 332364 31776
rect 332410 31764 332416 31776
rect 332468 31764 332474 31816
rect 310146 31696 310152 31748
rect 310204 31696 310210 31748
rect 327905 31739 327963 31745
rect 327905 31705 327917 31739
rect 327951 31736 327963 31739
rect 328086 31736 328092 31748
rect 327951 31708 328092 31736
rect 327951 31705 327963 31708
rect 327905 31699 327963 31705
rect 328086 31696 328092 31708
rect 328144 31696 328150 31748
rect 332318 31696 332324 31748
rect 332376 31696 332382 31748
rect 357066 31736 357072 31748
rect 357027 31708 357072 31736
rect 357066 31696 357072 31708
rect 357124 31696 357130 31748
rect 219710 31668 219716 31680
rect 219636 31640 219716 31668
rect 219710 31628 219716 31640
rect 219768 31628 219774 31680
rect 224954 31628 224960 31680
rect 225012 31628 225018 31680
rect 350350 31668 350356 31680
rect 350311 31640 350356 31668
rect 350350 31628 350356 31640
rect 350408 31628 350414 31680
rect 56410 31016 56416 31068
rect 56468 31056 56474 31068
rect 121730 31056 121736 31068
rect 56468 31028 121736 31056
rect 56468 31016 56474 31028
rect 121730 31016 121736 31028
rect 121788 31016 121794 31068
rect 150342 31016 150348 31068
rect 150400 31056 150406 31068
rect 187786 31056 187792 31068
rect 150400 31028 187792 31056
rect 150400 31016 150406 31028
rect 187786 31016 187792 31028
rect 187844 31016 187850 31068
rect 388990 31016 388996 31068
rect 389048 31056 389054 31068
rect 426434 31056 426440 31068
rect 389048 31028 426440 31056
rect 389048 31016 389054 31028
rect 426434 31016 426440 31028
rect 426492 31016 426498 31068
rect 427078 31016 427084 31068
rect 427136 31056 427142 31068
rect 478874 31056 478880 31068
rect 427136 31028 478880 31056
rect 427136 31016 427142 31028
rect 478874 31016 478880 31028
rect 478932 31016 478938 31068
rect 481542 31016 481548 31068
rect 481600 31056 481606 31068
rect 554866 31056 554872 31068
rect 481600 31028 554872 31056
rect 481600 31016 481606 31028
rect 554866 31016 554872 31028
rect 554924 31016 554930 31068
rect 504358 30268 504364 30320
rect 504416 30308 504422 30320
rect 580166 30308 580172 30320
rect 504416 30280 580172 30308
rect 504416 30268 504422 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 84102 29588 84108 29640
rect 84160 29628 84166 29640
rect 140774 29628 140780 29640
rect 84160 29600 140780 29628
rect 84160 29588 84166 29600
rect 140774 29588 140780 29600
rect 140832 29588 140838 29640
rect 146202 29588 146208 29640
rect 146260 29628 146266 29640
rect 186314 29628 186320 29640
rect 146260 29600 186320 29628
rect 146260 29588 146266 29600
rect 186314 29588 186320 29600
rect 186372 29588 186378 29640
rect 188982 29588 188988 29640
rect 189040 29628 189046 29640
rect 216674 29628 216680 29640
rect 189040 29600 216680 29628
rect 189040 29588 189046 29600
rect 216674 29588 216680 29600
rect 216732 29588 216738 29640
rect 386233 29631 386291 29637
rect 386233 29597 386245 29631
rect 386279 29628 386291 29631
rect 423674 29628 423680 29640
rect 386279 29600 423680 29628
rect 386279 29597 386291 29600
rect 386233 29591 386291 29597
rect 423674 29588 423680 29600
rect 423732 29588 423738 29640
rect 445018 29588 445024 29640
rect 445076 29628 445082 29640
rect 503714 29628 503720 29640
rect 445076 29600 503720 29628
rect 445076 29588 445082 29600
rect 503714 29588 503720 29600
rect 503772 29588 503778 29640
rect 153378 29044 153384 29096
rect 153436 29084 153442 29096
rect 153473 29087 153531 29093
rect 153473 29084 153485 29087
rect 153436 29056 153485 29084
rect 153436 29044 153442 29056
rect 153473 29053 153485 29056
rect 153519 29053 153531 29087
rect 172698 29084 172704 29096
rect 153473 29047 153531 29053
rect 172624 29056 172704 29084
rect 172624 29028 172652 29056
rect 172698 29044 172704 29056
rect 172756 29044 172762 29096
rect 284478 29084 284484 29096
rect 284439 29056 284484 29084
rect 284478 29044 284484 29056
rect 284536 29044 284542 29096
rect 31662 29016 31668 29028
rect 31623 28988 31668 29016
rect 31662 28976 31668 28988
rect 31720 28976 31726 29028
rect 111794 28976 111800 29028
rect 111852 29016 111858 29028
rect 112070 29016 112076 29028
rect 111852 28988 112076 29016
rect 111852 28976 111858 28988
rect 112070 28976 112076 28988
rect 112128 28976 112134 29028
rect 158809 29019 158867 29025
rect 158809 28985 158821 29019
rect 158855 29016 158867 29019
rect 158990 29016 158996 29028
rect 158855 28988 158996 29016
rect 158855 28985 158867 28988
rect 158809 28979 158867 28985
rect 158990 28976 158996 28988
rect 159048 28976 159054 29028
rect 172606 28976 172612 29028
rect 172664 28976 172670 29028
rect 207017 29019 207075 29025
rect 207017 28985 207029 29019
rect 207063 29016 207075 29019
rect 207106 29016 207112 29028
rect 207063 28988 207112 29016
rect 207063 28985 207075 28988
rect 207017 28979 207075 28985
rect 207106 28976 207112 28988
rect 207164 28976 207170 29028
rect 226610 29016 226616 29028
rect 226571 28988 226616 29016
rect 226610 28976 226616 28988
rect 226668 28976 226674 29028
rect 229370 29016 229376 29028
rect 229331 28988 229376 29016
rect 229370 28976 229376 28988
rect 229428 28976 229434 29028
rect 248690 28976 248696 29028
rect 248748 29016 248754 29028
rect 248966 29016 248972 29028
rect 248748 28988 248972 29016
rect 248748 28976 248754 28988
rect 248966 28976 248972 28988
rect 249024 28976 249030 29028
rect 161658 28948 161664 28960
rect 161619 28920 161664 28948
rect 161658 28908 161664 28920
rect 161716 28908 161722 28960
rect 171134 28948 171140 28960
rect 171095 28920 171140 28948
rect 171134 28908 171140 28920
rect 171192 28908 171198 28960
rect 224954 28948 224960 28960
rect 224915 28920 224960 28948
rect 224954 28908 224960 28920
rect 225012 28908 225018 28960
rect 271966 28948 271972 28960
rect 271927 28920 271972 28948
rect 271966 28908 271972 28920
rect 272024 28908 272030 28960
rect 284478 28948 284484 28960
rect 284439 28920 284484 28948
rect 284478 28908 284484 28920
rect 284536 28908 284542 28960
rect 287238 28948 287244 28960
rect 287199 28920 287244 28948
rect 287238 28908 287244 28920
rect 287296 28908 287302 28960
rect 212810 28880 212816 28892
rect 212771 28852 212816 28880
rect 212810 28840 212816 28852
rect 212868 28840 212874 28892
rect 424962 28296 424968 28348
rect 425020 28336 425026 28348
rect 476114 28336 476120 28348
rect 425020 28308 476120 28336
rect 425020 28296 425026 28308
rect 476114 28296 476120 28308
rect 476172 28296 476178 28348
rect 45462 28228 45468 28280
rect 45520 28268 45526 28280
rect 113358 28268 113364 28280
rect 45520 28240 113364 28268
rect 45520 28228 45526 28240
rect 113358 28228 113364 28240
rect 113416 28228 113422 28280
rect 142062 28228 142068 28280
rect 142120 28268 142126 28280
rect 178678 28268 178684 28280
rect 142120 28240 178684 28268
rect 142120 28228 142126 28240
rect 178678 28228 178684 28240
rect 178736 28228 178742 28280
rect 182082 28228 182088 28280
rect 182140 28268 182146 28280
rect 211338 28268 211344 28280
rect 182140 28240 211344 28268
rect 182140 28228 182146 28240
rect 211338 28228 211344 28240
rect 211396 28228 211402 28280
rect 384942 28228 384948 28280
rect 385000 28268 385006 28280
rect 419534 28268 419540 28280
rect 385000 28240 419540 28268
rect 385000 28228 385006 28240
rect 419534 28228 419540 28240
rect 419592 28228 419598 28280
rect 476022 28228 476028 28280
rect 476080 28268 476086 28280
rect 547874 28268 547880 28280
rect 476080 28240 547880 28268
rect 476080 28228 476086 28240
rect 547874 28228 547880 28240
rect 547932 28228 547938 28280
rect 429010 27724 429016 27736
rect 428971 27696 429016 27724
rect 429010 27684 429016 27696
rect 429068 27684 429074 27736
rect 176749 27659 176807 27665
rect 176749 27625 176761 27659
rect 176795 27656 176807 27659
rect 176930 27656 176936 27668
rect 176795 27628 176936 27656
rect 176795 27625 176807 27628
rect 176749 27619 176807 27625
rect 176930 27616 176936 27628
rect 176988 27616 176994 27668
rect 321094 27656 321100 27668
rect 321055 27628 321100 27656
rect 321094 27616 321100 27628
rect 321152 27616 321158 27668
rect 153286 27588 153292 27600
rect 153247 27560 153292 27588
rect 153286 27548 153292 27560
rect 153344 27548 153350 27600
rect 255406 27588 255412 27600
rect 255367 27560 255412 27588
rect 255406 27548 255412 27560
rect 255464 27548 255470 27600
rect 357158 27588 357164 27600
rect 357119 27560 357164 27588
rect 357158 27548 357164 27560
rect 357216 27548 357222 27600
rect 408218 27588 408224 27600
rect 408179 27560 408224 27588
rect 408218 27548 408224 27560
rect 408276 27548 408282 27600
rect 422294 27588 422300 27600
rect 422255 27560 422300 27588
rect 422294 27548 422300 27560
rect 422352 27548 422358 27600
rect 428734 27548 428740 27600
rect 428792 27588 428798 27600
rect 429010 27588 429016 27600
rect 428792 27560 429016 27588
rect 428792 27548 428798 27560
rect 429010 27548 429016 27560
rect 429068 27548 429074 27600
rect 431954 27588 431960 27600
rect 431915 27560 431960 27588
rect 431954 27548 431960 27560
rect 432012 27548 432018 27600
rect 310054 27480 310060 27532
rect 310112 27520 310118 27532
rect 310241 27523 310299 27529
rect 310241 27520 310253 27523
rect 310112 27492 310253 27520
rect 310112 27480 310118 27492
rect 310241 27489 310253 27492
rect 310287 27489 310299 27523
rect 310241 27483 310299 27489
rect 70302 26868 70308 26920
rect 70360 26908 70366 26920
rect 131114 26908 131120 26920
rect 70360 26880 131120 26908
rect 70360 26868 70366 26880
rect 131114 26868 131120 26880
rect 131172 26868 131178 26920
rect 132402 26868 132408 26920
rect 132460 26908 132466 26920
rect 175458 26908 175464 26920
rect 132460 26880 175464 26908
rect 132460 26868 132466 26880
rect 175458 26868 175464 26880
rect 175516 26868 175522 26920
rect 177942 26868 177948 26920
rect 178000 26908 178006 26920
rect 208486 26908 208492 26920
rect 178000 26880 208492 26908
rect 178000 26868 178006 26880
rect 208486 26868 208492 26880
rect 208544 26868 208550 26920
rect 382182 26868 382188 26920
rect 382240 26908 382246 26920
rect 416866 26908 416872 26920
rect 382240 26880 416872 26908
rect 382240 26868 382246 26880
rect 416866 26868 416872 26880
rect 416924 26868 416930 26920
rect 422202 26868 422208 26920
rect 422260 26908 422266 26920
rect 471974 26908 471980 26920
rect 422260 26880 471980 26908
rect 422260 26868 422266 26880
rect 471974 26868 471980 26880
rect 472032 26868 472038 26920
rect 488442 26868 488448 26920
rect 488500 26908 488506 26920
rect 564434 26908 564440 26920
rect 488500 26880 564440 26908
rect 488500 26868 488506 26880
rect 564434 26868 564440 26880
rect 564492 26868 564498 26920
rect 327902 26364 327908 26376
rect 327863 26336 327908 26364
rect 327902 26324 327908 26336
rect 327960 26324 327966 26376
rect 212810 26188 212816 26240
rect 212868 26228 212874 26240
rect 212905 26231 212963 26237
rect 212905 26228 212917 26231
rect 212868 26200 212917 26228
rect 212868 26188 212874 26200
rect 212905 26197 212917 26200
rect 212951 26197 212963 26231
rect 212905 26191 212963 26197
rect 327902 26188 327908 26240
rect 327960 26228 327966 26240
rect 328089 26231 328147 26237
rect 328089 26228 328101 26231
rect 327960 26200 328101 26228
rect 327960 26188 327966 26200
rect 328089 26197 328101 26200
rect 328135 26197 328147 26231
rect 328089 26191 328147 26197
rect 41322 25508 41328 25560
rect 41380 25548 41386 25560
rect 110690 25548 110696 25560
rect 41380 25520 110696 25548
rect 41380 25508 41386 25520
rect 110690 25508 110696 25520
rect 110748 25508 110754 25560
rect 129642 25508 129648 25560
rect 129700 25548 129706 25560
rect 173894 25548 173900 25560
rect 129700 25520 173900 25548
rect 129700 25508 129706 25520
rect 173894 25508 173900 25520
rect 173952 25508 173958 25560
rect 175182 25508 175188 25560
rect 175240 25548 175246 25560
rect 205726 25548 205732 25560
rect 175240 25520 205732 25548
rect 175240 25508 175246 25520
rect 205726 25508 205732 25520
rect 205784 25508 205790 25560
rect 373902 25508 373908 25560
rect 373960 25548 373966 25560
rect 405734 25548 405740 25560
rect 373960 25520 405740 25548
rect 373960 25508 373966 25520
rect 405734 25508 405740 25520
rect 405792 25508 405798 25560
rect 420178 25508 420184 25560
rect 420236 25548 420242 25560
rect 467926 25548 467932 25560
rect 420236 25520 467932 25548
rect 420236 25508 420242 25520
rect 467926 25508 467932 25520
rect 467984 25508 467990 25560
rect 471882 25508 471888 25560
rect 471940 25548 471946 25560
rect 540974 25548 540980 25560
rect 471940 25520 540980 25548
rect 471940 25508 471946 25520
rect 540974 25508 540980 25520
rect 541032 25508 541038 25560
rect 23382 24080 23388 24132
rect 23440 24120 23446 24132
rect 97994 24120 98000 24132
rect 23440 24092 98000 24120
rect 23440 24080 23446 24092
rect 97994 24080 98000 24092
rect 98052 24080 98058 24132
rect 106182 24080 106188 24132
rect 106240 24120 106246 24132
rect 156598 24120 156604 24132
rect 106240 24092 156604 24120
rect 106240 24080 106246 24092
rect 156598 24080 156604 24092
rect 156656 24080 156662 24132
rect 168190 24080 168196 24132
rect 168248 24120 168254 24132
rect 200758 24120 200764 24132
rect 168248 24092 200764 24120
rect 168248 24080 168254 24092
rect 200758 24080 200764 24092
rect 200816 24080 200822 24132
rect 202690 24080 202696 24132
rect 202748 24120 202754 24132
rect 226610 24120 226616 24132
rect 202748 24092 226616 24120
rect 202748 24080 202754 24092
rect 226610 24080 226616 24092
rect 226668 24080 226674 24132
rect 368290 24080 368296 24132
rect 368348 24120 368354 24132
rect 398834 24120 398840 24132
rect 368348 24092 398840 24120
rect 368348 24080 368354 24092
rect 398834 24080 398840 24092
rect 398892 24080 398898 24132
rect 416682 24080 416688 24132
rect 416740 24120 416746 24132
rect 465074 24120 465080 24132
rect 416740 24092 465080 24120
rect 416740 24080 416746 24092
rect 465074 24080 465080 24092
rect 465132 24080 465138 24132
rect 470502 24080 470508 24132
rect 470560 24120 470566 24132
rect 539594 24120 539600 24132
rect 470560 24092 539600 24120
rect 470560 24080 470566 24092
rect 539594 24080 539600 24092
rect 539652 24080 539658 24132
rect 30190 22720 30196 22772
rect 30248 22760 30254 22772
rect 103514 22760 103520 22772
rect 30248 22732 103520 22760
rect 30248 22720 30254 22732
rect 103514 22720 103520 22732
rect 103572 22720 103578 22772
rect 108942 22720 108948 22772
rect 109000 22760 109006 22772
rect 159082 22760 159088 22772
rect 109000 22732 159088 22760
rect 109000 22720 109006 22732
rect 159082 22720 159088 22732
rect 159140 22720 159146 22772
rect 164142 22720 164148 22772
rect 164200 22760 164206 22772
rect 198734 22760 198740 22772
rect 164200 22732 198740 22760
rect 164200 22720 164206 22732
rect 198734 22720 198740 22732
rect 198792 22720 198798 22772
rect 200022 22720 200028 22772
rect 200080 22760 200086 22772
rect 223574 22760 223580 22772
rect 200080 22732 223580 22760
rect 200080 22720 200086 22732
rect 223574 22720 223580 22732
rect 223632 22720 223638 22772
rect 353110 22720 353116 22772
rect 353168 22760 353174 22772
rect 376754 22760 376760 22772
rect 353168 22732 376760 22760
rect 353168 22720 353174 22732
rect 376754 22720 376760 22732
rect 376812 22720 376818 22772
rect 377398 22720 377404 22772
rect 377456 22760 377462 22772
rect 408494 22760 408500 22772
rect 377456 22732 408500 22760
rect 377456 22720 377462 22732
rect 408494 22720 408500 22732
rect 408552 22720 408558 22772
rect 416038 22720 416044 22772
rect 416096 22760 416102 22772
rect 460934 22760 460940 22772
rect 416096 22732 460940 22760
rect 416096 22720 416102 22732
rect 460934 22720 460940 22732
rect 460992 22720 460998 22772
rect 469858 22720 469864 22772
rect 469916 22760 469922 22772
rect 536926 22760 536932 22772
rect 469916 22732 536932 22760
rect 469916 22720 469922 22732
rect 536926 22720 536932 22732
rect 536984 22720 536990 22772
rect 254118 22244 254124 22296
rect 254176 22244 254182 22296
rect 229370 22216 229376 22228
rect 229331 22188 229376 22216
rect 229370 22176 229376 22188
rect 229428 22176 229434 22228
rect 254136 22160 254164 22244
rect 85942 22148 85948 22160
rect 85776 22120 85948 22148
rect 85776 22092 85804 22120
rect 85942 22108 85948 22120
rect 86000 22108 86006 22160
rect 165798 22148 165804 22160
rect 165724 22120 165804 22148
rect 165724 22092 165752 22120
rect 165798 22108 165804 22120
rect 165856 22108 165862 22160
rect 176930 22148 176936 22160
rect 176764 22120 176936 22148
rect 176764 22092 176792 22120
rect 176930 22108 176936 22120
rect 176988 22108 176994 22160
rect 230661 22151 230719 22157
rect 230661 22117 230673 22151
rect 230707 22148 230719 22151
rect 230750 22148 230756 22160
rect 230707 22120 230756 22148
rect 230707 22117 230719 22120
rect 230661 22111 230719 22117
rect 230750 22108 230756 22120
rect 230808 22108 230814 22160
rect 254118 22108 254124 22160
rect 254176 22108 254182 22160
rect 321094 22148 321100 22160
rect 321055 22120 321100 22148
rect 321094 22108 321100 22120
rect 321152 22108 321158 22160
rect 332318 22108 332324 22160
rect 332376 22108 332382 22160
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 79410 22080 79416 22092
rect 3200 22052 79416 22080
rect 3200 22040 3206 22052
rect 79410 22040 79416 22052
rect 79468 22040 79474 22092
rect 85758 22040 85764 22092
rect 85816 22040 85822 22092
rect 111886 22040 111892 22092
rect 111944 22080 111950 22092
rect 112070 22080 112076 22092
rect 111944 22052 112076 22080
rect 111944 22040 111950 22052
rect 112070 22040 112076 22052
rect 112128 22040 112134 22092
rect 165706 22040 165712 22092
rect 165764 22040 165770 22092
rect 176746 22040 176752 22092
rect 176804 22040 176810 22092
rect 332336 22024 332364 22108
rect 332318 21972 332324 22024
rect 332376 21972 332382 22024
rect 328086 21944 328092 21956
rect 328047 21916 328092 21944
rect 328086 21904 328092 21916
rect 328144 21904 328150 21956
rect 128262 21428 128268 21480
rect 128320 21468 128326 21480
rect 172606 21468 172612 21480
rect 128320 21440 172612 21468
rect 128320 21428 128326 21440
rect 172606 21428 172612 21440
rect 172664 21428 172670 21480
rect 86862 21360 86868 21412
rect 86920 21400 86926 21412
rect 143534 21400 143540 21412
rect 86920 21372 143540 21400
rect 86920 21360 86926 21372
rect 143534 21360 143540 21372
rect 143592 21360 143598 21412
rect 171042 21360 171048 21412
rect 171100 21400 171106 21412
rect 204346 21400 204352 21412
rect 171100 21372 204352 21400
rect 171100 21360 171106 21372
rect 204346 21360 204352 21372
rect 204404 21360 204410 21412
rect 206922 21360 206928 21412
rect 206980 21400 206986 21412
rect 229373 21403 229431 21409
rect 229373 21400 229385 21403
rect 206980 21372 229385 21400
rect 206980 21360 206986 21372
rect 229373 21369 229385 21372
rect 229419 21369 229431 21403
rect 229373 21363 229431 21369
rect 348970 21360 348976 21412
rect 349028 21400 349034 21412
rect 369854 21400 369860 21412
rect 349028 21372 369860 21400
rect 349028 21360 349034 21372
rect 369854 21360 369860 21372
rect 369912 21360 369918 21412
rect 371142 21360 371148 21412
rect 371200 21400 371206 21412
rect 401594 21400 401600 21412
rect 371200 21372 401600 21400
rect 371200 21360 371206 21372
rect 401594 21360 401600 21372
rect 401652 21360 401658 21412
rect 410978 21360 410984 21412
rect 411036 21400 411042 21412
rect 458174 21400 458180 21412
rect 411036 21372 458180 21400
rect 411036 21360 411042 21372
rect 458174 21360 458180 21372
rect 458232 21360 458238 21412
rect 463602 21360 463608 21412
rect 463660 21400 463666 21412
rect 529934 21400 529940 21412
rect 463660 21372 529940 21400
rect 463660 21360 463666 21372
rect 529934 21360 529940 21372
rect 529992 21360 529998 21412
rect 19242 19932 19248 19984
rect 19300 19972 19306 19984
rect 94130 19972 94136 19984
rect 19300 19944 94136 19972
rect 19300 19932 19306 19944
rect 94130 19932 94136 19944
rect 94188 19932 94194 19984
rect 102042 19932 102048 19984
rect 102100 19972 102106 19984
rect 154574 19972 154580 19984
rect 102100 19944 154580 19972
rect 102100 19932 102106 19944
rect 154574 19932 154580 19944
rect 154632 19932 154638 19984
rect 159910 19932 159916 19984
rect 159968 19972 159974 19984
rect 194594 19972 194600 19984
rect 159968 19944 194600 19972
rect 159968 19932 159974 19944
rect 194594 19932 194600 19944
rect 194652 19932 194658 19984
rect 195882 19932 195888 19984
rect 195940 19972 195946 19984
rect 222286 19972 222292 19984
rect 195940 19944 222292 19972
rect 195940 19932 195946 19944
rect 222286 19932 222292 19944
rect 222344 19932 222350 19984
rect 370498 19932 370504 19984
rect 370556 19972 370562 19984
rect 387794 19972 387800 19984
rect 370556 19944 387800 19972
rect 370556 19932 370562 19944
rect 387794 19932 387800 19944
rect 387852 19932 387858 19984
rect 409138 19932 409144 19984
rect 409196 19972 409202 19984
rect 454034 19972 454040 19984
rect 409196 19944 454040 19972
rect 409196 19932 409202 19944
rect 454034 19932 454040 19944
rect 454092 19932 454098 19984
rect 458082 19932 458088 19984
rect 458140 19972 458146 19984
rect 523034 19972 523040 19984
rect 458140 19944 523040 19972
rect 458140 19932 458146 19944
rect 523034 19932 523040 19944
rect 523092 19932 523098 19984
rect 224954 19428 224960 19440
rect 224915 19400 224960 19428
rect 224954 19388 224960 19400
rect 225012 19388 225018 19440
rect 161661 19363 161719 19369
rect 161661 19329 161673 19363
rect 161707 19360 161719 19363
rect 161842 19360 161848 19372
rect 161707 19332 161848 19360
rect 161707 19329 161719 19332
rect 161661 19323 161719 19329
rect 161842 19320 161848 19332
rect 161900 19320 161906 19372
rect 171137 19363 171195 19369
rect 171137 19329 171149 19363
rect 171183 19360 171195 19363
rect 171318 19360 171324 19372
rect 171183 19332 171324 19360
rect 171183 19329 171195 19332
rect 171137 19323 171195 19329
rect 171318 19320 171324 19332
rect 171376 19320 171382 19372
rect 207014 19320 207020 19372
rect 207072 19360 207078 19372
rect 207106 19360 207112 19372
rect 207072 19332 207112 19360
rect 207072 19320 207078 19332
rect 207106 19320 207112 19332
rect 207164 19320 207170 19372
rect 230658 19360 230664 19372
rect 230619 19332 230664 19360
rect 230658 19320 230664 19332
rect 230716 19320 230722 19372
rect 271966 19360 271972 19372
rect 271927 19332 271972 19360
rect 271966 19320 271972 19332
rect 272024 19320 272030 19372
rect 284478 19360 284484 19372
rect 284439 19332 284484 19360
rect 284478 19320 284484 19332
rect 284536 19320 284542 19372
rect 287241 19363 287299 19369
rect 287241 19329 287253 19363
rect 287287 19360 287299 19363
rect 287330 19360 287336 19372
rect 287287 19332 287336 19360
rect 287287 19329 287299 19332
rect 287241 19323 287299 19329
rect 287330 19320 287336 19332
rect 287388 19320 287394 19372
rect 31478 19252 31484 19304
rect 31536 19292 31542 19304
rect 31662 19292 31668 19304
rect 31536 19264 31668 19292
rect 31536 19252 31542 19264
rect 31662 19252 31668 19264
rect 31720 19252 31726 19304
rect 112070 19292 112076 19304
rect 112031 19264 112076 19292
rect 112070 19252 112076 19264
rect 112128 19252 112134 19304
rect 212902 19292 212908 19304
rect 212863 19264 212908 19292
rect 212902 19252 212908 19264
rect 212960 19252 212966 19304
rect 224954 19292 224960 19304
rect 224915 19264 224960 19292
rect 224954 19252 224960 19264
rect 225012 19252 225018 19304
rect 248598 19292 248604 19304
rect 248559 19264 248604 19292
rect 248598 19252 248604 19264
rect 248656 19252 248662 19304
rect 260834 19252 260840 19304
rect 260892 19292 260898 19304
rect 260892 19264 260937 19292
rect 260892 19252 260898 19264
rect 193122 18640 193128 18692
rect 193180 18680 193186 18692
rect 214558 18680 214564 18692
rect 193180 18652 214564 18680
rect 193180 18640 193186 18652
rect 214558 18640 214564 18652
rect 214616 18640 214622 18692
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 91094 18612 91100 18624
rect 13688 18584 91100 18612
rect 13688 18572 13694 18584
rect 91094 18572 91100 18584
rect 91152 18572 91158 18624
rect 99190 18572 99196 18624
rect 99248 18612 99254 18624
rect 151814 18612 151820 18624
rect 99248 18584 151820 18612
rect 99248 18572 99254 18584
rect 151814 18572 151820 18584
rect 151872 18572 151878 18624
rect 155862 18572 155868 18624
rect 155920 18612 155926 18624
rect 193214 18612 193220 18624
rect 155920 18584 193220 18612
rect 155920 18572 155926 18584
rect 193214 18572 193220 18584
rect 193272 18572 193278 18624
rect 217962 18572 217968 18624
rect 218020 18612 218026 18624
rect 237466 18612 237472 18624
rect 218020 18584 237472 18612
rect 218020 18572 218026 18584
rect 237466 18572 237472 18584
rect 237524 18572 237530 18624
rect 346210 18572 346216 18624
rect 346268 18612 346274 18624
rect 365714 18612 365720 18624
rect 346268 18584 365720 18612
rect 346268 18572 346274 18584
rect 365714 18572 365720 18584
rect 365772 18572 365778 18624
rect 367002 18572 367008 18624
rect 367060 18612 367066 18624
rect 395433 18615 395491 18621
rect 395433 18612 395445 18615
rect 367060 18584 395445 18612
rect 367060 18572 367066 18584
rect 395433 18581 395445 18584
rect 395479 18581 395491 18615
rect 395433 18575 395491 18581
rect 407022 18572 407028 18624
rect 407080 18612 407086 18624
rect 451366 18612 451372 18624
rect 407080 18584 451372 18612
rect 407080 18572 407086 18584
rect 451366 18572 451372 18584
rect 451424 18572 451430 18624
rect 478782 18572 478788 18624
rect 478840 18612 478846 18624
rect 550634 18612 550640 18624
rect 478840 18584 550640 18612
rect 478840 18572 478846 18584
rect 550634 18572 550640 18584
rect 550692 18572 550698 18624
rect 153289 18003 153347 18009
rect 153289 17969 153301 18003
rect 153335 18000 153347 18003
rect 153378 18000 153384 18012
rect 153335 17972 153384 18000
rect 153335 17969 153347 17972
rect 153289 17963 153347 17969
rect 153378 17960 153384 17972
rect 153436 17960 153442 18012
rect 255406 18000 255412 18012
rect 255367 17972 255412 18000
rect 255406 17960 255412 17972
rect 255464 17960 255470 18012
rect 321094 18000 321100 18012
rect 321055 17972 321100 18000
rect 321094 17960 321100 17972
rect 321152 17960 321158 18012
rect 357161 18003 357219 18009
rect 357161 17969 357173 18003
rect 357207 18000 357219 18003
rect 357250 18000 357256 18012
rect 357207 17972 357256 18000
rect 357207 17969 357219 17972
rect 357161 17963 357219 17969
rect 357250 17960 357256 17972
rect 357308 17960 357314 18012
rect 408221 18003 408279 18009
rect 408221 17969 408233 18003
rect 408267 18000 408279 18003
rect 408402 18000 408408 18012
rect 408267 17972 408408 18000
rect 408267 17969 408279 17972
rect 408221 17963 408279 17969
rect 408402 17960 408408 17972
rect 408460 17960 408466 18012
rect 431954 18000 431960 18012
rect 431915 17972 431960 18000
rect 431954 17960 431960 17972
rect 432012 17960 432018 18012
rect 505738 17892 505744 17944
rect 505796 17932 505802 17944
rect 579798 17932 579804 17944
rect 505796 17904 579804 17932
rect 505796 17892 505802 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 184842 17280 184848 17332
rect 184900 17320 184906 17332
rect 213914 17320 213920 17332
rect 184900 17292 213920 17320
rect 184900 17280 184906 17292
rect 213914 17280 213920 17292
rect 213972 17280 213978 17332
rect 9030 17212 9036 17264
rect 9088 17252 9094 17264
rect 84194 17252 84200 17264
rect 9088 17224 84200 17252
rect 9088 17212 9094 17224
rect 84194 17212 84200 17224
rect 84252 17212 84258 17264
rect 95142 17212 95148 17264
rect 95200 17252 95206 17264
rect 149054 17252 149060 17264
rect 95200 17224 149060 17252
rect 95200 17212 95206 17224
rect 149054 17212 149060 17224
rect 149112 17212 149118 17264
rect 151630 17212 151636 17264
rect 151688 17252 151694 17264
rect 190454 17252 190460 17264
rect 151688 17224 190460 17252
rect 151688 17212 151694 17224
rect 190454 17212 190460 17224
rect 190512 17212 190518 17264
rect 213457 17255 213515 17261
rect 213457 17221 213469 17255
rect 213503 17252 213515 17255
rect 234614 17252 234620 17264
rect 213503 17224 234620 17252
rect 213503 17221 213515 17224
rect 213457 17215 213515 17221
rect 234614 17212 234620 17224
rect 234672 17212 234678 17264
rect 340782 17212 340788 17264
rect 340840 17252 340846 17264
rect 358814 17252 358820 17264
rect 340840 17224 358820 17252
rect 340840 17212 340846 17224
rect 358814 17212 358820 17224
rect 358872 17212 358878 17264
rect 364150 17212 364156 17264
rect 364208 17252 364214 17264
rect 390554 17252 390560 17264
rect 364208 17224 390560 17252
rect 364208 17212 364214 17224
rect 390554 17212 390560 17224
rect 390612 17212 390618 17264
rect 404170 17212 404176 17264
rect 404228 17252 404234 17264
rect 447134 17252 447140 17264
rect 404228 17224 447140 17252
rect 404228 17212 404234 17224
rect 447134 17212 447140 17224
rect 447192 17212 447198 17264
rect 447778 17212 447784 17264
rect 447836 17252 447842 17264
rect 502426 17252 502432 17264
rect 447836 17224 502432 17252
rect 447836 17212 447842 17224
rect 502426 17212 502432 17224
rect 502484 17212 502490 17264
rect 408402 16844 408408 16856
rect 408363 16816 408408 16844
rect 408402 16804 408408 16816
rect 408460 16804 408466 16856
rect 350258 16600 350264 16652
rect 350316 16640 350322 16652
rect 350350 16640 350356 16652
rect 350316 16612 350356 16640
rect 350316 16600 350322 16612
rect 350350 16600 350356 16612
rect 350408 16600 350414 16652
rect 77202 15852 77208 15904
rect 77260 15892 77266 15904
rect 131758 15892 131764 15904
rect 77260 15864 131764 15892
rect 77260 15852 77266 15864
rect 131758 15852 131764 15864
rect 131816 15852 131822 15904
rect 148962 15852 148968 15904
rect 149020 15892 149026 15904
rect 185578 15892 185584 15904
rect 149020 15864 185584 15892
rect 149020 15852 149026 15864
rect 185578 15852 185584 15864
rect 185636 15852 185642 15904
rect 198642 15852 198648 15904
rect 198700 15892 198706 15904
rect 207658 15892 207664 15904
rect 198700 15864 207664 15892
rect 198700 15852 198706 15864
rect 207658 15852 207664 15864
rect 207716 15852 207722 15904
rect 211062 15852 211068 15904
rect 211120 15892 211126 15904
rect 231854 15892 231860 15904
rect 211120 15864 231860 15892
rect 211120 15852 211126 15864
rect 231854 15852 231860 15864
rect 231912 15852 231918 15904
rect 335170 15852 335176 15904
rect 335228 15892 335234 15904
rect 351914 15892 351920 15904
rect 335228 15864 351920 15892
rect 335228 15852 335234 15864
rect 351914 15852 351920 15864
rect 351972 15852 351978 15904
rect 355962 15852 355968 15904
rect 356020 15892 356026 15904
rect 380894 15892 380900 15904
rect 356020 15864 380900 15892
rect 356020 15852 356026 15864
rect 380894 15852 380900 15864
rect 380952 15852 380958 15904
rect 401502 15852 401508 15904
rect 401560 15892 401566 15904
rect 443086 15892 443092 15904
rect 401560 15864 443092 15892
rect 401560 15852 401566 15864
rect 443086 15852 443092 15864
rect 443144 15852 443150 15904
rect 464982 15852 464988 15904
rect 465040 15892 465046 15904
rect 532694 15892 532700 15904
rect 465040 15864 532700 15892
rect 465040 15852 465046 15864
rect 532694 15852 532700 15864
rect 532752 15852 532758 15904
rect 117130 14492 117136 14544
rect 117188 14532 117194 14544
rect 157978 14532 157984 14544
rect 117188 14504 157984 14532
rect 117188 14492 117194 14504
rect 157978 14492 157984 14504
rect 158036 14492 158042 14544
rect 66162 14424 66168 14476
rect 66220 14464 66226 14476
rect 120718 14464 120724 14476
rect 66220 14436 120724 14464
rect 66220 14424 66226 14436
rect 120718 14424 120724 14436
rect 120776 14424 120782 14476
rect 144822 14424 144828 14476
rect 144880 14464 144886 14476
rect 184934 14464 184940 14476
rect 144880 14436 184940 14464
rect 144880 14424 144886 14436
rect 184934 14424 184940 14436
rect 184992 14424 184998 14476
rect 191742 14424 191748 14476
rect 191800 14464 191806 14476
rect 218238 14464 218244 14476
rect 191800 14436 218244 14464
rect 191800 14424 191806 14436
rect 218238 14424 218244 14436
rect 218296 14424 218302 14476
rect 220541 14467 220599 14473
rect 220541 14433 220553 14467
rect 220587 14464 220599 14467
rect 240226 14464 240232 14476
rect 220587 14436 240232 14464
rect 220587 14433 220599 14436
rect 220541 14427 220599 14433
rect 240226 14424 240232 14436
rect 240284 14424 240290 14476
rect 344278 14424 344284 14476
rect 344336 14464 344342 14476
rect 357434 14464 357440 14476
rect 344336 14436 357440 14464
rect 344336 14424 344342 14436
rect 357434 14424 357440 14436
rect 357492 14424 357498 14476
rect 358722 14424 358728 14476
rect 358780 14464 358786 14476
rect 383654 14464 383660 14476
rect 358780 14436 383660 14464
rect 358780 14424 358786 14436
rect 383654 14424 383660 14436
rect 383712 14424 383718 14476
rect 398742 14424 398748 14476
rect 398800 14464 398806 14476
rect 440234 14464 440240 14476
rect 398800 14436 440240 14464
rect 398800 14424 398806 14436
rect 440234 14424 440240 14436
rect 440292 14424 440298 14476
rect 460842 14424 460848 14476
rect 460900 14464 460906 14476
rect 525794 14464 525800 14476
rect 460900 14436 525800 14464
rect 460900 14424 460906 14436
rect 525794 14424 525800 14436
rect 525852 14424 525858 14476
rect 375282 13132 375288 13184
rect 375340 13172 375346 13184
rect 408586 13172 408592 13184
rect 375340 13144 408592 13172
rect 375340 13132 375346 13144
rect 408586 13132 408592 13144
rect 408644 13132 408650 13184
rect 63402 13064 63408 13116
rect 63460 13104 63466 13116
rect 125594 13104 125600 13116
rect 63460 13076 125600 13104
rect 63460 13064 63466 13076
rect 125594 13064 125600 13076
rect 125652 13064 125658 13116
rect 141970 13064 141976 13116
rect 142028 13104 142034 13116
rect 182174 13104 182180 13116
rect 142028 13076 182180 13104
rect 142028 13064 142034 13076
rect 182174 13064 182180 13076
rect 182232 13064 182238 13116
rect 187602 13064 187608 13116
rect 187660 13104 187666 13116
rect 215478 13104 215484 13116
rect 187660 13076 215484 13104
rect 187660 13064 187666 13076
rect 215478 13064 215484 13076
rect 215536 13064 215542 13116
rect 219342 13064 219348 13116
rect 219400 13104 219406 13116
rect 238754 13104 238760 13116
rect 219400 13076 238760 13104
rect 219400 13064 219406 13076
rect 238754 13064 238760 13076
rect 238812 13064 238818 13116
rect 332318 13064 332324 13116
rect 332376 13104 332382 13116
rect 347774 13104 347780 13116
rect 332376 13076 347780 13104
rect 332376 13064 332382 13076
rect 347774 13064 347780 13076
rect 347832 13064 347838 13116
rect 350258 13064 350264 13116
rect 350316 13104 350322 13116
rect 374086 13104 374092 13116
rect 350316 13076 374092 13104
rect 350316 13064 350322 13076
rect 374086 13064 374092 13076
rect 374144 13064 374150 13116
rect 404262 13064 404268 13116
rect 404320 13104 404326 13116
rect 448514 13104 448520 13116
rect 404320 13076 448520 13104
rect 404320 13064 404326 13076
rect 448514 13064 448520 13076
rect 448572 13064 448578 13116
rect 452562 13064 452568 13116
rect 452620 13104 452626 13116
rect 514754 13104 514760 13116
rect 452620 13076 514760 13104
rect 452620 13064 452626 13076
rect 514754 13064 514760 13076
rect 514812 13064 514818 13116
rect 176746 12492 176752 12504
rect 176707 12464 176752 12492
rect 176746 12452 176752 12464
rect 176804 12452 176810 12504
rect 251358 12492 251364 12504
rect 251284 12464 251364 12492
rect 251284 12436 251312 12464
rect 251358 12452 251364 12464
rect 251416 12452 251422 12504
rect 398834 12452 398840 12504
rect 398892 12452 398898 12504
rect 402974 12452 402980 12504
rect 403032 12452 403038 12504
rect 251266 12384 251272 12436
rect 251324 12384 251330 12436
rect 396074 12384 396080 12436
rect 396132 12424 396138 12436
rect 396626 12424 396632 12436
rect 396132 12396 396632 12424
rect 396132 12384 396138 12396
rect 396626 12384 396632 12396
rect 396684 12384 396690 12436
rect 310241 12359 310299 12365
rect 310241 12325 310253 12359
rect 310287 12356 310299 12359
rect 310330 12356 310336 12368
rect 310287 12328 310336 12356
rect 310287 12325 310299 12328
rect 310241 12319 310299 12325
rect 310330 12316 310336 12328
rect 310388 12316 310394 12368
rect 397546 12316 397552 12368
rect 397604 12356 397610 12368
rect 397822 12356 397828 12368
rect 397604 12328 397828 12356
rect 397604 12316 397610 12328
rect 397822 12316 397828 12328
rect 397880 12316 397886 12368
rect 398852 12356 398880 12452
rect 401594 12384 401600 12436
rect 401652 12424 401658 12436
rect 402514 12424 402520 12436
rect 401652 12396 402520 12424
rect 401652 12384 401658 12396
rect 402514 12384 402520 12396
rect 402572 12384 402578 12436
rect 399018 12356 399024 12368
rect 398852 12328 399024 12356
rect 399018 12316 399024 12328
rect 399076 12316 399082 12368
rect 402992 12356 403020 12452
rect 404354 12384 404360 12436
rect 404412 12424 404418 12436
rect 404906 12424 404912 12436
rect 404412 12396 404912 12424
rect 404412 12384 404418 12396
rect 404906 12384 404912 12396
rect 404964 12384 404970 12436
rect 409874 12384 409880 12436
rect 409932 12424 409938 12436
rect 410886 12424 410892 12436
rect 409932 12396 410892 12424
rect 409932 12384 409938 12396
rect 410886 12384 410892 12396
rect 410944 12384 410950 12436
rect 411346 12384 411352 12436
rect 411404 12424 411410 12436
rect 412082 12424 412088 12436
rect 411404 12396 412088 12424
rect 411404 12384 411410 12396
rect 412082 12384 412088 12396
rect 412140 12384 412146 12436
rect 412634 12384 412640 12436
rect 412692 12424 412698 12436
rect 413278 12424 413284 12436
rect 412692 12396 413284 12424
rect 412692 12384 412698 12396
rect 413278 12384 413284 12396
rect 413336 12384 413342 12436
rect 414014 12384 414020 12436
rect 414072 12424 414078 12436
rect 414474 12424 414480 12436
rect 414072 12396 414480 12424
rect 414072 12384 414078 12396
rect 414474 12384 414480 12396
rect 414532 12384 414538 12436
rect 419534 12384 419540 12436
rect 419592 12424 419598 12436
rect 420362 12424 420368 12436
rect 419592 12396 420368 12424
rect 419592 12384 419598 12396
rect 420362 12384 420368 12396
rect 420420 12384 420426 12436
rect 420914 12384 420920 12436
rect 420972 12424 420978 12436
rect 421558 12424 421564 12436
rect 420972 12396 421564 12424
rect 420972 12384 420978 12396
rect 421558 12384 421564 12396
rect 421616 12384 421622 12436
rect 426434 12384 426440 12436
rect 426492 12424 426498 12436
rect 427538 12424 427544 12436
rect 426492 12396 427544 12424
rect 426492 12384 426498 12396
rect 427538 12384 427544 12396
rect 427596 12384 427602 12436
rect 427814 12384 427820 12436
rect 427872 12424 427878 12436
rect 428734 12424 428740 12436
rect 427872 12396 428740 12424
rect 427872 12384 427878 12396
rect 428734 12384 428740 12396
rect 428792 12384 428798 12436
rect 429194 12384 429200 12436
rect 429252 12424 429258 12436
rect 429930 12424 429936 12436
rect 429252 12396 429936 12424
rect 429252 12384 429258 12396
rect 429930 12384 429936 12396
rect 429988 12384 429994 12436
rect 430574 12384 430580 12436
rect 430632 12424 430638 12436
rect 431126 12424 431132 12436
rect 430632 12396 431132 12424
rect 430632 12384 430638 12396
rect 431126 12384 431132 12396
rect 431184 12384 431190 12436
rect 434714 12384 434720 12436
rect 434772 12424 434778 12436
rect 435818 12424 435824 12436
rect 434772 12396 435824 12424
rect 434772 12384 434778 12396
rect 435818 12384 435824 12396
rect 435876 12384 435882 12436
rect 403710 12356 403716 12368
rect 402992 12328 403716 12356
rect 403710 12316 403716 12328
rect 403768 12316 403774 12368
rect 112070 11880 112076 11892
rect 112031 11852 112076 11880
rect 112070 11840 112076 11852
rect 112128 11840 112134 11892
rect 59262 11704 59268 11756
rect 59320 11744 59326 11756
rect 122834 11744 122840 11756
rect 59320 11716 122840 11744
rect 59320 11704 59326 11716
rect 122834 11704 122840 11716
rect 122892 11704 122898 11756
rect 137922 11704 137928 11756
rect 137980 11744 137986 11756
rect 179414 11744 179420 11756
rect 137980 11716 179420 11744
rect 137980 11704 137986 11716
rect 179414 11704 179420 11716
rect 179472 11704 179478 11756
rect 183738 11704 183744 11756
rect 183796 11744 183802 11756
rect 212902 11744 212908 11756
rect 183796 11716 212908 11744
rect 183796 11704 183802 11716
rect 212902 11704 212908 11716
rect 212960 11704 212966 11756
rect 215846 11704 215852 11756
rect 215904 11744 215910 11756
rect 236086 11744 236092 11756
rect 215904 11716 236092 11744
rect 215904 11704 215910 11716
rect 236086 11704 236092 11716
rect 236144 11704 236150 11756
rect 331030 11704 331036 11756
rect 331088 11744 331094 11756
rect 345014 11744 345020 11756
rect 331088 11716 345020 11744
rect 331088 11704 331094 11716
rect 345014 11704 345020 11716
rect 345072 11704 345078 11756
rect 347038 11704 347044 11756
rect 347096 11744 347102 11756
rect 362954 11744 362960 11756
rect 347096 11716 362960 11744
rect 347096 11704 347102 11716
rect 362954 11704 362960 11716
rect 363012 11704 363018 11756
rect 365622 11704 365628 11756
rect 365680 11744 365686 11756
rect 394234 11744 394240 11756
rect 365680 11716 394240 11744
rect 365680 11704 365686 11716
rect 394234 11704 394240 11716
rect 394292 11704 394298 11756
rect 395982 11704 395988 11756
rect 396040 11744 396046 11756
rect 437014 11744 437020 11756
rect 396040 11716 437020 11744
rect 396040 11704 396046 11716
rect 437014 11704 437020 11716
rect 437072 11704 437078 11756
rect 449802 11704 449808 11756
rect 449860 11744 449866 11756
rect 512086 11744 512092 11756
rect 449860 11716 512092 11744
rect 449860 11704 449866 11716
rect 512086 11704 512092 11716
rect 512144 11704 512150 11756
rect 48222 10276 48228 10328
rect 48280 10316 48286 10328
rect 115934 10316 115940 10328
rect 48280 10288 115940 10316
rect 48280 10276 48286 10288
rect 115934 10276 115940 10288
rect 115992 10276 115998 10328
rect 133782 10276 133788 10328
rect 133840 10316 133846 10328
rect 176749 10319 176807 10325
rect 176749 10316 176761 10319
rect 133840 10288 176761 10316
rect 133840 10276 133846 10288
rect 176749 10285 176761 10288
rect 176795 10285 176807 10319
rect 176749 10279 176807 10285
rect 180150 10276 180156 10328
rect 180208 10316 180214 10328
rect 211154 10316 211160 10328
rect 180208 10288 211160 10316
rect 180208 10276 180214 10288
rect 211154 10276 211160 10288
rect 211212 10276 211218 10328
rect 212258 10276 212264 10328
rect 212316 10316 212322 10328
rect 233326 10316 233332 10328
rect 212316 10288 233332 10316
rect 212316 10276 212322 10288
rect 233326 10276 233332 10288
rect 233384 10276 233390 10328
rect 233694 10276 233700 10328
rect 233752 10316 233758 10328
rect 248601 10319 248659 10325
rect 248601 10316 248613 10319
rect 233752 10288 248613 10316
rect 233752 10276 233758 10288
rect 248601 10285 248613 10288
rect 248647 10285 248659 10319
rect 248601 10279 248659 10285
rect 329742 10276 329748 10328
rect 329800 10316 329806 10328
rect 343634 10316 343640 10328
rect 329800 10288 343640 10316
rect 329800 10276 329806 10288
rect 343634 10276 343640 10288
rect 343692 10276 343698 10328
rect 362862 10276 362868 10328
rect 362920 10316 362926 10328
rect 390646 10316 390652 10328
rect 362920 10288 390652 10316
rect 362920 10276 362926 10288
rect 390646 10276 390652 10288
rect 390704 10276 390710 10328
rect 393222 10276 393228 10328
rect 393280 10316 393286 10328
rect 433518 10316 433524 10328
rect 393280 10288 433524 10316
rect 393280 10276 393286 10288
rect 433518 10276 433524 10288
rect 433576 10276 433582 10328
rect 447042 10276 447048 10328
rect 447100 10316 447106 10328
rect 507854 10316 507860 10328
rect 447100 10288 507860 10316
rect 447100 10276 447106 10288
rect 507854 10276 507860 10288
rect 507912 10276 507918 10328
rect 328086 9732 328092 9784
rect 328144 9732 328150 9784
rect 213454 9704 213460 9716
rect 213415 9676 213460 9704
rect 213454 9664 213460 9676
rect 213512 9664 213518 9716
rect 220538 9704 220544 9716
rect 220499 9676 220544 9704
rect 220538 9664 220544 9676
rect 220596 9664 220602 9716
rect 224957 9707 225015 9713
rect 224957 9673 224969 9707
rect 225003 9704 225015 9707
rect 225046 9704 225052 9716
rect 225003 9676 225052 9704
rect 225003 9673 225015 9676
rect 224957 9667 225015 9673
rect 225046 9664 225052 9676
rect 225104 9664 225110 9716
rect 260837 9707 260895 9713
rect 260837 9673 260849 9707
rect 260883 9704 260895 9707
rect 261018 9704 261024 9716
rect 260883 9676 261024 9704
rect 260883 9673 260895 9676
rect 260837 9667 260895 9673
rect 261018 9664 261024 9676
rect 261076 9664 261082 9716
rect 328104 9648 328132 9732
rect 395430 9704 395436 9716
rect 395391 9676 395436 9704
rect 395430 9664 395436 9676
rect 395488 9664 395494 9716
rect 408402 9704 408408 9716
rect 408363 9676 408408 9704
rect 408402 9664 408408 9676
rect 408460 9664 408466 9716
rect 422297 9707 422355 9713
rect 422297 9673 422309 9707
rect 422343 9704 422355 9707
rect 422754 9704 422760 9716
rect 422343 9676 422760 9704
rect 422343 9673 422355 9676
rect 422297 9667 422355 9673
rect 422754 9664 422760 9676
rect 422812 9664 422818 9716
rect 31481 9639 31539 9645
rect 31481 9605 31493 9639
rect 31527 9636 31539 9639
rect 31662 9636 31668 9648
rect 31527 9608 31668 9636
rect 31527 9605 31539 9608
rect 31481 9599 31539 9605
rect 31662 9596 31668 9608
rect 31720 9596 31726 9648
rect 85758 9636 85764 9648
rect 85719 9608 85764 9636
rect 85758 9596 85764 9608
rect 85816 9596 85822 9648
rect 151541 9639 151599 9645
rect 151541 9605 151553 9639
rect 151587 9636 151599 9639
rect 151630 9636 151636 9648
rect 151587 9608 151636 9636
rect 151587 9605 151599 9608
rect 151541 9599 151599 9605
rect 151630 9596 151636 9608
rect 151688 9596 151694 9648
rect 271966 9636 271972 9648
rect 271927 9608 271972 9636
rect 271966 9596 271972 9608
rect 272024 9596 272030 9648
rect 283650 9596 283656 9648
rect 283708 9636 283714 9648
rect 284478 9636 284484 9648
rect 283708 9608 284484 9636
rect 283708 9596 283714 9608
rect 284478 9596 284484 9608
rect 284536 9596 284542 9648
rect 328086 9596 328092 9648
rect 328144 9596 328150 9648
rect 357434 9596 357440 9648
rect 357492 9636 357498 9648
rect 358541 9639 358599 9645
rect 358541 9636 358553 9639
rect 357492 9608 358553 9636
rect 357492 9596 357498 9608
rect 358541 9605 358553 9608
rect 358587 9605 358599 9639
rect 358541 9599 358599 9605
rect 358814 9596 358820 9648
rect 358872 9636 358878 9648
rect 359737 9639 359795 9645
rect 359737 9636 359749 9639
rect 358872 9608 359749 9636
rect 358872 9596 358878 9608
rect 359737 9605 359749 9608
rect 359783 9605 359795 9639
rect 359737 9599 359795 9605
rect 397822 9596 397828 9648
rect 397880 9596 397886 9648
rect 399018 9596 399024 9648
rect 399076 9596 399082 9648
rect 403710 9596 403716 9648
rect 403768 9596 403774 9648
rect 406102 9636 406108 9648
rect 406063 9608 406108 9636
rect 406102 9596 406108 9608
rect 406160 9596 406166 9648
rect 407298 9636 407304 9648
rect 407259 9608 407304 9636
rect 407298 9596 407304 9608
rect 407356 9596 407362 9648
rect 414474 9636 414480 9648
rect 414435 9608 414480 9636
rect 414474 9596 414480 9608
rect 414532 9596 414538 9648
rect 428918 9636 428924 9648
rect 428879 9608 428924 9636
rect 428918 9596 428924 9608
rect 428976 9596 428982 9648
rect 431126 9636 431132 9648
rect 431087 9608 431132 9636
rect 431126 9596 431132 9608
rect 431184 9596 431190 9648
rect 432322 9636 432328 9648
rect 432283 9608 432328 9636
rect 432322 9596 432328 9608
rect 432380 9596 432386 9648
rect 321094 9568 321100 9580
rect 321055 9540 321100 9568
rect 321094 9528 321100 9540
rect 321152 9528 321158 9580
rect 397840 9512 397868 9596
rect 399036 9512 399064 9596
rect 403728 9512 403756 9596
rect 397822 9460 397828 9512
rect 397880 9460 397886 9512
rect 399018 9460 399024 9512
rect 399076 9460 399082 9512
rect 403710 9460 403716 9512
rect 403768 9460 403774 9512
rect 130194 8984 130200 9036
rect 130252 9024 130258 9036
rect 175274 9024 175280 9036
rect 130252 8996 175280 9024
rect 130252 8984 130258 8996
rect 175274 8984 175280 8996
rect 175332 8984 175338 9036
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 77938 8956 77944 8968
rect 2924 8928 77944 8956
rect 2924 8916 2930 8928
rect 77938 8916 77944 8928
rect 77996 8916 78002 8968
rect 79042 8916 79048 8968
rect 79100 8956 79106 8968
rect 138014 8956 138020 8968
rect 79100 8928 138020 8956
rect 79100 8916 79106 8928
rect 138014 8916 138020 8928
rect 138072 8916 138078 8968
rect 176562 8916 176568 8968
rect 176620 8956 176626 8968
rect 208394 8956 208400 8968
rect 176620 8928 208400 8956
rect 176620 8916 176626 8928
rect 208394 8916 208400 8928
rect 208452 8916 208458 8968
rect 208670 8916 208676 8968
rect 208728 8956 208734 8968
rect 230750 8956 230756 8968
rect 208728 8928 230756 8956
rect 208728 8916 208734 8928
rect 230750 8916 230756 8928
rect 230808 8916 230814 8968
rect 237190 8916 237196 8968
rect 237248 8956 237254 8968
rect 251266 8956 251272 8968
rect 237248 8928 251272 8956
rect 237248 8916 237254 8928
rect 251266 8916 251272 8928
rect 251324 8916 251330 8968
rect 338758 8916 338764 8968
rect 338816 8956 338822 8968
rect 356146 8956 356152 8968
rect 338816 8928 356152 8956
rect 338816 8916 338822 8928
rect 356146 8916 356152 8928
rect 356204 8916 356210 8968
rect 360010 8916 360016 8968
rect 360068 8956 360074 8968
rect 387058 8956 387064 8968
rect 360068 8928 387064 8956
rect 360068 8916 360074 8928
rect 387058 8916 387064 8928
rect 387116 8916 387122 8968
rect 389082 8916 389088 8968
rect 389140 8956 389146 8968
rect 426342 8956 426348 8968
rect 389140 8928 426348 8956
rect 389140 8916 389146 8928
rect 426342 8916 426348 8928
rect 426400 8916 426406 8968
rect 440142 8916 440148 8968
rect 440200 8956 440206 8968
rect 497734 8956 497740 8968
rect 440200 8928 497740 8956
rect 440200 8916 440206 8928
rect 497734 8916 497740 8928
rect 497792 8916 497798 8968
rect 499482 8916 499488 8968
rect 499540 8956 499546 8968
rect 580994 8956 581000 8968
rect 499540 8928 581000 8956
rect 499540 8916 499546 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 337378 8508 337384 8560
rect 337436 8548 337442 8560
rect 340690 8548 340696 8560
rect 337436 8520 340696 8548
rect 337436 8508 337442 8520
rect 340690 8508 340696 8520
rect 340748 8508 340754 8560
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 79318 8276 79324 8288
rect 4120 8248 79324 8276
rect 4120 8236 4126 8248
rect 79318 8236 79324 8248
rect 79376 8236 79382 8288
rect 169386 7624 169392 7676
rect 169444 7664 169450 7676
rect 202874 7664 202880 7676
rect 169444 7636 202880 7664
rect 169444 7624 169450 7636
rect 202874 7624 202880 7636
rect 202932 7624 202938 7676
rect 390554 7624 390560 7676
rect 390612 7664 390618 7676
rect 391842 7664 391848 7676
rect 390612 7636 391848 7664
rect 390612 7624 390618 7636
rect 391842 7624 391848 7636
rect 391900 7624 391906 7676
rect 408494 7624 408500 7676
rect 408552 7664 408558 7676
rect 409690 7664 409696 7676
rect 408552 7636 409696 7664
rect 408552 7624 408558 7636
rect 409690 7624 409696 7636
rect 409748 7624 409754 7676
rect 71866 7556 71872 7608
rect 71924 7596 71930 7608
rect 132494 7596 132500 7608
rect 71924 7568 132500 7596
rect 71924 7556 71930 7568
rect 132494 7556 132500 7568
rect 132552 7556 132558 7608
rect 134886 7556 134892 7608
rect 134944 7596 134950 7608
rect 178218 7596 178224 7608
rect 134944 7568 178224 7596
rect 134944 7556 134950 7568
rect 178218 7556 178224 7568
rect 178276 7556 178282 7608
rect 205082 7556 205088 7608
rect 205140 7596 205146 7608
rect 229094 7596 229100 7608
rect 205140 7568 229100 7596
rect 205140 7556 205146 7568
rect 229094 7556 229100 7568
rect 229152 7556 229158 7608
rect 230106 7556 230112 7608
rect 230164 7596 230170 7608
rect 247126 7596 247132 7608
rect 230164 7568 247132 7596
rect 230164 7556 230170 7568
rect 247126 7556 247132 7568
rect 247184 7556 247190 7608
rect 324130 7556 324136 7608
rect 324188 7596 324194 7608
rect 337102 7596 337108 7608
rect 324188 7568 337108 7596
rect 324188 7556 324194 7568
rect 337102 7556 337108 7568
rect 337160 7556 337166 7608
rect 344922 7556 344928 7608
rect 344980 7596 344986 7608
rect 365806 7596 365812 7608
rect 344980 7568 365812 7596
rect 344980 7556 344986 7568
rect 365806 7556 365812 7568
rect 365864 7556 365870 7608
rect 380802 7556 380808 7608
rect 380860 7596 380866 7608
rect 415670 7596 415676 7608
rect 380860 7568 415676 7596
rect 380860 7556 380866 7568
rect 415670 7556 415676 7568
rect 415728 7556 415734 7608
rect 416774 7556 416780 7608
rect 416832 7596 416838 7608
rect 417970 7596 417976 7608
rect 416832 7568 417976 7596
rect 416832 7556 416838 7568
rect 417970 7556 417976 7568
rect 418028 7556 418034 7608
rect 438118 7556 438124 7608
rect 438176 7596 438182 7608
rect 494146 7596 494152 7608
rect 438176 7568 494152 7596
rect 438176 7556 438182 7568
rect 494146 7556 494152 7568
rect 494204 7556 494210 7608
rect 496722 7556 496728 7608
rect 496780 7596 496786 7608
rect 577406 7596 577412 7608
rect 496780 7568 577412 7596
rect 496780 7556 496786 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 132586 6196 132592 6248
rect 132644 6236 132650 6248
rect 142798 6236 142804 6248
rect 132644 6208 142804 6236
rect 132644 6196 132650 6208
rect 142798 6196 142804 6208
rect 142856 6196 142862 6248
rect 194410 6196 194416 6248
rect 194468 6236 194474 6248
rect 220814 6236 220820 6248
rect 194468 6208 220820 6236
rect 194468 6196 194474 6208
rect 220814 6196 220820 6208
rect 220872 6196 220878 6248
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 75178 6168 75184 6180
rect 7708 6140 75184 6168
rect 7708 6128 7714 6140
rect 75178 6128 75184 6140
rect 75236 6128 75242 6180
rect 112346 6128 112352 6180
rect 112404 6168 112410 6180
rect 161842 6168 161848 6180
rect 112404 6140 161848 6168
rect 112404 6128 112410 6140
rect 161842 6128 161848 6140
rect 161900 6128 161906 6180
rect 162302 6128 162308 6180
rect 162360 6168 162366 6180
rect 197354 6168 197360 6180
rect 162360 6140 197360 6168
rect 162360 6128 162366 6140
rect 197354 6128 197360 6140
rect 197412 6128 197418 6180
rect 222930 6128 222936 6180
rect 222988 6168 222994 6180
rect 239398 6168 239404 6180
rect 222988 6140 239404 6168
rect 222988 6128 222994 6140
rect 239398 6128 239404 6140
rect 239456 6128 239462 6180
rect 240778 6128 240784 6180
rect 240836 6168 240842 6180
rect 254118 6168 254124 6180
rect 240836 6140 254124 6168
rect 240836 6128 240842 6140
rect 254118 6128 254124 6140
rect 254176 6128 254182 6180
rect 321097 6171 321155 6177
rect 321097 6137 321109 6171
rect 321143 6168 321155 6171
rect 321143 6140 331260 6168
rect 321143 6137 321155 6140
rect 321097 6131 321155 6137
rect 331232 6032 331260 6140
rect 333238 6128 333244 6180
rect 333296 6168 333302 6180
rect 347866 6168 347872 6180
rect 333296 6140 347872 6168
rect 333296 6128 333302 6140
rect 347866 6128 347872 6140
rect 347924 6128 347930 6180
rect 357158 6128 357164 6180
rect 357216 6168 357222 6180
rect 383470 6168 383476 6180
rect 357216 6140 383476 6168
rect 357216 6128 357222 6140
rect 383470 6128 383476 6140
rect 383528 6128 383534 6180
rect 383562 6128 383568 6180
rect 383620 6168 383626 6180
rect 419166 6168 419172 6180
rect 383620 6140 419172 6168
rect 383620 6128 383626 6140
rect 419166 6128 419172 6140
rect 419224 6128 419230 6180
rect 434622 6128 434628 6180
rect 434680 6168 434686 6180
rect 490558 6168 490564 6180
rect 434680 6140 490564 6168
rect 434680 6128 434686 6140
rect 490558 6128 490564 6140
rect 490616 6128 490622 6180
rect 502978 6128 502984 6180
rect 503036 6168 503042 6180
rect 561950 6168 561956 6180
rect 503036 6140 561956 6168
rect 503036 6128 503042 6140
rect 561950 6128 561956 6140
rect 562008 6128 562014 6180
rect 333606 6032 333612 6044
rect 331232 6004 333612 6032
rect 333606 5992 333612 6004
rect 333664 5992 333670 6044
rect 433334 5992 433340 6044
rect 433392 6032 433398 6044
rect 434622 6032 434628 6044
rect 433392 6004 434628 6032
rect 433392 5992 433398 6004
rect 434622 5992 434628 6004
rect 434680 5992 434686 6044
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 8938 5556 8944 5568
rect 1728 5528 8944 5556
rect 1728 5516 1734 5528
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 326338 5448 326344 5500
rect 326396 5488 326402 5500
rect 330018 5488 330024 5500
rect 326396 5460 330024 5488
rect 326396 5448 326402 5460
rect 330018 5448 330024 5460
rect 330076 5448 330082 5500
rect 165890 4836 165896 4888
rect 165948 4876 165954 4888
rect 167638 4876 167644 4888
rect 165948 4848 167644 4876
rect 165948 4836 165954 4848
rect 167638 4836 167644 4848
rect 167696 4836 167702 4888
rect 201494 4836 201500 4888
rect 201552 4876 201558 4888
rect 226334 4876 226340 4888
rect 201552 4848 226340 4876
rect 201552 4836 201558 4848
rect 226334 4836 226340 4848
rect 226392 4836 226398 4888
rect 310238 4836 310244 4888
rect 310296 4876 310302 4888
rect 318058 4876 318064 4888
rect 310296 4848 318064 4876
rect 310296 4836 310302 4848
rect 318058 4836 318064 4848
rect 318116 4836 318122 4888
rect 376018 4836 376024 4888
rect 376076 4876 376082 4888
rect 401318 4876 401324 4888
rect 376076 4848 401324 4876
rect 376076 4836 376082 4848
rect 401318 4836 401324 4848
rect 401376 4836 401382 4888
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 81434 4808 81440 4820
rect 1452 4780 81440 4808
rect 1452 4768 1458 4780
rect 81434 4768 81440 4780
rect 81492 4768 81498 4820
rect 99282 4768 99288 4820
rect 99340 4808 99346 4820
rect 124858 4808 124864 4820
rect 99340 4780 124864 4808
rect 99340 4768 99346 4780
rect 124858 4768 124864 4780
rect 124916 4768 124922 4820
rect 126606 4768 126612 4820
rect 126664 4808 126670 4820
rect 172514 4808 172520 4820
rect 126664 4780 172520 4808
rect 126664 4768 126670 4780
rect 172514 4768 172520 4780
rect 172572 4768 172578 4820
rect 172974 4768 172980 4820
rect 173032 4808 173038 4820
rect 203518 4808 203524 4820
rect 173032 4780 203524 4808
rect 173032 4768 173038 4780
rect 203518 4768 203524 4780
rect 203576 4768 203582 4820
rect 226518 4768 226524 4820
rect 226576 4808 226582 4820
rect 244366 4808 244372 4820
rect 226576 4780 244372 4808
rect 226576 4768 226582 4780
rect 244366 4768 244372 4780
rect 244424 4768 244430 4820
rect 244458 4768 244464 4820
rect 244516 4808 244522 4820
rect 256694 4808 256700 4820
rect 244516 4780 256700 4808
rect 244516 4768 244522 4780
rect 256694 4768 256700 4780
rect 256752 4768 256758 4820
rect 335262 4768 335268 4820
rect 335320 4808 335326 4820
rect 351362 4808 351368 4820
rect 335320 4780 351368 4808
rect 335320 4768 335326 4780
rect 351362 4768 351368 4780
rect 351420 4768 351426 4820
rect 353202 4768 353208 4820
rect 353260 4808 353266 4820
rect 376386 4808 376392 4820
rect 353260 4780 376392 4808
rect 353260 4768 353266 4780
rect 376386 4768 376392 4780
rect 376444 4768 376450 4820
rect 387702 4768 387708 4820
rect 387760 4808 387766 4820
rect 425146 4808 425152 4820
rect 387760 4780 425152 4808
rect 387760 4768 387766 4780
rect 425146 4768 425152 4780
rect 425204 4768 425210 4820
rect 428921 4811 428979 4817
rect 428921 4777 428933 4811
rect 428967 4808 428979 4811
rect 483474 4808 483480 4820
rect 428967 4780 483480 4808
rect 428967 4777 428979 4780
rect 428921 4771 428979 4777
rect 483474 4768 483480 4780
rect 483532 4768 483538 4820
rect 507118 4768 507124 4820
rect 507176 4808 507182 4820
rect 544102 4808 544108 4820
rect 507176 4780 544108 4808
rect 507176 4768 507182 4780
rect 544102 4768 544108 4780
rect 544160 4768 544166 4820
rect 545758 4768 545764 4820
rect 545816 4808 545822 4820
rect 579798 4808 579804 4820
rect 545816 4780 579804 4808
rect 545816 4768 545822 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 317230 4700 317236 4752
rect 317288 4740 317294 4752
rect 326430 4740 326436 4752
rect 317288 4712 326436 4740
rect 317288 4700 317294 4712
rect 326430 4700 326436 4712
rect 326488 4700 326494 4752
rect 483658 4156 483664 4208
rect 483716 4196 483722 4208
rect 486970 4196 486976 4208
rect 483716 4168 486976 4196
rect 483716 4156 483722 4168
rect 486970 4156 486976 4168
rect 487028 4156 487034 4208
rect 502426 4156 502432 4208
rect 502484 4196 502490 4208
rect 503622 4196 503628 4208
rect 502484 4168 503628 4196
rect 502484 4156 502490 4168
rect 503622 4156 503628 4168
rect 503680 4156 503686 4208
rect 536926 4156 536932 4208
rect 536984 4196 536990 4208
rect 538122 4196 538128 4208
rect 536984 4168 538128 4196
rect 536984 4156 536990 4168
rect 538122 4156 538128 4168
rect 538180 4156 538186 4208
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 10410 4128 10416 4140
rect 8904 4100 10416 4128
rect 8904 4088 8910 4100
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 13722 4128 13728 4140
rect 12492 4100 13728 4128
rect 12492 4088 12498 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17862 4128 17868 4140
rect 17276 4100 17868 4128
rect 17276 4088 17282 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 19242 4128 19248 4140
rect 18380 4100 19248 4128
rect 18380 4088 18386 4100
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20622 4128 20628 4140
rect 19576 4100 20628 4128
rect 19576 4088 19582 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 24302 4088 24308 4140
rect 24360 4128 24366 4140
rect 24762 4128 24768 4140
rect 24360 4100 24768 4128
rect 24360 4088 24366 4100
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 27890 4088 27896 4140
rect 27948 4128 27954 4140
rect 28902 4128 28908 4140
rect 27948 4100 28908 4128
rect 27948 4088 27954 4100
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 33870 4088 33876 4140
rect 33928 4128 33934 4140
rect 34422 4128 34428 4140
rect 33928 4100 34428 4128
rect 33928 4088 33934 4100
rect 34422 4088 34428 4100
rect 34480 4088 34486 4140
rect 37366 4088 37372 4140
rect 37424 4128 37430 4140
rect 38562 4128 38568 4140
rect 37424 4100 38568 4128
rect 37424 4088 37430 4100
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 42702 4128 42708 4140
rect 42208 4100 42708 4128
rect 42208 4088 42214 4100
rect 42702 4088 42708 4100
rect 42760 4088 42766 4140
rect 44542 4088 44548 4140
rect 44600 4128 44606 4140
rect 45462 4128 45468 4140
rect 44600 4100 45468 4128
rect 44600 4088 44606 4100
rect 45462 4088 45468 4100
rect 45520 4088 45526 4140
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 46992 4100 112208 4128
rect 46992 4088 46998 4100
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 9030 4060 9036 4072
rect 4120 4032 9036 4060
rect 4120 4020 4126 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 112070 4060 112076 4072
rect 43404 4032 112076 4060
rect 43404 4020 43410 4032
rect 112070 4020 112076 4032
rect 112128 4020 112134 4072
rect 112180 4060 112208 4100
rect 113542 4088 113548 4140
rect 113600 4128 113606 4140
rect 114462 4128 114468 4140
rect 113600 4100 114468 4128
rect 113600 4088 113606 4100
rect 114462 4088 114468 4100
rect 114520 4088 114526 4140
rect 115934 4088 115940 4140
rect 115992 4128 115998 4140
rect 117222 4128 117228 4140
rect 115992 4100 117228 4128
rect 115992 4088 115998 4100
rect 117222 4088 117228 4100
rect 117280 4088 117286 4140
rect 149238 4088 149244 4140
rect 149296 4128 149302 4140
rect 150342 4128 150348 4140
rect 149296 4100 150348 4128
rect 149296 4088 149302 4100
rect 150342 4088 150348 4100
rect 150400 4088 150406 4140
rect 153930 4088 153936 4140
rect 153988 4128 153994 4140
rect 154482 4128 154488 4140
rect 153988 4100 154488 4128
rect 153988 4088 153994 4100
rect 154482 4088 154488 4100
rect 154540 4088 154546 4140
rect 158714 4088 158720 4140
rect 158772 4128 158778 4140
rect 159910 4128 159916 4140
rect 158772 4100 159916 4128
rect 158772 4088 158778 4100
rect 159910 4088 159916 4100
rect 159968 4088 159974 4140
rect 163498 4088 163504 4140
rect 163556 4128 163562 4140
rect 164142 4128 164148 4140
rect 163556 4100 164148 4128
rect 163556 4088 163562 4100
rect 164142 4088 164148 4100
rect 164200 4088 164206 4140
rect 166997 4131 167055 4137
rect 166997 4128 167009 4131
rect 164252 4100 167009 4128
rect 114554 4060 114560 4072
rect 112180 4032 114560 4060
rect 114554 4020 114560 4032
rect 114612 4020 114618 4072
rect 125410 4020 125416 4072
rect 125468 4060 125474 4072
rect 164252 4060 164280 4100
rect 166997 4097 167009 4100
rect 167043 4097 167055 4131
rect 166997 4091 167055 4097
rect 167086 4088 167092 4140
rect 167144 4128 167150 4140
rect 168190 4128 168196 4140
rect 167144 4100 168196 4128
rect 167144 4088 167150 4100
rect 168190 4088 168196 4100
rect 168248 4088 168254 4140
rect 170582 4088 170588 4140
rect 170640 4128 170646 4140
rect 171042 4128 171048 4140
rect 170640 4100 171048 4128
rect 170640 4088 170646 4100
rect 171042 4088 171048 4100
rect 171100 4088 171106 4140
rect 174170 4088 174176 4140
rect 174228 4128 174234 4140
rect 175182 4128 175188 4140
rect 174228 4100 175188 4128
rect 174228 4088 174234 4100
rect 175182 4088 175188 4100
rect 175240 4088 175246 4140
rect 235994 4088 236000 4140
rect 236052 4128 236058 4140
rect 251174 4128 251180 4140
rect 236052 4100 251180 4128
rect 236052 4088 236058 4100
rect 251174 4088 251180 4100
rect 251232 4088 251238 4140
rect 252738 4088 252744 4140
rect 252796 4128 252802 4140
rect 262214 4128 262220 4140
rect 252796 4100 262220 4128
rect 252796 4088 252802 4100
rect 262214 4088 262220 4100
rect 262272 4088 262278 4140
rect 271690 4088 271696 4140
rect 271748 4128 271754 4140
rect 276014 4128 276020 4140
rect 271748 4100 276020 4128
rect 271748 4088 271754 4100
rect 276014 4088 276020 4100
rect 276072 4088 276078 4140
rect 277670 4088 277676 4140
rect 277728 4128 277734 4140
rect 280338 4128 280344 4140
rect 277728 4100 280344 4128
rect 277728 4088 277734 4100
rect 280338 4088 280344 4100
rect 280396 4088 280402 4140
rect 284754 4088 284760 4140
rect 284812 4128 284818 4140
rect 285674 4128 285680 4140
rect 284812 4100 285680 4128
rect 284812 4088 284818 4100
rect 285674 4088 285680 4100
rect 285732 4088 285738 4140
rect 288526 4088 288532 4140
rect 288584 4128 288590 4140
rect 289538 4128 289544 4140
rect 288584 4100 289544 4128
rect 288584 4088 288590 4100
rect 289538 4088 289544 4100
rect 289596 4088 289602 4140
rect 289906 4088 289912 4140
rect 289964 4128 289970 4140
rect 290734 4128 290740 4140
rect 289964 4100 290740 4128
rect 289964 4088 289970 4100
rect 290734 4088 290740 4100
rect 290792 4088 290798 4140
rect 291286 4088 291292 4140
rect 291344 4128 291350 4140
rect 291930 4128 291936 4140
rect 291344 4100 291936 4128
rect 291344 4088 291350 4100
rect 291930 4088 291936 4100
rect 291988 4088 291994 4140
rect 295242 4088 295248 4140
rect 295300 4128 295306 4140
rect 296714 4128 296720 4140
rect 295300 4100 296720 4128
rect 295300 4088 295306 4100
rect 296714 4088 296720 4100
rect 296772 4088 296778 4140
rect 303522 4088 303528 4140
rect 303580 4128 303586 4140
rect 307386 4128 307392 4140
rect 303580 4100 307392 4128
rect 303580 4088 303586 4100
rect 307386 4088 307392 4100
rect 307444 4088 307450 4140
rect 402882 4088 402888 4140
rect 402940 4128 402946 4140
rect 446582 4128 446588 4140
rect 402940 4100 446588 4128
rect 402940 4088 402946 4100
rect 446582 4088 446588 4100
rect 446640 4088 446646 4140
rect 474642 4088 474648 4140
rect 474700 4128 474706 4140
rect 546494 4128 546500 4140
rect 474700 4100 546500 4128
rect 474700 4088 474706 4100
rect 546494 4088 546500 4100
rect 546552 4088 546558 4140
rect 168374 4060 168380 4072
rect 125468 4032 164280 4060
rect 164344 4032 168380 4060
rect 125468 4020 125474 4032
rect 36170 3952 36176 4004
rect 36228 3992 36234 4004
rect 107654 3992 107660 4004
rect 36228 3964 107660 3992
rect 36228 3952 36234 3964
rect 107654 3952 107660 3964
rect 107712 3952 107718 4004
rect 121822 3952 121828 4004
rect 121880 3992 121886 4004
rect 164344 3992 164372 4032
rect 168374 4020 168380 4032
rect 168432 4020 168438 4072
rect 200390 4020 200396 4072
rect 200448 4060 200454 4072
rect 225046 4060 225052 4072
rect 200448 4032 225052 4060
rect 200448 4020 200454 4032
rect 225046 4020 225052 4032
rect 225104 4020 225110 4072
rect 227806 4020 227812 4072
rect 227864 4060 227870 4072
rect 244274 4060 244280 4072
rect 227864 4032 244280 4060
rect 227864 4020 227870 4032
rect 244274 4020 244280 4032
rect 244332 4020 244338 4072
rect 249150 4020 249156 4072
rect 249208 4060 249214 4072
rect 259454 4060 259460 4072
rect 249208 4032 259460 4060
rect 249208 4020 249214 4032
rect 259454 4020 259460 4032
rect 259512 4020 259518 4072
rect 275278 4020 275284 4072
rect 275336 4060 275342 4072
rect 278682 4060 278688 4072
rect 275336 4032 278688 4060
rect 275336 4020 275342 4032
rect 278682 4020 278688 4032
rect 278740 4020 278746 4072
rect 278866 4020 278872 4072
rect 278924 4060 278930 4072
rect 281534 4060 281540 4072
rect 278924 4032 281540 4060
rect 278924 4020 278930 4032
rect 281534 4020 281540 4032
rect 281592 4020 281598 4072
rect 282454 4020 282460 4072
rect 282512 4060 282518 4072
rect 284294 4060 284300 4072
rect 282512 4032 284300 4060
rect 282512 4020 282518 4032
rect 284294 4020 284300 4032
rect 284352 4020 284358 4072
rect 296622 4020 296628 4072
rect 296680 4060 296686 4072
rect 297910 4060 297916 4072
rect 296680 4032 297916 4060
rect 296680 4020 296686 4032
rect 297910 4020 297916 4032
rect 297968 4020 297974 4072
rect 306282 4020 306288 4072
rect 306340 4060 306346 4072
rect 310974 4060 310980 4072
rect 306340 4032 310980 4060
rect 306340 4020 306346 4032
rect 310974 4020 310980 4032
rect 311032 4020 311038 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 322842 4060 322848 4072
rect 314620 4032 322848 4060
rect 314620 4020 314626 4032
rect 322842 4020 322848 4032
rect 322900 4020 322906 4072
rect 408402 4020 408408 4072
rect 408460 4060 408466 4072
rect 453666 4060 453672 4072
rect 408460 4032 453672 4060
rect 408460 4020 408466 4032
rect 453666 4020 453672 4032
rect 453724 4020 453730 4072
rect 477402 4020 477408 4072
rect 477460 4060 477466 4072
rect 550082 4060 550088 4072
rect 477460 4032 550088 4060
rect 477460 4020 477466 4032
rect 550082 4020 550088 4032
rect 550140 4020 550146 4072
rect 121880 3964 164372 3992
rect 121880 3952 121886 3964
rect 203886 3952 203892 4004
rect 203944 3992 203950 4004
rect 227714 3992 227720 4004
rect 203944 3964 227720 3992
rect 203944 3952 203950 3964
rect 227714 3952 227720 3964
rect 227772 3952 227778 4004
rect 231302 3952 231308 4004
rect 231360 3992 231366 4004
rect 247034 3992 247040 4004
rect 231360 3964 247040 3992
rect 231360 3952 231366 3964
rect 247034 3952 247040 3964
rect 247092 3952 247098 4004
rect 247954 3952 247960 4004
rect 248012 3992 248018 4004
rect 259546 3992 259552 4004
rect 248012 3964 259552 3992
rect 248012 3952 248018 3964
rect 259546 3952 259552 3964
rect 259604 3952 259610 4004
rect 304902 3952 304908 4004
rect 304960 3992 304966 4004
rect 309778 3992 309784 4004
rect 304960 3964 309784 3992
rect 304960 3952 304966 3964
rect 309778 3952 309784 3964
rect 309836 3952 309842 4004
rect 313090 3952 313096 4004
rect 313148 3992 313154 4004
rect 320450 3992 320456 4004
rect 313148 3964 320456 3992
rect 313148 3952 313154 3964
rect 320450 3952 320456 3964
rect 320508 3952 320514 4004
rect 321462 3952 321468 4004
rect 321520 3992 321526 4004
rect 332410 3992 332416 4004
rect 321520 3964 332416 3992
rect 321520 3952 321526 3964
rect 332410 3952 332416 3964
rect 332468 3952 332474 4004
rect 346302 3952 346308 4004
rect 346360 3992 346366 4004
rect 368014 3992 368020 4004
rect 346360 3964 368020 3992
rect 346360 3952 346366 3964
rect 368014 3952 368020 3964
rect 368072 3952 368078 4004
rect 405642 3952 405648 4004
rect 405700 3992 405706 4004
rect 450170 3992 450176 4004
rect 405700 3964 450176 3992
rect 405700 3952 405706 3964
rect 450170 3952 450176 3964
rect 450228 3952 450234 4004
rect 480162 3952 480168 4004
rect 480220 3992 480226 4004
rect 553578 3992 553584 4004
rect 480220 3964 553584 3992
rect 480220 3952 480226 3964
rect 553578 3952 553584 3964
rect 553636 3952 553642 4004
rect 39758 3884 39764 3936
rect 39816 3924 39822 3936
rect 110414 3924 110420 3936
rect 39816 3896 110420 3924
rect 39816 3884 39822 3896
rect 110414 3884 110420 3896
rect 110472 3884 110478 3936
rect 118234 3884 118240 3936
rect 118292 3924 118298 3936
rect 157337 3927 157395 3933
rect 157337 3924 157349 3927
rect 118292 3896 157349 3924
rect 118292 3884 118298 3896
rect 157337 3893 157349 3896
rect 157383 3893 157395 3927
rect 164234 3924 164240 3936
rect 157337 3887 157395 3893
rect 157444 3896 164240 3924
rect 29086 3816 29092 3868
rect 29144 3856 29150 3868
rect 30282 3856 30288 3868
rect 29144 3828 30288 3856
rect 29144 3816 29150 3828
rect 30282 3816 30288 3828
rect 30340 3816 30346 3868
rect 32674 3816 32680 3868
rect 32732 3856 32738 3868
rect 32732 3828 99512 3856
rect 32732 3816 32738 3828
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 99374 3788 99380 3800
rect 25556 3760 99380 3788
rect 25556 3748 25562 3760
rect 99374 3748 99380 3760
rect 99432 3748 99438 3800
rect 99484 3788 99512 3828
rect 114738 3816 114744 3868
rect 114796 3856 114802 3868
rect 157444 3856 157472 3896
rect 164234 3884 164240 3896
rect 164292 3884 164298 3936
rect 166997 3927 167055 3933
rect 166997 3893 167009 3927
rect 167043 3924 167055 3927
rect 171318 3924 171324 3936
rect 167043 3896 171324 3924
rect 167043 3893 167055 3896
rect 166997 3887 167055 3893
rect 171318 3884 171324 3896
rect 171376 3884 171382 3936
rect 193214 3884 193220 3936
rect 193272 3924 193278 3936
rect 219526 3924 219532 3936
rect 193272 3896 219532 3924
rect 193272 3884 193278 3896
rect 219526 3884 219532 3896
rect 219584 3884 219590 3936
rect 225322 3884 225328 3936
rect 225380 3924 225386 3936
rect 242894 3924 242900 3936
rect 225380 3896 242900 3924
rect 225380 3884 225386 3896
rect 242894 3884 242900 3896
rect 242952 3884 242958 3936
rect 243170 3884 243176 3936
rect 243228 3924 243234 3936
rect 255406 3924 255412 3936
rect 243228 3896 255412 3924
rect 243228 3884 243234 3896
rect 255406 3884 255412 3896
rect 255464 3884 255470 3936
rect 259822 3884 259828 3936
rect 259880 3924 259886 3936
rect 267734 3924 267740 3936
rect 259880 3896 267740 3924
rect 259880 3884 259886 3896
rect 267734 3884 267740 3896
rect 267792 3884 267798 3936
rect 303430 3884 303436 3936
rect 303488 3924 303494 3936
rect 308582 3924 308588 3936
rect 303488 3896 308588 3924
rect 303488 3884 303494 3896
rect 308582 3884 308588 3896
rect 308640 3884 308646 3936
rect 311802 3884 311808 3936
rect 311860 3924 311866 3936
rect 319254 3924 319260 3936
rect 311860 3896 319260 3924
rect 311860 3884 311866 3896
rect 319254 3884 319260 3896
rect 319312 3884 319318 3936
rect 324222 3884 324228 3936
rect 324280 3924 324286 3936
rect 335906 3924 335912 3936
rect 324280 3896 335912 3924
rect 324280 3884 324286 3896
rect 335906 3884 335912 3896
rect 335964 3884 335970 3936
rect 343542 3884 343548 3936
rect 343600 3924 343606 3936
rect 364518 3924 364524 3936
rect 343600 3896 364524 3924
rect 343600 3884 343606 3896
rect 364518 3884 364524 3896
rect 364576 3884 364582 3936
rect 371602 3924 371608 3936
rect 365640 3896 371608 3924
rect 114796 3828 157472 3856
rect 114796 3816 114802 3828
rect 157518 3816 157524 3868
rect 157576 3856 157582 3868
rect 158622 3856 158628 3868
rect 157576 3828 158628 3856
rect 157576 3816 157582 3828
rect 158622 3816 158628 3828
rect 158680 3816 158686 3868
rect 196802 3816 196808 3868
rect 196860 3856 196866 3868
rect 222194 3856 222200 3868
rect 196860 3828 222200 3856
rect 196860 3816 196866 3828
rect 222194 3816 222200 3828
rect 222252 3816 222258 3868
rect 228910 3816 228916 3868
rect 228968 3856 228974 3868
rect 245654 3856 245660 3868
rect 228968 3828 245660 3856
rect 228968 3816 228974 3828
rect 245654 3816 245660 3828
rect 245712 3816 245718 3868
rect 246758 3816 246764 3868
rect 246816 3856 246822 3868
rect 258350 3856 258356 3868
rect 246816 3828 258356 3856
rect 246816 3816 246822 3828
rect 258350 3816 258356 3828
rect 258408 3816 258414 3868
rect 262214 3816 262220 3868
rect 262272 3856 262278 3868
rect 269298 3856 269304 3868
rect 262272 3828 269304 3856
rect 262272 3816 262278 3828
rect 269298 3816 269304 3828
rect 269356 3816 269362 3868
rect 328362 3816 328368 3868
rect 328420 3856 328426 3868
rect 341886 3856 341892 3868
rect 328420 3828 341892 3856
rect 328420 3816 328426 3828
rect 341886 3816 341892 3828
rect 341944 3816 341950 3868
rect 349062 3816 349068 3868
rect 349120 3856 349126 3868
rect 365640 3856 365668 3896
rect 371602 3884 371608 3896
rect 371660 3884 371666 3936
rect 411162 3884 411168 3936
rect 411220 3924 411226 3936
rect 457254 3924 457260 3936
rect 411220 3896 457260 3924
rect 411220 3884 411226 3896
rect 457254 3884 457260 3896
rect 457312 3884 457318 3936
rect 482922 3884 482928 3936
rect 482980 3924 482986 3936
rect 557166 3924 557172 3936
rect 482980 3896 557172 3924
rect 482980 3884 482986 3896
rect 557166 3884 557172 3896
rect 557224 3884 557230 3936
rect 349120 3828 365668 3856
rect 349120 3816 349126 3828
rect 365714 3816 365720 3868
rect 365772 3856 365778 3868
rect 366910 3856 366916 3868
rect 365772 3828 366916 3856
rect 365772 3816 365778 3828
rect 366910 3816 366916 3828
rect 366968 3816 366974 3868
rect 413922 3816 413928 3868
rect 413980 3856 413986 3868
rect 460842 3856 460848 3868
rect 413980 3828 460848 3856
rect 413980 3816 413986 3828
rect 460842 3816 460848 3828
rect 460900 3816 460906 3868
rect 485682 3816 485688 3868
rect 485740 3856 485746 3868
rect 560754 3856 560760 3868
rect 485740 3828 560760 3856
rect 485740 3816 485746 3828
rect 560754 3816 560760 3828
rect 560812 3816 560818 3868
rect 104894 3788 104900 3800
rect 99484 3760 104900 3788
rect 104894 3748 104900 3760
rect 104952 3748 104958 3800
rect 111150 3748 111156 3800
rect 111208 3788 111214 3800
rect 161474 3788 161480 3800
rect 111208 3760 161480 3788
rect 111208 3748 111214 3760
rect 161474 3748 161480 3760
rect 161532 3748 161538 3800
rect 189626 3748 189632 3800
rect 189684 3788 189690 3800
rect 218054 3788 218060 3800
rect 189684 3760 218060 3788
rect 189684 3748 189690 3760
rect 218054 3748 218060 3760
rect 218112 3748 218118 3800
rect 241974 3748 241980 3800
rect 242032 3788 242038 3800
rect 255314 3788 255320 3800
rect 242032 3760 255320 3788
rect 242032 3748 242038 3760
rect 255314 3748 255320 3760
rect 255372 3748 255378 3800
rect 256234 3748 256240 3800
rect 256292 3788 256298 3800
rect 264974 3788 264980 3800
rect 256292 3760 264980 3788
rect 256292 3748 256298 3760
rect 264974 3748 264980 3760
rect 265032 3748 265038 3800
rect 276474 3748 276480 3800
rect 276532 3788 276538 3800
rect 280154 3788 280160 3800
rect 276532 3760 280160 3788
rect 276532 3748 276538 3760
rect 280154 3748 280160 3760
rect 280212 3748 280218 3800
rect 317322 3748 317328 3800
rect 317380 3788 317386 3800
rect 327626 3788 327632 3800
rect 317380 3760 327632 3788
rect 317380 3748 317386 3760
rect 327626 3748 327632 3760
rect 327684 3748 327690 3800
rect 328086 3748 328092 3800
rect 328144 3788 328150 3800
rect 343082 3788 343088 3800
rect 328144 3760 343088 3788
rect 328144 3748 328150 3760
rect 343082 3748 343088 3760
rect 343140 3748 343146 3800
rect 351822 3748 351828 3800
rect 351880 3788 351886 3800
rect 375190 3788 375196 3800
rect 351880 3760 375196 3788
rect 351880 3748 351886 3760
rect 375190 3748 375196 3760
rect 375248 3748 375254 3800
rect 415118 3748 415124 3800
rect 415176 3788 415182 3800
rect 464430 3788 464436 3800
rect 415176 3760 464436 3788
rect 415176 3748 415182 3760
rect 464430 3748 464436 3760
rect 464488 3748 464494 3800
rect 487062 3748 487068 3800
rect 487120 3788 487126 3800
rect 564342 3788 564348 3800
rect 487120 3760 564348 3788
rect 487120 3748 487126 3760
rect 564342 3748 564348 3760
rect 564400 3748 564406 3800
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 96614 3720 96620 3732
rect 20772 3692 96620 3720
rect 20772 3680 20778 3692
rect 96614 3680 96620 3692
rect 96672 3680 96678 3732
rect 107470 3680 107476 3732
rect 107528 3720 107534 3732
rect 158806 3720 158812 3732
rect 107528 3692 158812 3720
rect 107528 3680 107534 3692
rect 158806 3680 158812 3692
rect 158864 3680 158870 3732
rect 186038 3680 186044 3732
rect 186096 3720 186102 3732
rect 215294 3720 215300 3732
rect 186096 3692 215300 3720
rect 186096 3680 186102 3692
rect 215294 3680 215300 3692
rect 215352 3680 215358 3732
rect 218146 3680 218152 3732
rect 218204 3720 218210 3732
rect 237374 3720 237380 3732
rect 218204 3692 237380 3720
rect 218204 3680 218210 3692
rect 237374 3680 237380 3692
rect 237432 3680 237438 3732
rect 239582 3680 239588 3732
rect 239640 3720 239646 3732
rect 252646 3720 252652 3732
rect 239640 3692 252652 3720
rect 239640 3680 239646 3692
rect 252646 3680 252652 3692
rect 252704 3680 252710 3732
rect 257430 3680 257436 3732
rect 257488 3720 257494 3732
rect 266354 3720 266360 3732
rect 257488 3692 266360 3720
rect 257488 3680 257494 3692
rect 266354 3680 266360 3692
rect 266412 3680 266418 3732
rect 269298 3680 269304 3732
rect 269356 3720 269362 3732
rect 274634 3720 274640 3732
rect 269356 3692 274640 3720
rect 269356 3680 269362 3692
rect 274634 3680 274640 3692
rect 274692 3680 274698 3732
rect 318702 3680 318708 3732
rect 318760 3720 318766 3732
rect 328822 3720 328828 3732
rect 318760 3692 328828 3720
rect 318760 3680 318766 3692
rect 328822 3680 328828 3692
rect 328880 3680 328886 3732
rect 331122 3680 331128 3732
rect 331180 3720 331186 3732
rect 346670 3720 346676 3732
rect 331180 3692 346676 3720
rect 331180 3680 331186 3692
rect 346670 3680 346676 3692
rect 346728 3680 346734 3732
rect 354582 3680 354588 3732
rect 354640 3720 354646 3732
rect 378778 3720 378784 3732
rect 354640 3692 378784 3720
rect 354640 3680 354646 3692
rect 378778 3680 378784 3692
rect 378836 3680 378842 3732
rect 420822 3680 420828 3732
rect 420880 3720 420886 3732
rect 471514 3720 471520 3732
rect 420880 3692 471520 3720
rect 420880 3680 420886 3692
rect 471514 3680 471520 3692
rect 471572 3680 471578 3732
rect 489822 3680 489828 3732
rect 489880 3720 489886 3732
rect 567838 3720 567844 3732
rect 489880 3692 567844 3720
rect 489880 3680 489886 3692
rect 567838 3680 567844 3692
rect 567896 3680 567902 3732
rect 16022 3612 16028 3664
rect 16080 3652 16086 3664
rect 92474 3652 92480 3664
rect 16080 3624 92480 3652
rect 16080 3612 16086 3624
rect 92474 3612 92480 3624
rect 92532 3612 92538 3664
rect 103974 3612 103980 3664
rect 104032 3652 104038 3664
rect 155954 3652 155960 3664
rect 104032 3624 155960 3652
rect 104032 3612 104038 3624
rect 155954 3612 155960 3624
rect 156012 3612 156018 3664
rect 157337 3655 157395 3661
rect 157337 3621 157349 3655
rect 157383 3652 157395 3655
rect 165798 3652 165804 3664
rect 157383 3624 165804 3652
rect 157383 3621 157395 3624
rect 157337 3615 157395 3621
rect 165798 3612 165804 3624
rect 165856 3612 165862 3664
rect 182542 3612 182548 3664
rect 182600 3652 182606 3664
rect 212534 3652 212540 3664
rect 182600 3624 212540 3652
rect 182600 3612 182606 3624
rect 212534 3612 212540 3624
rect 212592 3612 212598 3664
rect 221734 3612 221740 3664
rect 221792 3652 221798 3664
rect 240134 3652 240140 3664
rect 221792 3624 240140 3652
rect 221792 3612 221798 3624
rect 240134 3612 240140 3624
rect 240192 3612 240198 3664
rect 245562 3612 245568 3664
rect 245620 3652 245626 3664
rect 258074 3652 258080 3664
rect 245620 3624 258080 3652
rect 245620 3612 245626 3624
rect 258074 3612 258080 3624
rect 258132 3612 258138 3664
rect 268102 3612 268108 3664
rect 268160 3652 268166 3664
rect 273254 3652 273260 3664
rect 268160 3624 273260 3652
rect 268160 3612 268166 3624
rect 273254 3612 273260 3624
rect 273312 3612 273318 3664
rect 320082 3612 320088 3664
rect 320140 3652 320146 3664
rect 331214 3652 331220 3664
rect 320140 3624 331220 3652
rect 320140 3612 320146 3624
rect 331214 3612 331220 3624
rect 331272 3612 331278 3664
rect 333882 3612 333888 3664
rect 333940 3652 333946 3664
rect 350258 3652 350264 3664
rect 333940 3624 350264 3652
rect 333940 3612 333946 3624
rect 350258 3612 350264 3624
rect 350316 3612 350322 3664
rect 357342 3612 357348 3664
rect 357400 3612 357406 3664
rect 360102 3612 360108 3664
rect 360160 3652 360166 3664
rect 385862 3652 385868 3664
rect 360160 3624 385868 3652
rect 360160 3612 360166 3624
rect 385862 3612 385868 3624
rect 385920 3612 385926 3664
rect 418062 3612 418068 3664
rect 418120 3652 418126 3664
rect 467834 3652 467840 3664
rect 418120 3624 467840 3652
rect 418120 3612 418126 3624
rect 467834 3612 467840 3624
rect 467892 3612 467898 3664
rect 492582 3612 492588 3664
rect 492640 3652 492646 3664
rect 571334 3652 571340 3664
rect 492640 3624 571340 3652
rect 492640 3612 492646 3624
rect 571334 3612 571340 3624
rect 571392 3612 571398 3664
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10962 3584 10968 3596
rect 10100 3556 10968 3584
rect 10100 3544 10106 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 89714 3584 89720 3596
rect 11296 3556 89720 3584
rect 11296 3544 11302 3556
rect 89714 3544 89720 3556
rect 89772 3544 89778 3596
rect 100478 3544 100484 3596
rect 100536 3584 100542 3596
rect 102229 3587 102287 3593
rect 100536 3556 102180 3584
rect 100536 3544 100542 3556
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6512 3488 74672 3516
rect 6512 3476 6518 3488
rect 38580 3420 45692 3448
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 5316 3352 9689 3380
rect 5316 3340 5322 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 22189 3383 22247 3389
rect 22189 3349 22201 3383
rect 22235 3380 22247 3383
rect 31665 3383 31723 3389
rect 31665 3380 31677 3383
rect 22235 3352 31677 3380
rect 22235 3349 22247 3352
rect 22189 3343 22247 3349
rect 31665 3349 31677 3352
rect 31711 3349 31723 3383
rect 31665 3343 31723 3349
rect 31849 3383 31907 3389
rect 31849 3349 31861 3383
rect 31895 3380 31907 3383
rect 38580 3380 38608 3420
rect 31895 3352 38608 3380
rect 31895 3349 31907 3352
rect 31849 3343 31907 3349
rect 19245 3315 19303 3321
rect 19245 3281 19257 3315
rect 19291 3312 19303 3315
rect 22005 3315 22063 3321
rect 22005 3312 22017 3315
rect 19291 3284 22017 3312
rect 19291 3281 19303 3284
rect 19245 3275 19303 3281
rect 22005 3281 22017 3284
rect 22051 3281 22063 3315
rect 45664 3312 45692 3420
rect 45738 3408 45744 3460
rect 45796 3448 45802 3460
rect 46842 3448 46848 3460
rect 45796 3420 46848 3448
rect 45796 3408 45802 3420
rect 46842 3408 46848 3420
rect 46900 3408 46906 3460
rect 50522 3408 50528 3460
rect 50580 3448 50586 3460
rect 50982 3448 50988 3460
rect 50580 3420 50988 3448
rect 50580 3408 50586 3420
rect 50982 3408 50988 3420
rect 51040 3408 51046 3460
rect 51626 3408 51632 3460
rect 51684 3448 51690 3460
rect 52362 3448 52368 3460
rect 51684 3420 52368 3448
rect 51684 3408 51690 3420
rect 52362 3408 52368 3420
rect 52420 3408 52426 3460
rect 52822 3408 52828 3460
rect 52880 3448 52886 3460
rect 53742 3448 53748 3460
rect 52880 3420 53748 3448
rect 52880 3408 52886 3420
rect 53742 3408 53748 3420
rect 53800 3408 53806 3460
rect 54018 3408 54024 3460
rect 54076 3448 54082 3460
rect 55122 3448 55128 3460
rect 54076 3420 55128 3448
rect 54076 3408 54082 3420
rect 55122 3408 55128 3420
rect 55180 3408 55186 3460
rect 68278 3408 68284 3460
rect 68336 3448 68342 3460
rect 68922 3448 68928 3460
rect 68336 3420 68928 3448
rect 68336 3408 68342 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 69474 3408 69480 3460
rect 69532 3448 69538 3460
rect 70302 3448 70308 3460
rect 69532 3420 70308 3448
rect 69532 3408 69538 3420
rect 70302 3408 70308 3420
rect 70360 3408 70366 3460
rect 70670 3408 70676 3460
rect 70728 3448 70734 3460
rect 71682 3448 71688 3460
rect 70728 3420 71688 3448
rect 70728 3408 70734 3420
rect 71682 3408 71688 3420
rect 71740 3408 71746 3460
rect 74644 3448 74672 3488
rect 76650 3476 76656 3528
rect 76708 3516 76714 3528
rect 77202 3516 77208 3528
rect 76708 3488 77208 3516
rect 76708 3476 76714 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 77846 3476 77852 3528
rect 77904 3516 77910 3528
rect 78582 3516 78588 3528
rect 77904 3488 78588 3516
rect 77904 3476 77910 3488
rect 78582 3476 78588 3488
rect 78640 3476 78646 3528
rect 81434 3476 81440 3528
rect 81492 3516 81498 3528
rect 82630 3516 82636 3528
rect 81492 3488 82636 3516
rect 81492 3476 81498 3488
rect 82630 3476 82636 3488
rect 82688 3476 82694 3528
rect 84930 3476 84936 3528
rect 84988 3516 84994 3528
rect 85482 3516 85488 3528
rect 84988 3488 85488 3516
rect 84988 3476 84994 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 86126 3476 86132 3528
rect 86184 3516 86190 3528
rect 86862 3516 86868 3528
rect 86184 3488 86868 3516
rect 86184 3476 86190 3488
rect 86862 3476 86868 3488
rect 86920 3476 86926 3528
rect 88518 3476 88524 3528
rect 88576 3516 88582 3528
rect 89622 3516 89628 3528
rect 88576 3488 89628 3516
rect 88576 3476 88582 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 94498 3476 94504 3528
rect 94556 3516 94562 3528
rect 95142 3516 95148 3528
rect 94556 3488 95148 3516
rect 94556 3476 94562 3488
rect 95142 3476 95148 3488
rect 95200 3476 95206 3528
rect 95694 3476 95700 3528
rect 95752 3516 95758 3528
rect 96522 3516 96528 3528
rect 95752 3488 96528 3516
rect 95752 3476 95758 3488
rect 96522 3476 96528 3488
rect 96580 3476 96586 3528
rect 98086 3476 98092 3528
rect 98144 3516 98150 3528
rect 99190 3516 99196 3528
rect 98144 3488 99196 3516
rect 98144 3476 98150 3488
rect 99190 3476 99196 3488
rect 99248 3476 99254 3528
rect 101582 3476 101588 3528
rect 101640 3516 101646 3528
rect 102042 3516 102048 3528
rect 101640 3488 102048 3516
rect 101640 3476 101646 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 102152 3516 102180 3556
rect 102229 3553 102241 3587
rect 102275 3584 102287 3587
rect 150342 3584 150348 3596
rect 102275 3556 150348 3584
rect 102275 3553 102287 3556
rect 102229 3547 102287 3553
rect 150342 3544 150348 3556
rect 150400 3544 150406 3596
rect 175366 3544 175372 3596
rect 175424 3584 175430 3596
rect 207106 3584 207112 3596
rect 175424 3556 207112 3584
rect 175424 3544 175430 3556
rect 207106 3544 207112 3556
rect 207164 3544 207170 3596
rect 207474 3544 207480 3596
rect 207532 3584 207538 3596
rect 230474 3584 230480 3596
rect 207532 3556 230480 3584
rect 207532 3544 207538 3556
rect 230474 3544 230480 3556
rect 230532 3544 230538 3596
rect 232498 3544 232504 3596
rect 232556 3584 232562 3596
rect 248414 3584 248420 3596
rect 232556 3556 248420 3584
rect 232556 3544 232562 3556
rect 248414 3544 248420 3556
rect 248472 3544 248478 3596
rect 251450 3544 251456 3596
rect 251508 3584 251514 3596
rect 262306 3584 262312 3596
rect 251508 3556 262312 3584
rect 251508 3544 251514 3556
rect 262306 3544 262312 3556
rect 262364 3544 262370 3596
rect 263410 3544 263416 3596
rect 263468 3584 263474 3596
rect 263468 3556 264560 3584
rect 263468 3544 263474 3556
rect 102152 3488 145604 3516
rect 85761 3451 85819 3457
rect 85761 3448 85773 3451
rect 71792 3420 74580 3448
rect 74644 3420 85773 3448
rect 58802 3340 58808 3392
rect 58860 3380 58866 3392
rect 59262 3380 59268 3392
rect 58860 3352 59268 3380
rect 58860 3340 58866 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 62390 3340 62396 3392
rect 62448 3380 62454 3392
rect 63402 3380 63408 3392
rect 62448 3352 63408 3380
rect 62448 3340 62454 3352
rect 63402 3340 63408 3352
rect 63460 3340 63466 3392
rect 71792 3380 71820 3420
rect 74552 3380 74580 3420
rect 85761 3417 85773 3420
rect 85807 3417 85819 3451
rect 85761 3411 85819 3417
rect 93302 3408 93308 3460
rect 93360 3448 93366 3460
rect 145576 3448 145604 3488
rect 145650 3476 145656 3528
rect 145708 3516 145714 3528
rect 146202 3516 146208 3528
rect 145708 3488 146208 3516
rect 145708 3476 145714 3488
rect 146202 3476 146208 3488
rect 146260 3476 146266 3528
rect 146846 3476 146852 3528
rect 146904 3516 146910 3528
rect 147582 3516 147588 3528
rect 146904 3488 147588 3516
rect 146904 3476 146910 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 150434 3476 150440 3528
rect 150492 3516 150498 3528
rect 151722 3516 151728 3528
rect 150492 3488 151728 3516
rect 150492 3476 150498 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 164694 3476 164700 3528
rect 164752 3516 164758 3528
rect 165522 3516 165528 3528
rect 164752 3488 165528 3516
rect 164752 3476 164758 3488
rect 165522 3476 165528 3488
rect 165580 3476 165586 3528
rect 178954 3476 178960 3528
rect 179012 3516 179018 3528
rect 209958 3516 209964 3528
rect 179012 3488 209964 3516
rect 179012 3476 179018 3488
rect 209958 3476 209964 3488
rect 210016 3476 210022 3528
rect 224865 3519 224923 3525
rect 224865 3485 224877 3519
rect 224911 3516 224923 3519
rect 224957 3519 225015 3525
rect 224957 3516 224969 3519
rect 224911 3488 224969 3516
rect 224911 3485 224923 3488
rect 224865 3479 224923 3485
rect 224957 3485 224969 3488
rect 225003 3485 225015 3519
rect 236178 3516 236184 3528
rect 224957 3479 225015 3485
rect 234724 3488 236184 3516
rect 153470 3448 153476 3460
rect 93360 3420 145052 3448
rect 145576 3420 153476 3448
rect 93360 3408 93366 3420
rect 63512 3352 71820 3380
rect 74460 3352 74580 3380
rect 63512 3312 63540 3352
rect 45664 3284 63540 3312
rect 22005 3275 22063 3281
rect 63586 3272 63592 3324
rect 63644 3312 63650 3324
rect 64782 3312 64788 3324
rect 63644 3284 64788 3312
rect 63644 3272 63650 3284
rect 64782 3272 64788 3284
rect 64840 3272 64846 3324
rect 55214 3204 55220 3256
rect 55272 3244 55278 3256
rect 56502 3244 56508 3256
rect 55272 3216 56508 3244
rect 55272 3204 55278 3216
rect 56502 3204 56508 3216
rect 56560 3204 56566 3256
rect 74460 3244 74488 3352
rect 96890 3340 96896 3392
rect 96948 3380 96954 3392
rect 102229 3383 102287 3389
rect 102229 3380 102241 3383
rect 96948 3352 102241 3380
rect 96948 3340 96954 3352
rect 102229 3349 102241 3352
rect 102275 3349 102287 3383
rect 102229 3343 102287 3349
rect 105170 3340 105176 3392
rect 105228 3380 105234 3392
rect 106182 3380 106188 3392
rect 105228 3352 106188 3380
rect 105228 3340 105234 3352
rect 106182 3340 106188 3352
rect 106240 3340 106246 3392
rect 106366 3340 106372 3392
rect 106424 3380 106430 3392
rect 107562 3380 107568 3392
rect 106424 3352 107568 3380
rect 106424 3340 106430 3352
rect 107562 3340 107568 3352
rect 107620 3340 107626 3392
rect 119430 3340 119436 3392
rect 119488 3380 119494 3392
rect 119982 3380 119988 3392
rect 119488 3352 119988 3380
rect 119488 3340 119494 3352
rect 119982 3340 119988 3352
rect 120040 3340 120046 3392
rect 120626 3340 120632 3392
rect 120684 3380 120690 3392
rect 121362 3380 121368 3392
rect 120684 3352 121368 3380
rect 120684 3340 120690 3352
rect 121362 3340 121368 3352
rect 121420 3340 121426 3392
rect 123018 3340 123024 3392
rect 123076 3380 123082 3392
rect 124122 3380 124128 3392
rect 123076 3352 124128 3380
rect 123076 3340 123082 3352
rect 124122 3340 124128 3352
rect 124180 3340 124186 3392
rect 124214 3340 124220 3392
rect 124272 3380 124278 3392
rect 125502 3380 125508 3392
rect 124272 3352 125508 3380
rect 124272 3340 124278 3352
rect 125502 3340 125508 3352
rect 125560 3340 125566 3392
rect 127802 3340 127808 3392
rect 127860 3380 127866 3392
rect 128262 3380 128268 3392
rect 127860 3352 128268 3380
rect 127860 3340 127866 3352
rect 128262 3340 128268 3352
rect 128320 3340 128326 3392
rect 128998 3340 129004 3392
rect 129056 3380 129062 3392
rect 129642 3380 129648 3392
rect 129056 3352 129648 3380
rect 129056 3340 129062 3352
rect 129642 3340 129648 3352
rect 129700 3340 129706 3392
rect 131390 3340 131396 3392
rect 131448 3380 131454 3392
rect 132402 3380 132408 3392
rect 131448 3352 132408 3380
rect 131448 3340 131454 3352
rect 132402 3340 132408 3352
rect 132460 3340 132466 3392
rect 136082 3340 136088 3392
rect 136140 3380 136146 3392
rect 136542 3380 136548 3392
rect 136140 3352 136548 3380
rect 136140 3340 136146 3352
rect 136542 3340 136548 3352
rect 136600 3340 136606 3392
rect 137278 3340 137284 3392
rect 137336 3380 137342 3392
rect 137922 3380 137928 3392
rect 137336 3352 137928 3380
rect 137336 3340 137342 3352
rect 137922 3340 137928 3352
rect 137980 3340 137986 3392
rect 138474 3340 138480 3392
rect 138532 3380 138538 3392
rect 139302 3380 139308 3392
rect 138532 3352 139308 3380
rect 138532 3340 138538 3352
rect 139302 3340 139308 3352
rect 139360 3340 139366 3392
rect 139670 3340 139676 3392
rect 139728 3380 139734 3392
rect 140682 3380 140688 3392
rect 139728 3352 140688 3380
rect 139728 3340 139734 3352
rect 140682 3340 140688 3352
rect 140740 3340 140746 3392
rect 140866 3340 140872 3392
rect 140924 3380 140930 3392
rect 141970 3380 141976 3392
rect 140924 3352 141976 3380
rect 140924 3340 140930 3352
rect 141970 3340 141976 3352
rect 142028 3340 142034 3392
rect 145024 3380 145052 3420
rect 153470 3408 153476 3420
rect 153528 3408 153534 3460
rect 171778 3408 171784 3460
rect 171836 3448 171842 3460
rect 204438 3448 204444 3460
rect 171836 3420 204444 3448
rect 171836 3408 171842 3420
rect 204438 3408 204444 3420
rect 204496 3408 204502 3460
rect 209866 3408 209872 3460
rect 209924 3448 209930 3460
rect 211062 3448 211068 3460
rect 209924 3420 211068 3448
rect 209924 3408 209930 3420
rect 211062 3408 211068 3420
rect 211120 3408 211126 3460
rect 233418 3448 233424 3460
rect 211816 3420 233424 3448
rect 148042 3380 148048 3392
rect 145024 3352 148048 3380
rect 148042 3340 148048 3352
rect 148100 3340 148106 3392
rect 188430 3340 188436 3392
rect 188488 3380 188494 3392
rect 188982 3380 188988 3392
rect 188488 3352 188988 3380
rect 188488 3340 188494 3352
rect 188982 3340 188988 3352
rect 189040 3340 189046 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 191742 3380 191748 3392
rect 190880 3352 191748 3380
rect 190880 3340 190886 3352
rect 191742 3340 191748 3352
rect 191800 3340 191806 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 193122 3380 193128 3392
rect 192076 3352 193128 3380
rect 192076 3340 192082 3352
rect 193122 3340 193128 3352
rect 193180 3340 193186 3392
rect 197998 3340 198004 3392
rect 198056 3380 198062 3392
rect 198642 3380 198648 3392
rect 198056 3352 198648 3380
rect 198056 3340 198062 3352
rect 198642 3340 198648 3352
rect 198700 3340 198706 3392
rect 199194 3340 199200 3392
rect 199252 3380 199258 3392
rect 200022 3380 200028 3392
rect 199252 3352 200028 3380
rect 199252 3340 199258 3352
rect 200022 3340 200028 3352
rect 200080 3340 200086 3392
rect 211816 3380 211844 3420
rect 233418 3408 233424 3420
rect 233476 3408 233482 3460
rect 233513 3451 233571 3457
rect 233513 3417 233525 3451
rect 233559 3448 233571 3451
rect 234724 3448 234752 3488
rect 236178 3476 236184 3488
rect 236236 3476 236242 3528
rect 238386 3476 238392 3528
rect 238444 3516 238450 3528
rect 252554 3516 252560 3528
rect 238444 3488 252560 3516
rect 238444 3476 238450 3488
rect 252554 3476 252560 3488
rect 252612 3476 252618 3528
rect 253842 3476 253848 3528
rect 253900 3516 253906 3528
rect 263594 3516 263600 3528
rect 253900 3488 263600 3516
rect 253900 3476 253906 3488
rect 263594 3476 263600 3488
rect 263652 3476 263658 3528
rect 264532 3516 264560 3556
rect 264606 3544 264612 3596
rect 264664 3584 264670 3596
rect 270494 3584 270500 3596
rect 264664 3556 270500 3584
rect 264664 3544 264670 3556
rect 270494 3544 270500 3556
rect 270552 3544 270558 3596
rect 285950 3544 285956 3596
rect 286008 3584 286014 3596
rect 287054 3584 287060 3596
rect 286008 3556 287060 3584
rect 286008 3544 286014 3556
rect 287054 3544 287060 3556
rect 287112 3544 287118 3596
rect 313182 3544 313188 3596
rect 313240 3584 313246 3596
rect 321646 3584 321652 3596
rect 313240 3556 321652 3584
rect 313240 3544 313246 3556
rect 321646 3544 321652 3556
rect 321704 3544 321710 3596
rect 322934 3544 322940 3596
rect 322992 3584 322998 3596
rect 334710 3584 334716 3596
rect 322992 3556 334716 3584
rect 322992 3544 322998 3556
rect 334710 3544 334716 3556
rect 334768 3544 334774 3596
rect 336550 3544 336556 3596
rect 336608 3584 336614 3596
rect 347685 3587 347743 3593
rect 347685 3584 347697 3587
rect 336608 3556 347697 3584
rect 336608 3544 336614 3556
rect 347685 3553 347697 3556
rect 347731 3553 347743 3587
rect 347685 3547 347743 3553
rect 347774 3544 347780 3596
rect 347832 3584 347838 3596
rect 349062 3584 349068 3596
rect 347832 3556 349068 3584
rect 347832 3544 347838 3556
rect 349062 3544 349068 3556
rect 349120 3544 349126 3596
rect 357360 3584 357388 3612
rect 382366 3584 382372 3596
rect 357360 3556 382372 3584
rect 382366 3544 382372 3556
rect 382424 3544 382430 3596
rect 426066 3544 426072 3596
rect 426124 3584 426130 3596
rect 478690 3584 478696 3596
rect 426124 3556 478696 3584
rect 426124 3544 426130 3556
rect 478690 3544 478696 3556
rect 478748 3544 478754 3596
rect 495158 3544 495164 3596
rect 495216 3584 495222 3596
rect 568761 3587 568819 3593
rect 568761 3584 568773 3587
rect 495216 3556 568773 3584
rect 495216 3544 495222 3556
rect 568761 3553 568773 3556
rect 568807 3553 568819 3587
rect 568761 3547 568819 3553
rect 571426 3544 571432 3596
rect 571484 3584 571490 3596
rect 572622 3584 572628 3596
rect 571484 3556 572628 3584
rect 571484 3544 571490 3556
rect 572622 3544 572628 3556
rect 572680 3544 572686 3596
rect 270586 3516 270592 3528
rect 264532 3488 270592 3516
rect 270586 3476 270592 3488
rect 270644 3476 270650 3528
rect 272886 3476 272892 3528
rect 272944 3516 272950 3528
rect 277394 3516 277400 3528
rect 272944 3488 277400 3516
rect 272944 3476 272950 3488
rect 277394 3476 277400 3488
rect 277452 3476 277458 3528
rect 300762 3476 300768 3528
rect 300820 3516 300826 3528
rect 303798 3516 303804 3528
rect 300820 3488 303804 3516
rect 300820 3476 300826 3488
rect 303798 3476 303804 3488
rect 303856 3476 303862 3528
rect 306190 3476 306196 3528
rect 306248 3516 306254 3528
rect 312170 3516 312176 3528
rect 306248 3488 312176 3516
rect 306248 3476 306254 3488
rect 312170 3476 312176 3488
rect 312228 3476 312234 3528
rect 315942 3476 315948 3528
rect 316000 3516 316006 3528
rect 325234 3516 325240 3528
rect 316000 3488 325240 3516
rect 316000 3476 316006 3488
rect 325234 3476 325240 3488
rect 325292 3476 325298 3528
rect 325510 3476 325516 3528
rect 325568 3516 325574 3528
rect 338298 3516 338304 3528
rect 325568 3488 338304 3516
rect 325568 3476 325574 3488
rect 338298 3476 338304 3488
rect 338356 3476 338362 3528
rect 339402 3476 339408 3528
rect 339460 3516 339466 3528
rect 357342 3516 357348 3528
rect 339460 3488 357348 3516
rect 339460 3476 339466 3488
rect 357342 3476 357348 3488
rect 357400 3476 357406 3528
rect 364242 3476 364248 3528
rect 364300 3516 364306 3528
rect 393038 3516 393044 3528
rect 364300 3488 393044 3516
rect 364300 3476 364306 3488
rect 393038 3476 393044 3488
rect 393096 3476 393102 3528
rect 423582 3476 423588 3528
rect 423640 3516 423646 3528
rect 475102 3516 475108 3528
rect 423640 3488 475108 3516
rect 423640 3476 423646 3488
rect 475102 3476 475108 3488
rect 475160 3476 475166 3528
rect 494054 3476 494060 3528
rect 494112 3516 494118 3528
rect 495342 3516 495348 3528
rect 494112 3488 495348 3516
rect 494112 3476 494118 3488
rect 495342 3476 495348 3488
rect 495400 3476 495406 3528
rect 498102 3476 498108 3528
rect 498160 3516 498166 3528
rect 578602 3516 578608 3528
rect 498160 3488 578608 3516
rect 498160 3476 498166 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 233559 3420 234752 3448
rect 233559 3417 233571 3420
rect 233513 3411 233571 3417
rect 234798 3408 234804 3460
rect 234856 3448 234862 3460
rect 249794 3448 249800 3460
rect 234856 3420 249800 3448
rect 234856 3408 234862 3420
rect 249794 3408 249800 3420
rect 249852 3408 249858 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 265066 3448 265072 3460
rect 255096 3420 265072 3448
rect 255096 3408 255102 3420
rect 265066 3408 265072 3420
rect 265124 3408 265130 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 273346 3448 273352 3460
rect 267056 3420 273352 3448
rect 267056 3408 267062 3420
rect 273346 3408 273352 3420
rect 273404 3408 273410 3460
rect 280062 3408 280068 3460
rect 280120 3448 280126 3460
rect 282914 3448 282920 3460
rect 280120 3420 282920 3448
rect 280120 3408 280126 3420
rect 282914 3408 282920 3420
rect 282972 3408 282978 3460
rect 292482 3408 292488 3460
rect 292540 3448 292546 3460
rect 293126 3448 293132 3460
rect 292540 3420 293132 3448
rect 292540 3408 292546 3420
rect 293126 3408 293132 3420
rect 293184 3408 293190 3460
rect 314470 3408 314476 3460
rect 314528 3448 314534 3460
rect 324038 3448 324044 3460
rect 314528 3420 324044 3448
rect 314528 3408 314534 3420
rect 324038 3408 324044 3420
rect 324096 3408 324102 3460
rect 325602 3408 325608 3460
rect 325660 3448 325666 3460
rect 339494 3448 339500 3460
rect 325660 3420 339500 3448
rect 325660 3408 325666 3420
rect 339494 3408 339500 3420
rect 339552 3408 339558 3460
rect 342162 3408 342168 3460
rect 342220 3448 342226 3460
rect 360930 3448 360936 3460
rect 342220 3420 360936 3448
rect 342220 3408 342226 3420
rect 360930 3408 360936 3420
rect 360988 3408 360994 3460
rect 361482 3408 361488 3460
rect 361540 3448 361546 3460
rect 389450 3448 389456 3460
rect 361540 3420 389456 3448
rect 361540 3408 361546 3420
rect 389450 3408 389456 3420
rect 389508 3408 389514 3460
rect 429102 3408 429108 3460
rect 429160 3448 429166 3460
rect 482278 3448 482284 3460
rect 429160 3420 482284 3448
rect 429160 3408 429166 3420
rect 482278 3408 482284 3420
rect 482336 3408 482342 3460
rect 500862 3408 500868 3460
rect 500920 3448 500926 3460
rect 582190 3448 582196 3460
rect 500920 3420 582196 3448
rect 500920 3408 500926 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 211080 3352 211844 3380
rect 211080 3324 211108 3352
rect 217042 3340 217048 3392
rect 217100 3380 217106 3392
rect 217962 3380 217968 3392
rect 217100 3352 217968 3380
rect 217100 3340 217106 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 224126 3340 224132 3392
rect 224184 3380 224190 3392
rect 241606 3380 241612 3392
rect 224184 3352 241612 3380
rect 224184 3340 224190 3352
rect 241606 3340 241612 3352
rect 241664 3340 241670 3392
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 261018 3380 261024 3392
rect 250404 3352 261024 3380
rect 250404 3340 250410 3352
rect 261018 3340 261024 3352
rect 261076 3340 261082 3392
rect 270494 3340 270500 3392
rect 270552 3380 270558 3392
rect 276106 3380 276112 3392
rect 270552 3352 276112 3380
rect 270552 3340 270558 3352
rect 276106 3340 276112 3352
rect 276164 3340 276170 3392
rect 299290 3340 299296 3392
rect 299348 3380 299354 3392
rect 302602 3380 302608 3392
rect 299348 3352 302608 3380
rect 299348 3340 299354 3352
rect 302602 3340 302608 3352
rect 302660 3340 302666 3392
rect 347685 3383 347743 3389
rect 347685 3349 347697 3383
rect 347731 3380 347743 3383
rect 353754 3380 353760 3392
rect 347731 3352 353760 3380
rect 347731 3349 347743 3352
rect 347685 3343 347743 3349
rect 353754 3340 353760 3352
rect 353812 3340 353818 3392
rect 451274 3340 451280 3392
rect 451332 3380 451338 3392
rect 452470 3380 452476 3392
rect 451332 3352 452476 3380
rect 451332 3340 451338 3352
rect 452470 3340 452476 3352
rect 452528 3340 452534 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 511994 3340 512000 3392
rect 512052 3380 512058 3392
rect 513190 3380 513196 3392
rect 512052 3352 513196 3380
rect 512052 3340 512058 3352
rect 513190 3340 513196 3352
rect 513248 3340 513254 3392
rect 528554 3340 528560 3392
rect 528612 3380 528618 3392
rect 529842 3380 529848 3392
rect 528612 3352 529848 3380
rect 528612 3340 528618 3352
rect 529842 3340 529848 3352
rect 529900 3340 529906 3392
rect 568761 3383 568819 3389
rect 568761 3349 568773 3383
rect 568807 3380 568819 3383
rect 575014 3380 575020 3392
rect 568807 3352 575020 3380
rect 568807 3349 568819 3352
rect 568761 3343 568819 3349
rect 575014 3340 575020 3352
rect 575072 3340 575078 3392
rect 102778 3272 102784 3324
rect 102836 3312 102842 3324
rect 103422 3312 103428 3324
rect 102836 3284 103428 3312
rect 102836 3272 102842 3284
rect 103422 3272 103428 3284
rect 103480 3272 103486 3324
rect 211062 3272 211068 3324
rect 211120 3272 211126 3324
rect 214650 3272 214656 3324
rect 214708 3312 214714 3324
rect 224865 3315 224923 3321
rect 224865 3312 224877 3315
rect 214708 3284 224877 3312
rect 214708 3272 214714 3284
rect 224865 3281 224877 3284
rect 224911 3281 224923 3315
rect 224865 3275 224923 3281
rect 224957 3315 225015 3321
rect 224957 3281 224969 3315
rect 225003 3312 225015 3315
rect 233513 3315 233571 3321
rect 233513 3312 233525 3315
rect 225003 3284 233525 3312
rect 225003 3281 225015 3284
rect 224957 3275 225015 3281
rect 233513 3281 233525 3284
rect 233559 3281 233571 3315
rect 233513 3275 233571 3281
rect 258626 3272 258632 3324
rect 258684 3312 258690 3324
rect 266538 3312 266544 3324
rect 258684 3284 266544 3312
rect 258684 3272 258690 3284
rect 266538 3272 266544 3284
rect 266596 3272 266602 3324
rect 302050 3272 302056 3324
rect 302108 3312 302114 3324
rect 306190 3312 306196 3324
rect 302108 3284 306196 3312
rect 302108 3272 302114 3284
rect 306190 3272 306196 3284
rect 306248 3272 306254 3324
rect 307662 3272 307668 3324
rect 307720 3312 307726 3324
rect 314562 3312 314568 3324
rect 307720 3284 314568 3312
rect 307720 3272 307726 3284
rect 314562 3272 314568 3284
rect 314620 3272 314626 3324
rect 574738 3272 574744 3324
rect 574796 3312 574802 3324
rect 576210 3312 576216 3324
rect 574796 3284 576216 3312
rect 574796 3272 574802 3284
rect 576210 3272 576216 3284
rect 576268 3272 576274 3324
rect 85666 3244 85672 3256
rect 74460 3216 85672 3244
rect 85666 3204 85672 3216
rect 85724 3204 85730 3256
rect 181346 3204 181352 3256
rect 181404 3244 181410 3256
rect 182082 3244 182088 3256
rect 181404 3216 182088 3244
rect 181404 3204 181410 3216
rect 182082 3204 182088 3216
rect 182140 3204 182146 3256
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 19245 3179 19303 3185
rect 19245 3176 19257 3179
rect 9723 3148 19257 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 19245 3145 19257 3148
rect 19291 3145 19303 3179
rect 19245 3139 19303 3145
rect 80238 3136 80244 3188
rect 80296 3176 80302 3188
rect 81342 3176 81348 3188
rect 80296 3148 81348 3176
rect 80296 3136 80302 3148
rect 81342 3136 81348 3148
rect 81400 3136 81406 3188
rect 148042 3136 148048 3188
rect 148100 3176 148106 3188
rect 148962 3176 148968 3188
rect 148100 3148 148968 3176
rect 148100 3136 148106 3148
rect 148962 3136 148968 3148
rect 149020 3136 149026 3188
rect 155126 3136 155132 3188
rect 155184 3176 155190 3188
rect 155862 3176 155868 3188
rect 155184 3148 155868 3176
rect 155184 3136 155190 3148
rect 155862 3136 155868 3148
rect 155920 3136 155926 3188
rect 265802 3136 265808 3188
rect 265860 3176 265866 3188
rect 271969 3179 272027 3185
rect 271969 3176 271981 3179
rect 265860 3148 271981 3176
rect 265860 3136 265866 3148
rect 271969 3145 271981 3148
rect 272015 3145 272027 3179
rect 271969 3139 272027 3145
rect 293862 3136 293868 3188
rect 293920 3176 293926 3188
rect 294322 3176 294328 3188
rect 293920 3148 294328 3176
rect 293920 3136 293926 3148
rect 294322 3136 294328 3148
rect 294380 3136 294386 3188
rect 302142 3136 302148 3188
rect 302200 3176 302206 3188
rect 304994 3176 305000 3188
rect 302200 3148 305000 3176
rect 302200 3136 302206 3148
rect 304994 3136 305000 3148
rect 305052 3136 305058 3188
rect 26694 3068 26700 3120
rect 26752 3108 26758 3120
rect 27522 3108 27528 3120
rect 26752 3080 27528 3108
rect 26752 3068 26758 3080
rect 27522 3068 27528 3080
rect 27580 3068 27586 3120
rect 298002 3068 298008 3120
rect 298060 3108 298066 3120
rect 300302 3108 300308 3120
rect 298060 3080 300308 3108
rect 298060 3068 298066 3080
rect 300302 3068 300308 3080
rect 300360 3068 300366 3120
rect 34974 3000 34980 3052
rect 35032 3040 35038 3052
rect 35802 3040 35808 3052
rect 35032 3012 35808 3040
rect 35032 3000 35038 3012
rect 35802 3000 35808 3012
rect 35860 3000 35866 3052
rect 89714 3000 89720 3052
rect 89772 3040 89778 3052
rect 91002 3040 91008 3052
rect 89772 3012 91008 3040
rect 89772 3000 89778 3012
rect 91002 3000 91008 3012
rect 91060 3000 91066 3052
rect 261018 3000 261024 3052
rect 261076 3040 261082 3052
rect 269114 3040 269120 3052
rect 261076 3012 269120 3040
rect 261076 3000 261082 3012
rect 269114 3000 269120 3012
rect 269172 3000 269178 3052
rect 274082 3000 274088 3052
rect 274140 3040 274146 3052
rect 277578 3040 277584 3052
rect 274140 3012 277584 3040
rect 274140 3000 274146 3012
rect 277578 3000 277584 3012
rect 277636 3000 277642 3052
rect 281258 3000 281264 3052
rect 281316 3040 281322 3052
rect 283098 3040 283104 3052
rect 281316 3012 283104 3040
rect 281316 3000 281322 3012
rect 283098 3000 283104 3012
rect 283156 3000 283162 3052
rect 299382 3000 299388 3052
rect 299440 3040 299446 3052
rect 301406 3040 301412 3052
rect 299440 3012 301412 3040
rect 299440 3000 299446 3012
rect 301406 3000 301412 3012
rect 301464 3000 301470 3052
rect 309042 3000 309048 3052
rect 309100 3040 309106 3052
rect 315758 3040 315764 3052
rect 309100 3012 315764 3040
rect 309100 3000 309106 3012
rect 315758 3000 315764 3012
rect 315816 3000 315822 3052
rect 307570 2932 307576 2984
rect 307628 2972 307634 2984
rect 313366 2972 313372 2984
rect 307628 2944 313372 2972
rect 307628 2932 307634 2944
rect 313366 2932 313372 2944
rect 313424 2932 313430 2984
rect 87322 2864 87328 2916
rect 87380 2904 87386 2916
rect 88242 2904 88248 2916
rect 87380 2876 88248 2904
rect 87380 2864 87386 2876
rect 88242 2864 88248 2876
rect 88300 2864 88306 2916
rect 156322 2864 156328 2916
rect 156380 2904 156386 2916
rect 157242 2904 157248 2916
rect 156380 2876 157248 2904
rect 156380 2864 156386 2876
rect 157242 2864 157248 2876
rect 157300 2864 157306 2916
rect 296530 2864 296536 2916
rect 296588 2904 296594 2916
rect 299106 2904 299112 2916
rect 296588 2876 299112 2904
rect 296588 2864 296594 2876
rect 299106 2864 299112 2876
rect 299164 2864 299170 2916
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 1394 2836 1400 2848
rect 624 2808 1400 2836
rect 624 2796 630 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 14826 2796 14832 2848
rect 14884 2836 14890 2848
rect 15102 2836 15108 2848
rect 14884 2808 15108 2836
rect 14884 2796 14890 2808
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23382 2836 23388 2848
rect 23164 2808 23388 2836
rect 23164 2796 23170 2808
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 40954 2796 40960 2848
rect 41012 2836 41018 2848
rect 41322 2836 41328 2848
rect 41012 2808 41328 2836
rect 41012 2796 41018 2808
rect 41322 2796 41328 2808
rect 41380 2796 41386 2848
rect 83826 2796 83832 2848
rect 83884 2836 83890 2848
rect 84102 2836 84108 2848
rect 83884 2808 84108 2836
rect 83884 2796 83890 2808
rect 84102 2796 84108 2808
rect 84160 2796 84166 2848
rect 177761 2839 177819 2845
rect 177761 2805 177773 2839
rect 177807 2836 177819 2839
rect 177942 2836 177948 2848
rect 177807 2808 177948 2836
rect 177807 2805 177819 2808
rect 177761 2799 177819 2805
rect 177942 2796 177948 2808
rect 178000 2796 178006 2848
rect 310422 2660 310428 2712
rect 310480 2700 310486 2712
rect 316954 2700 316960 2712
rect 310480 2672 316960 2700
rect 310480 2660 310486 2672
rect 316954 2660 316960 2672
rect 317012 2660 317018 2712
rect 206278 1096 206284 1148
rect 206336 1136 206342 1148
rect 206922 1136 206928 1148
rect 206336 1108 206928 1136
rect 206336 1096 206342 1108
rect 206922 1096 206928 1108
rect 206980 1096 206986 1148
rect 31478 592 31484 604
rect 31439 564 31484 592
rect 31478 552 31484 564
rect 31536 552 31542 604
rect 109954 552 109960 604
rect 110012 592 110018 604
rect 110322 592 110328 604
rect 110012 564 110328 592
rect 110012 552 110018 564
rect 110322 552 110328 564
rect 110380 552 110386 604
rect 151538 592 151544 604
rect 151499 564 151544 592
rect 151538 552 151544 564
rect 151596 552 151602 604
rect 161106 552 161112 604
rect 161164 592 161170 604
rect 161382 592 161388 604
rect 161164 564 161388 592
rect 161164 552 161170 564
rect 161382 552 161388 564
rect 161440 552 161446 604
rect 177758 592 177764 604
rect 177719 564 177764 592
rect 177758 552 177764 564
rect 177816 552 177822 604
rect 287146 552 287152 604
rect 287204 592 287210 604
rect 287330 592 287336 604
rect 287204 564 287336 592
rect 287204 552 287210 564
rect 287330 552 287336 564
rect 287388 552 287394 604
rect 351914 552 351920 604
rect 351972 592 351978 604
rect 352558 592 352564 604
rect 351972 564 352564 592
rect 351972 552 351978 564
rect 352558 552 352564 564
rect 352616 552 352622 604
rect 358538 592 358544 604
rect 358499 564 358544 592
rect 358538 552 358544 564
rect 358596 552 358602 604
rect 359734 592 359740 604
rect 359695 564 359740 592
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 406102 592 406108 604
rect 406063 564 406108 592
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 407298 592 407304 604
rect 407259 564 407304 592
rect 407298 552 407304 564
rect 407356 552 407362 604
rect 414474 592 414480 604
rect 414435 564 414480 592
rect 414474 552 414480 564
rect 414532 552 414538 604
rect 431126 592 431132 604
rect 431087 564 431132 592
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 432322 592 432328 604
rect 432283 564 432328 592
rect 432322 552 432328 564
rect 432380 552 432386 604
<< via1 >>
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 364984 699660 365036 699712
rect 365628 699660 365680 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 504364 696940 504416 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 348700 695487 348752 695496
rect 348700 695453 348709 695487
rect 348709 695453 348743 695487
rect 348743 695453 348752 695487
rect 348700 695444 348752 695453
rect 72700 694084 72752 694136
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 412824 692724 412876 692776
rect 542544 692724 542596 692776
rect 542728 692724 542780 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 348792 685856 348844 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 429200 684428 429252 684480
rect 429844 684428 429896 684480
rect 558920 684428 558972 684480
rect 559656 684428 559708 684480
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 412640 683068 412692 683120
rect 429200 683068 429252 683120
rect 542360 683068 542412 683120
rect 558920 683068 558972 683120
rect 3516 681708 3568 681760
rect 8944 681708 8996 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 348700 676175 348752 676184
rect 348700 676141 348709 676175
rect 348709 676141 348743 676175
rect 348743 676141 348752 676175
rect 348700 676132 348752 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 494060 673480 494112 673532
rect 494244 673480 494296 673532
rect 514024 673480 514076 673532
rect 580172 673480 580224 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 219072 666544 219124 666596
rect 348792 666544 348844 666596
rect 413100 666544 413152 666596
rect 429660 666544 429712 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 348884 659608 348936 659660
rect 349068 659608 349120 659660
rect 73068 656820 73120 656872
rect 219348 656820 219400 656872
rect 349068 656820 349120 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 284024 654100 284076 654152
rect 284208 654100 284260 654152
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 14464 652740 14516 652792
rect 525064 650020 525116 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 348976 647275 349028 647284
rect 348976 647241 348985 647275
rect 348985 647241 349019 647275
rect 349019 647241 349028 647275
rect 348976 647232 349028 647241
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 72976 640364 73028 640416
rect 219256 640364 219308 640416
rect 348976 640364 349028 640416
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 72792 640228 72844 640280
rect 219072 640228 219124 640280
rect 348792 640228 348844 640280
rect 72792 637551 72844 637560
rect 72792 637517 72801 637551
rect 72801 637517 72835 637551
rect 72835 637517 72844 637551
rect 72792 637508 72844 637517
rect 219072 637551 219124 637560
rect 219072 637517 219081 637551
rect 219081 637517 219115 637551
rect 219115 637517 219124 637551
rect 219072 637508 219124 637517
rect 348792 637551 348844 637560
rect 348792 637517 348801 637551
rect 348801 637517 348835 637551
rect 348835 637517 348844 637551
rect 348792 637508 348844 637517
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 284024 634788 284076 634840
rect 284208 634788 284260 634840
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 73068 627920 73120 627972
rect 219348 627920 219400 627972
rect 349068 627920 349120 627972
rect 519544 626560 519596 626612
rect 580172 626560 580224 626612
rect 3240 623772 3292 623824
rect 10324 623772 10376 623824
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 284024 615476 284076 615528
rect 284208 615476 284260 615528
rect 477500 615476 477552 615528
rect 477684 615476 477736 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 137744 604120 137796 604172
rect 224132 604120 224184 604172
rect 106188 604052 106240 604104
rect 210608 604052 210660 604104
rect 89628 603984 89680 604036
rect 197084 603984 197136 604036
rect 235908 603984 235960 604036
rect 291844 603984 291896 604036
rect 73068 603916 73120 603968
rect 183468 603916 183520 603968
rect 219348 603916 219400 603968
rect 278320 603916 278372 603968
rect 41328 603848 41380 603900
rect 169944 603848 169996 603900
rect 202788 603848 202840 603900
rect 264796 603848 264848 603900
rect 300768 603848 300820 603900
rect 332508 603848 332560 603900
rect 427360 603848 427412 603900
rect 462320 603848 462372 603900
rect 468024 603848 468076 603900
rect 527180 603848 527232 603900
rect 24768 603780 24820 603832
rect 156420 603780 156472 603832
rect 171048 603780 171100 603832
rect 251272 603780 251324 603832
rect 284024 603780 284076 603832
rect 318984 603780 319036 603832
rect 440884 603780 440936 603832
rect 477684 603780 477736 603832
rect 481548 603780 481600 603832
rect 542452 603780 542504 603832
rect 8024 603712 8076 603764
rect 142896 603712 142948 603764
rect 154304 603712 154356 603764
rect 237656 603712 237708 603764
rect 267648 603712 267700 603764
rect 305460 603712 305512 603764
rect 332324 603712 332376 603764
rect 346032 603712 346084 603764
rect 349068 603712 349120 603764
rect 359648 603712 359700 603764
rect 386696 603712 386748 603764
rect 397460 603712 397512 603764
rect 400220 603712 400272 603764
rect 412732 603712 412784 603764
rect 413836 603712 413888 603764
rect 429292 603712 429344 603764
rect 454408 603712 454460 603764
rect 494244 603712 494296 603764
rect 495072 603712 495124 603764
rect 559012 603712 559064 603764
rect 365628 603236 365680 603288
rect 373172 603236 373224 603288
rect 560944 603100 560996 603152
rect 580172 603100 580224 603152
rect 8944 596096 8996 596148
rect 78680 596096 78732 596148
rect 3332 594804 3384 594856
rect 9036 594804 9088 594856
rect 520924 592016 520976 592068
rect 579896 592016 579948 592068
rect 3424 585080 3476 585132
rect 78680 585080 78732 585132
rect 504364 581612 504416 581664
rect 514024 581612 514076 581664
rect 514024 579640 514076 579692
rect 580172 579640 580224 579692
rect 505008 575424 505060 575476
rect 580264 575424 580316 575476
rect 14464 573996 14516 574048
rect 78680 573996 78732 574048
rect 9036 567808 9088 567860
rect 79324 567808 79376 567860
rect 3424 567196 3476 567248
rect 8944 567196 8996 567248
rect 10324 561620 10376 561672
rect 78680 561620 78732 561672
rect 509884 556180 509936 556232
rect 580172 556180 580224 556232
rect 503812 553324 503864 553376
rect 525064 553324 525116 553376
rect 3516 550536 3568 550588
rect 78680 550536 78732 550588
rect 505744 545096 505796 545148
rect 580172 545096 580224 545148
rect 505008 542308 505060 542360
rect 580356 542308 580408 542360
rect 504364 537480 504416 537532
rect 519544 537480 519596 537532
rect 519544 532720 519596 532772
rect 580172 532720 580224 532772
rect 8944 527076 8996 527128
rect 78680 527076 78732 527128
rect 504640 521568 504692 521620
rect 560944 521568 560996 521620
rect 3424 514700 3476 514752
rect 78680 514700 78732 514752
rect 505008 510552 505060 510604
rect 520924 510552 520976 510604
rect 578240 509600 578292 509652
rect 579988 509600 580040 509652
rect 504364 508512 504416 508564
rect 578240 508512 578292 508564
rect 3516 503616 3568 503668
rect 78680 503616 78732 503668
rect 505008 499468 505060 499520
rect 514024 499468 514076 499520
rect 3424 492600 3476 492652
rect 78680 492600 78732 492652
rect 505008 487432 505060 487484
rect 509884 487432 509936 487484
rect 514024 485800 514076 485852
rect 579896 485800 579948 485852
rect 3516 480156 3568 480208
rect 78680 480156 78732 480208
rect 503720 477232 503772 477284
rect 505744 477232 505796 477284
rect 3424 469140 3476 469192
rect 78680 469140 78732 469192
rect 505008 466352 505060 466404
rect 519544 466352 519596 466404
rect 505744 462340 505796 462392
rect 580172 462340 580224 462392
rect 3424 452548 3476 452600
rect 78680 452548 78732 452600
rect 505008 444320 505060 444372
rect 580264 444320 580316 444372
rect 504364 438880 504416 438932
rect 580172 438880 580224 438932
rect 3148 438812 3200 438864
rect 79324 438812 79376 438864
rect 504640 434664 504692 434716
rect 514024 434664 514076 434716
rect 3240 425008 3292 425060
rect 79324 425008 79376 425060
rect 503720 423444 503772 423496
rect 505744 423444 505796 423496
rect 505008 412564 505060 412616
rect 580356 412564 580408 412616
rect 3148 395972 3200 396024
rect 79416 395972 79468 396024
rect 514024 391960 514076 392012
rect 579896 391960 579948 392012
rect 505008 390464 505060 390516
rect 580448 390464 580500 390516
rect 3240 380808 3292 380860
rect 79508 380808 79560 380860
rect 503904 379448 503956 379500
rect 580264 379448 580316 379500
rect 505008 368432 505060 368484
rect 514024 368432 514076 368484
rect 3148 367004 3200 367056
rect 79324 367004 79376 367056
rect 505008 357348 505060 357400
rect 580264 357348 580316 357400
rect 505008 347692 505060 347744
rect 580356 347692 580408 347744
rect 3424 338036 3476 338088
rect 79416 338036 79468 338088
rect 504548 336676 504600 336728
rect 580264 336676 580316 336728
rect 3240 324232 3292 324284
rect 79692 324232 79744 324284
rect 505008 322872 505060 322924
rect 580172 322872 580224 322924
rect 8944 316004 8996 316056
rect 78680 316004 78732 316056
rect 504088 311788 504140 311840
rect 580172 311788 580224 311840
rect 3332 309068 3384 309120
rect 79324 309068 79376 309120
rect 504548 299412 504600 299464
rect 579804 299412 579856 299464
rect 3424 295264 3476 295316
rect 79600 295264 79652 295316
rect 17224 281528 17276 281580
rect 78680 281528 78732 281580
rect 3424 280100 3476 280152
rect 79508 280100 79560 280152
rect 504364 275952 504416 276004
rect 580172 275952 580224 276004
rect 3148 266296 3200 266348
rect 79416 266296 79468 266348
rect 504456 264868 504508 264920
rect 580172 264868 580224 264920
rect 504364 252492 504416 252544
rect 579804 252492 579856 252544
rect 3240 252424 3292 252476
rect 8944 252424 8996 252476
rect 28264 247052 28316 247104
rect 78680 247052 78732 247104
rect 3424 237328 3476 237380
rect 79324 237328 79376 237380
rect 504548 229032 504600 229084
rect 580172 229032 580224 229084
rect 14464 223592 14516 223644
rect 78680 223592 78732 223644
rect 3148 223524 3200 223576
rect 79600 223524 79652 223576
rect 504456 217948 504508 218000
rect 580172 217948 580224 218000
rect 8944 211148 8996 211200
rect 78680 211148 78732 211200
rect 3424 208292 3476 208344
rect 17224 208292 17276 208344
rect 504364 205572 504416 205624
rect 579804 205572 579856 205624
rect 3148 194488 3200 194540
rect 79508 194488 79560 194540
rect 19984 189048 20036 189100
rect 78680 189048 78732 189100
rect 504640 182112 504692 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 79416 180752 79468 180804
rect 17224 176672 17276 176724
rect 78680 176672 78732 176724
rect 504548 171028 504600 171080
rect 580172 171028 580224 171080
rect 3516 165520 3568 165572
rect 28264 165520 28316 165572
rect 504456 158652 504508 158704
rect 579804 158652 579856 158704
rect 3148 151716 3200 151768
rect 79324 151716 79376 151768
rect 10324 142128 10376 142180
rect 78680 142128 78732 142180
rect 505008 139408 505060 139460
rect 519544 139408 519596 139460
rect 3240 136552 3292 136604
rect 14464 136552 14516 136604
rect 504364 135192 504416 135244
rect 580172 135192 580224 135244
rect 504824 124108 504876 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 8944 122748 8996 122800
rect 504732 111732 504784 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 79692 108944 79744 108996
rect 157984 100648 158036 100700
rect 165988 100648 166040 100700
rect 302516 100648 302568 100700
rect 303528 100648 303580 100700
rect 309416 100648 309468 100700
rect 310428 100648 310480 100700
rect 311900 100648 311952 100700
rect 313096 100648 313148 100700
rect 313648 100648 313700 100700
rect 314568 100648 314620 100700
rect 316224 100648 316276 100700
rect 317236 100648 317288 100700
rect 317880 100648 317932 100700
rect 318708 100648 318760 100700
rect 323032 100648 323084 100700
rect 324228 100648 324280 100700
rect 324780 100648 324832 100700
rect 325516 100648 325568 100700
rect 327264 100648 327316 100700
rect 328368 100648 328420 100700
rect 329012 100648 329064 100700
rect 329748 100648 329800 100700
rect 329840 100648 329892 100700
rect 331036 100648 331088 100700
rect 331588 100648 331640 100700
rect 333244 100648 333296 100700
rect 334164 100648 334216 100700
rect 335268 100648 335320 100700
rect 335820 100648 335872 100700
rect 336556 100648 336608 100700
rect 338396 100648 338448 100700
rect 339408 100648 339460 100700
rect 345204 100648 345256 100700
rect 346216 100648 346268 100700
rect 353760 100648 353812 100700
rect 354588 100648 354640 100700
rect 356336 100648 356388 100700
rect 357348 100648 357400 100700
rect 374276 100648 374328 100700
rect 375196 100648 375248 100700
rect 383660 100648 383712 100700
rect 384948 100648 385000 100700
rect 421196 100648 421248 100700
rect 422208 100648 422260 100700
rect 425428 100648 425480 100700
rect 426256 100648 426308 100700
rect 426348 100648 426400 100700
rect 427084 100648 427136 100700
rect 430580 100648 430632 100700
rect 431868 100648 431920 100700
rect 432328 100648 432380 100700
rect 433984 100648 434036 100700
rect 434904 100648 434956 100700
rect 436008 100648 436060 100700
rect 439136 100648 439188 100700
rect 440148 100648 440200 100700
rect 444288 100648 444340 100700
rect 445024 100648 445076 100700
rect 445944 100648 445996 100700
rect 446956 100648 447008 100700
rect 448520 100648 448572 100700
rect 449716 100648 449768 100700
rect 452752 100648 452804 100700
rect 453856 100648 453908 100700
rect 466460 100648 466512 100700
rect 467748 100648 467800 100700
rect 468116 100648 468168 100700
rect 469864 100648 469916 100700
rect 475016 100648 475068 100700
rect 475936 100648 475988 100700
rect 305092 100580 305144 100632
rect 306288 100580 306340 100632
rect 340972 100580 341024 100632
rect 342168 100580 342220 100632
rect 342628 100580 342680 100632
rect 347044 100580 347096 100632
rect 347780 100580 347832 100632
rect 348976 100580 349028 100632
rect 352012 100580 352064 100632
rect 353208 100580 353260 100632
rect 371700 100580 371752 100632
rect 372528 100580 372580 100632
rect 387892 100580 387944 100632
rect 389088 100580 389140 100632
rect 423772 100580 423824 100632
rect 424968 100580 425020 100632
rect 470692 100580 470744 100632
rect 471888 100580 471940 100632
rect 369952 100512 370004 100564
rect 376024 100512 376076 100564
rect 200764 100376 200816 100428
rect 201776 100376 201828 100428
rect 337568 100104 337620 100156
rect 338764 100104 338816 100156
rect 447692 100104 447744 100156
rect 448428 100104 448480 100156
rect 485228 100104 485280 100156
rect 502984 100104 503036 100156
rect 75184 100036 75236 100088
rect 87420 100036 87472 100088
rect 124864 100036 124916 100088
rect 153200 100036 153252 100088
rect 167644 100036 167696 100088
rect 200948 100036 201000 100088
rect 360568 100036 360620 100088
rect 370504 100036 370556 100088
rect 472440 100036 472492 100088
rect 507124 100036 507176 100088
rect 8944 99968 8996 100020
rect 83188 99968 83240 100020
rect 88248 99968 88300 100020
rect 118976 99968 119028 100020
rect 120724 99968 120776 100020
rect 129280 99968 129332 100020
rect 131764 99968 131816 100020
rect 136916 99968 136968 100020
rect 142804 99968 142856 100020
rect 177028 99968 177080 100020
rect 178684 99968 178736 100020
rect 183928 99968 183980 100020
rect 207664 99968 207716 100020
rect 224040 99968 224092 100020
rect 326436 99968 326488 100020
rect 337384 99968 337436 100020
rect 346952 99968 347004 100020
rect 368572 99968 368624 100020
rect 375932 99968 375984 100020
rect 377404 99968 377456 100020
rect 377680 99968 377732 100020
rect 411352 99968 411404 100020
rect 431408 99968 431460 100020
rect 483664 99968 483716 100020
rect 498016 99968 498068 100020
rect 545764 99968 545816 100020
rect 358912 99832 358964 99884
rect 360108 99832 360160 99884
rect 381084 99832 381136 99884
rect 382188 99832 382240 99884
rect 418620 99764 418672 99816
rect 420184 99764 420236 99816
rect 450268 99764 450320 99816
rect 451924 99764 451976 99816
rect 376852 99628 376904 99680
rect 378048 99628 378100 99680
rect 339224 99492 339276 99544
rect 344284 99492 344336 99544
rect 318800 99424 318852 99476
rect 326344 99424 326396 99476
rect 397276 99424 397328 99476
rect 399484 99424 399536 99476
rect 413560 99424 413612 99476
rect 416044 99424 416096 99476
rect 427176 99424 427228 99476
rect 431224 99424 431276 99476
rect 443368 99424 443420 99476
rect 447784 99424 447836 99476
rect 77944 99356 77996 99408
rect 84016 99356 84068 99408
rect 91744 99356 91796 99408
rect 94228 99356 94280 99408
rect 106924 99356 106976 99408
rect 112168 99356 112220 99408
rect 129004 99356 129056 99408
rect 130108 99356 130160 99408
rect 156604 99356 156656 99408
rect 157432 99356 157484 99408
rect 160100 99356 160152 99408
rect 160836 99356 160888 99408
rect 185584 99356 185636 99408
rect 188160 99356 188212 99408
rect 203524 99356 203576 99408
rect 206100 99356 206152 99408
rect 214564 99356 214616 99408
rect 219716 99356 219768 99408
rect 239404 99356 239456 99408
rect 241980 99356 242032 99408
rect 293132 99356 293184 99408
rect 293868 99356 293920 99408
rect 294052 99356 294104 99408
rect 295156 99356 295208 99408
rect 295708 99356 295760 99408
rect 296628 99356 296680 99408
rect 298284 99356 298336 99408
rect 299388 99356 299440 99408
rect 300860 99356 300912 99408
rect 302148 99356 302200 99408
rect 363144 99356 363196 99408
rect 364156 99356 364208 99408
rect 364892 99356 364944 99408
rect 365628 99356 365680 99408
rect 365720 99356 365772 99408
rect 367008 99356 367060 99408
rect 389640 99356 389692 99408
rect 386144 99288 386196 99340
rect 386328 99288 386380 99340
rect 390468 99356 390520 99408
rect 391204 99356 391256 99408
rect 392216 99356 392268 99408
rect 393136 99356 393188 99408
rect 394700 99356 394752 99408
rect 395896 99356 395948 99408
rect 396448 99356 396500 99408
rect 397368 99356 397420 99408
rect 399024 99356 399076 99408
rect 400036 99356 400088 99408
rect 400680 99356 400732 99408
rect 401508 99356 401560 99408
rect 401600 99356 401652 99408
rect 402796 99356 402848 99408
rect 403256 99356 403308 99408
rect 404176 99356 404228 99408
rect 405832 99356 405884 99408
rect 407028 99356 407080 99408
rect 408408 99356 408460 99408
rect 409144 99356 409196 99408
rect 410064 99356 410116 99408
rect 411168 99356 411220 99408
rect 411812 99356 411864 99408
rect 412548 99356 412600 99408
rect 412640 99356 412692 99408
rect 413928 99356 413980 99408
rect 416964 99356 417016 99408
rect 417976 99356 418028 99408
rect 436560 99356 436612 99408
rect 438124 99356 438176 99408
rect 458732 99356 458784 99408
rect 459468 99356 459520 99408
rect 459652 99356 459704 99408
rect 460848 99356 460900 99408
rect 461308 99356 461360 99408
rect 462228 99356 462280 99408
rect 463884 99356 463936 99408
rect 464896 99356 464948 99408
rect 477500 99356 477552 99408
rect 478788 99356 478840 99408
rect 479248 99356 479300 99408
rect 480168 99356 480220 99408
rect 481824 99356 481876 99408
rect 482928 99356 482980 99408
rect 483480 99356 483532 99408
rect 484308 99356 484360 99408
rect 484400 99356 484452 99408
rect 485688 99356 485740 99408
rect 486056 99356 486108 99408
rect 486976 99356 487028 99408
rect 488632 99356 488684 99408
rect 489736 99356 489788 99408
rect 490380 99356 490432 99408
rect 491944 99356 491996 99408
rect 492864 99356 492916 99408
rect 493876 99356 493928 99408
rect 494612 99356 494664 99408
rect 495348 99356 495400 99408
rect 495440 99356 495492 99408
rect 496636 99356 496688 99408
rect 497188 99356 497240 99408
rect 498108 99356 498160 99408
rect 499764 99356 499816 99408
rect 500868 99356 500920 99408
rect 390468 99220 390520 99272
rect 399852 98676 399904 98728
rect 443000 98676 443052 98728
rect 52368 98608 52420 98660
rect 88248 98608 88300 98660
rect 336648 98608 336700 98660
rect 354680 98608 354732 98660
rect 367468 98608 367520 98660
rect 397460 98608 397512 98660
rect 428004 98608 428056 98660
rect 429108 98608 429160 98660
rect 441712 98608 441764 98660
rect 500960 98608 501012 98660
rect 194600 97928 194652 97980
rect 195612 97928 195664 97980
rect 372620 97316 372672 97368
rect 56508 97248 56560 97300
rect 121552 97248 121604 97300
rect 349528 97248 349580 97300
rect 404360 97248 404412 97300
rect 454500 97248 454552 97300
rect 518900 97248 518952 97300
rect 372620 97180 372672 97232
rect 218336 96840 218388 96892
rect 218888 96840 218940 96892
rect 211436 96704 211488 96756
rect 212080 96704 212132 96756
rect 356888 96636 356940 96688
rect 356980 96636 357032 96688
rect 468760 96636 468812 96688
rect 468852 96636 468904 96688
rect 173164 96568 173216 96620
rect 178408 96568 178460 96620
rect 208676 96568 208728 96620
rect 208860 96568 208912 96620
rect 328184 96568 328236 96620
rect 328276 96568 328328 96620
rect 468852 96543 468904 96552
rect 468852 96509 468861 96543
rect 468861 96509 468895 96543
rect 468895 96509 468904 96543
rect 468852 96500 468904 96509
rect 73068 95888 73120 95940
rect 134340 95888 134392 95940
rect 354496 95888 354548 95940
rect 379520 95888 379572 95940
rect 385316 95888 385368 95940
rect 422300 95888 422352 95940
rect 457076 95888 457128 95940
rect 521660 95888 521712 95940
rect 320456 95276 320508 95328
rect 321468 95276 321520 95328
rect 164424 95208 164476 95260
rect 165160 95208 165212 95260
rect 215576 95208 215628 95260
rect 216312 95208 216364 95260
rect 230848 95208 230900 95260
rect 231676 95208 231728 95260
rect 255872 95208 255924 95260
rect 256424 95208 256476 95260
rect 258356 95208 258408 95260
rect 259000 95208 259052 95260
rect 321192 95208 321244 95260
rect 321376 95208 321428 95260
rect 407580 95208 407632 95260
rect 408224 95208 408276 95260
rect 410892 95208 410944 95260
rect 411076 95208 411128 95260
rect 428832 95208 428884 95260
rect 429016 95208 429068 95260
rect 408224 95115 408276 95124
rect 408224 95081 408233 95115
rect 408233 95081 408267 95115
rect 408267 95081 408276 95115
rect 408224 95072 408276 95081
rect 92480 94528 92532 94580
rect 93124 94528 93176 94580
rect 99380 94528 99432 94580
rect 99932 94528 99984 94580
rect 114560 94528 114612 94580
rect 115204 94528 115256 94580
rect 117320 94528 117372 94580
rect 117780 94528 117832 94580
rect 122840 94528 122892 94580
rect 123852 94528 123904 94580
rect 125600 94528 125652 94580
rect 126428 94528 126480 94580
rect 132500 94528 132552 94580
rect 133236 94528 133288 94580
rect 135260 94528 135312 94580
rect 135812 94528 135864 94580
rect 139400 94528 139452 94580
rect 140044 94528 140096 94580
rect 140780 94528 140832 94580
rect 141700 94528 141752 94580
rect 146300 94528 146352 94580
rect 146852 94528 146904 94580
rect 150440 94528 150492 94580
rect 151084 94528 151136 94580
rect 168380 94528 168432 94580
rect 169116 94528 169168 94580
rect 182180 94528 182232 94580
rect 182732 94528 182784 94580
rect 197360 94528 197412 94580
rect 198004 94528 198056 94580
rect 222200 94528 222252 94580
rect 222844 94528 222896 94580
rect 233332 94528 233384 94580
rect 233884 94528 233936 94580
rect 236092 94528 236144 94580
rect 236460 94528 236512 94580
rect 237380 94528 237432 94580
rect 238116 94528 238168 94580
rect 240140 94528 240192 94580
rect 240692 94528 240744 94580
rect 247040 94528 247092 94580
rect 247684 94528 247736 94580
rect 264980 94528 265032 94580
rect 265532 94528 265584 94580
rect 276020 94528 276072 94580
rect 276572 94528 276624 94580
rect 13728 94460 13780 94512
rect 90824 94460 90876 94512
rect 378508 94460 378560 94512
rect 412640 94460 412692 94512
rect 414388 94460 414440 94512
rect 462320 94460 462372 94512
rect 462412 94460 462464 94512
rect 528560 94460 528612 94512
rect 3424 93780 3476 93832
rect 19984 93780 20036 93832
rect 251548 93780 251600 93832
rect 258356 93780 258408 93832
rect 22008 93100 22060 93152
rect 97172 93100 97224 93152
rect 467656 93100 467708 93152
rect 536840 93100 536892 93152
rect 415032 92463 415084 92472
rect 415032 92429 415041 92463
rect 415041 92429 415075 92463
rect 415075 92429 415084 92463
rect 415032 92420 415084 92429
rect 422116 92463 422168 92472
rect 422116 92429 422125 92463
rect 422125 92429 422159 92463
rect 422159 92429 422168 92463
rect 422116 92420 422168 92429
rect 179420 92352 179472 92404
rect 180156 92352 180208 92404
rect 244280 92352 244332 92404
rect 245108 92352 245160 92404
rect 262220 92352 262272 92404
rect 262956 92352 263008 92404
rect 273260 92352 273312 92404
rect 273996 92352 274048 92404
rect 88248 91740 88300 91792
rect 144092 91740 144144 91792
rect 475936 91740 475988 91792
rect 546592 91740 546644 91792
rect 270500 91536 270552 91588
rect 271420 91536 271472 91588
rect 259460 91264 259512 91316
rect 260380 91264 260432 91316
rect 27528 90312 27580 90364
rect 100852 90312 100904 90364
rect 139308 90312 139360 90364
rect 180800 90312 180852 90364
rect 400036 90312 400088 90364
rect 441620 90312 441672 90364
rect 480076 90312 480128 90364
rect 554780 90312 554832 90364
rect 175556 89768 175608 89820
rect 118792 89700 118844 89752
rect 119528 89700 119580 89752
rect 129740 89700 129792 89752
rect 130384 89700 130436 89752
rect 158904 89700 158956 89752
rect 159640 89700 159692 89752
rect 160100 89700 160152 89752
rect 165712 89700 165764 89752
rect 166356 89700 166408 89752
rect 169944 89700 169996 89752
rect 170404 89700 170456 89752
rect 175464 89700 175516 89752
rect 332324 89700 332376 89752
rect 332508 89700 332560 89752
rect 379244 89700 379296 89752
rect 379428 89700 379480 89752
rect 451004 89700 451056 89752
rect 451188 89700 451240 89752
rect 172888 89675 172940 89684
rect 172888 89641 172897 89675
rect 172897 89641 172931 89675
rect 172931 89641 172940 89675
rect 172888 89632 172940 89641
rect 469036 89632 469088 89684
rect 160192 89564 160244 89616
rect 34428 88952 34480 89004
rect 105544 88952 105596 89004
rect 397368 88952 397420 89004
rect 437480 88952 437532 89004
rect 482836 88952 482888 89004
rect 557540 88952 557592 89004
rect 504640 88272 504692 88324
rect 580172 88272 580224 88324
rect 38568 87592 38620 87644
rect 108304 87592 108356 87644
rect 178132 87091 178184 87100
rect 178132 87057 178141 87091
rect 178141 87057 178175 87091
rect 178175 87057 178184 87091
rect 178132 87048 178184 87057
rect 218336 87116 218388 87168
rect 95608 86980 95660 87032
rect 218244 86980 218296 87032
rect 224868 86980 224920 87032
rect 225328 86980 225380 87032
rect 230848 87023 230900 87032
rect 230848 86989 230857 87023
rect 230857 86989 230891 87023
rect 230891 86989 230900 87023
rect 230848 86980 230900 86989
rect 248880 86980 248932 87032
rect 248972 86980 249024 87032
rect 86132 86955 86184 86964
rect 86132 86921 86141 86955
rect 86141 86921 86175 86955
rect 86175 86921 86184 86955
rect 86132 86912 86184 86921
rect 88524 86955 88576 86964
rect 88524 86921 88533 86955
rect 88533 86921 88567 86955
rect 88567 86921 88576 86955
rect 88524 86912 88576 86921
rect 110604 86912 110656 86964
rect 124312 86912 124364 86964
rect 129924 86912 129976 86964
rect 142252 86912 142304 86964
rect 184020 86955 184072 86964
rect 184020 86921 184029 86955
rect 184029 86921 184063 86955
rect 184063 86921 184072 86955
rect 184020 86912 184072 86921
rect 196072 86912 196124 86964
rect 200304 86955 200356 86964
rect 200304 86921 200313 86955
rect 200313 86921 200347 86955
rect 200347 86921 200356 86955
rect 200304 86912 200356 86921
rect 252744 86912 252796 86964
rect 290096 86912 290148 86964
rect 310152 86955 310204 86964
rect 310152 86921 310161 86955
rect 310161 86921 310195 86955
rect 310195 86921 310204 86955
rect 310152 86912 310204 86921
rect 95700 86844 95752 86896
rect 49608 86232 49660 86284
rect 117412 86232 117464 86284
rect 491944 86232 491996 86284
rect 568580 86232 568632 86284
rect 229284 85552 229336 85604
rect 229652 85552 229704 85604
rect 230848 85595 230900 85604
rect 230848 85561 230857 85595
rect 230857 85561 230891 85595
rect 230891 85561 230900 85595
rect 230848 85552 230900 85561
rect 284576 85552 284628 85604
rect 284760 85552 284812 85604
rect 321192 85552 321244 85604
rect 321284 85552 321336 85604
rect 408224 85595 408276 85604
rect 408224 85561 408233 85595
rect 408233 85561 408267 85595
rect 408267 85561 408276 85595
rect 408224 85552 408276 85561
rect 428832 85552 428884 85604
rect 428924 85552 428976 85604
rect 160192 85527 160244 85536
rect 160192 85493 160201 85527
rect 160201 85493 160235 85527
rect 160235 85493 160244 85527
rect 160192 85484 160244 85493
rect 164424 85527 164476 85536
rect 164424 85493 164433 85527
rect 164433 85493 164467 85527
rect 164467 85493 164476 85527
rect 164424 85484 164476 85493
rect 169944 85527 169996 85536
rect 169944 85493 169953 85527
rect 169953 85493 169987 85527
rect 169987 85493 169996 85527
rect 169944 85484 169996 85493
rect 178132 85527 178184 85536
rect 178132 85493 178141 85527
rect 178141 85493 178175 85527
rect 178175 85493 178184 85527
rect 178132 85484 178184 85493
rect 215484 85484 215536 85536
rect 218244 85484 218296 85536
rect 224868 85527 224920 85536
rect 224868 85493 224877 85527
rect 224877 85493 224911 85527
rect 224911 85493 224920 85527
rect 224868 85484 224920 85493
rect 226524 85527 226576 85536
rect 226524 85493 226533 85527
rect 226533 85493 226567 85527
rect 226567 85493 226576 85527
rect 226524 85484 226576 85493
rect 426072 85484 426124 85536
rect 426164 85484 426216 85536
rect 469036 85484 469088 85536
rect 53748 84804 53800 84856
rect 118792 84804 118844 84856
rect 493876 84804 493928 84856
rect 571432 84804 571484 84856
rect 241612 84192 241664 84244
rect 241796 84192 241848 84244
rect 251456 84235 251508 84244
rect 251456 84201 251465 84235
rect 251465 84201 251499 84235
rect 251499 84201 251508 84235
rect 251456 84192 251508 84201
rect 258264 84235 258316 84244
rect 258264 84201 258273 84235
rect 258273 84201 258307 84235
rect 258307 84201 258316 84235
rect 258264 84192 258316 84201
rect 64788 83444 64840 83496
rect 126980 83444 127032 83496
rect 438768 83444 438820 83496
rect 495440 83444 495492 83496
rect 496636 83444 496688 83496
rect 574744 83444 574796 83496
rect 421932 82900 421984 82952
rect 415032 82875 415084 82884
rect 415032 82841 415041 82875
rect 415041 82841 415075 82875
rect 415075 82841 415084 82875
rect 415032 82832 415084 82841
rect 67548 82084 67600 82136
rect 129004 82084 129056 82136
rect 212724 82084 212776 82136
rect 213092 82084 213144 82136
rect 390192 82084 390244 82136
rect 390376 82084 390428 82136
rect 453856 82084 453908 82136
rect 516140 82084 516192 82136
rect 422024 81379 422076 81388
rect 422024 81345 422033 81379
rect 422033 81345 422067 81379
rect 422067 81345 422076 81379
rect 422024 81336 422076 81345
rect 154948 80724 155000 80776
rect 172888 80724 172940 80776
rect 428648 80724 428700 80776
rect 71688 80656 71740 80708
rect 132592 80656 132644 80708
rect 455328 80656 455380 80708
rect 520280 80656 520332 80708
rect 205732 80180 205784 80232
rect 206468 80180 206520 80232
rect 272156 80180 272208 80232
rect 287428 80180 287480 80232
rect 357072 80180 357124 80232
rect 161756 80112 161808 80164
rect 248880 80155 248932 80164
rect 248880 80121 248889 80155
rect 248889 80121 248923 80155
rect 248923 80121 248932 80155
rect 248880 80112 248932 80121
rect 350264 80112 350316 80164
rect 100760 80044 100812 80096
rect 101496 80044 101548 80096
rect 147680 80044 147732 80096
rect 147864 80044 147916 80096
rect 161664 80044 161716 80096
rect 176660 80044 176712 80096
rect 177120 80044 177172 80096
rect 328000 80044 328052 80096
rect 3424 79976 3476 80028
rect 17224 79976 17276 80028
rect 183744 79976 183796 80028
rect 310244 79976 310296 80028
rect 332508 80044 332560 80096
rect 379336 80112 379388 80164
rect 415032 80044 415084 80096
rect 433064 80044 433116 80096
rect 433248 80044 433300 80096
rect 439872 80044 439924 80096
rect 332416 79976 332468 80028
rect 357072 79976 357124 80028
rect 379336 79976 379388 80028
rect 328092 79908 328144 79960
rect 415124 79908 415176 79960
rect 439964 79908 440016 79960
rect 17868 79296 17920 79348
rect 91744 79296 91796 79348
rect 92388 79296 92440 79348
rect 147772 79296 147824 79348
rect 460756 79296 460808 79348
rect 527180 79296 527232 79348
rect 223672 78548 223724 78600
rect 224132 78548 224184 78600
rect 74448 77936 74500 77988
rect 135352 77936 135404 77988
rect 478696 77936 478748 77988
rect 552020 77936 552072 77988
rect 258264 77324 258316 77376
rect 85856 77256 85908 77308
rect 87236 77256 87288 77308
rect 87604 77256 87656 77308
rect 88524 77299 88576 77308
rect 88524 77265 88533 77299
rect 88533 77265 88567 77299
rect 88567 77265 88576 77299
rect 88524 77256 88576 77265
rect 103612 77256 103664 77308
rect 104072 77256 104124 77308
rect 106280 77256 106332 77308
rect 106648 77256 106700 77308
rect 110512 77299 110564 77308
rect 110512 77265 110521 77299
rect 110521 77265 110555 77299
rect 110555 77265 110564 77299
rect 110512 77256 110564 77265
rect 111800 77256 111852 77308
rect 112076 77256 112128 77308
rect 124220 77299 124272 77308
rect 124220 77265 124229 77299
rect 124229 77265 124263 77299
rect 124263 77265 124272 77299
rect 124220 77256 124272 77265
rect 129832 77299 129884 77308
rect 129832 77265 129841 77299
rect 129841 77265 129875 77299
rect 129875 77265 129884 77299
rect 129832 77256 129884 77265
rect 142160 77299 142212 77308
rect 142160 77265 142169 77299
rect 142169 77265 142203 77299
rect 142203 77265 142212 77299
rect 142160 77256 142212 77265
rect 195980 77299 196032 77308
rect 195980 77265 195989 77299
rect 195989 77265 196023 77299
rect 196023 77265 196032 77299
rect 195980 77256 196032 77265
rect 200304 77299 200356 77308
rect 200304 77265 200313 77299
rect 200313 77265 200347 77299
rect 200347 77265 200356 77299
rect 200304 77256 200356 77265
rect 248604 77256 248656 77308
rect 252652 77299 252704 77308
rect 252652 77265 252661 77299
rect 252661 77265 252695 77299
rect 252695 77265 252704 77299
rect 252652 77256 252704 77265
rect 272064 77299 272116 77308
rect 272064 77265 272073 77299
rect 272073 77265 272107 77299
rect 272107 77265 272116 77299
rect 272064 77256 272116 77265
rect 277584 77256 277636 77308
rect 277676 77256 277728 77308
rect 278872 77256 278924 77308
rect 278964 77256 279016 77308
rect 284576 77324 284628 77376
rect 287336 77299 287388 77308
rect 287336 77265 287345 77299
rect 287345 77265 287379 77299
rect 287379 77265 287388 77299
rect 287336 77256 287388 77265
rect 290004 77299 290056 77308
rect 290004 77265 290013 77299
rect 290013 77265 290047 77299
rect 290047 77265 290056 77299
rect 290004 77256 290056 77265
rect 136732 77231 136784 77240
rect 136732 77197 136741 77231
rect 136741 77197 136775 77231
rect 136775 77197 136784 77231
rect 136732 77188 136784 77197
rect 183744 77231 183796 77240
rect 183744 77197 183753 77231
rect 183753 77197 183787 77231
rect 183787 77197 183796 77231
rect 183744 77188 183796 77197
rect 258264 77188 258316 77240
rect 284392 77188 284444 77240
rect 439964 77231 440016 77240
rect 439964 77197 439973 77231
rect 439973 77197 440007 77231
rect 440007 77197 440016 77231
rect 439964 77188 440016 77197
rect 504548 77188 504600 77240
rect 580172 77188 580224 77240
rect 142160 77163 142212 77172
rect 142160 77129 142169 77163
rect 142169 77129 142203 77163
rect 142203 77129 142212 77163
rect 142160 77120 142212 77129
rect 230848 76644 230900 76696
rect 28908 76508 28960 76560
rect 100760 76508 100812 76560
rect 230848 76508 230900 76560
rect 408132 75964 408184 76016
rect 408224 75964 408276 76016
rect 160192 75939 160244 75948
rect 160192 75905 160201 75939
rect 160201 75905 160235 75939
rect 160235 75905 160244 75939
rect 160192 75896 160244 75905
rect 164424 75939 164476 75948
rect 164424 75905 164433 75939
rect 164433 75905 164467 75939
rect 164467 75905 164476 75939
rect 164424 75896 164476 75905
rect 169944 75939 169996 75948
rect 169944 75905 169953 75939
rect 169953 75905 169987 75939
rect 169987 75905 169996 75939
rect 169944 75896 169996 75905
rect 172612 75939 172664 75948
rect 172612 75905 172621 75939
rect 172621 75905 172655 75939
rect 172655 75905 172664 75939
rect 172612 75896 172664 75905
rect 178408 75896 178460 75948
rect 215392 75939 215444 75948
rect 215392 75905 215401 75939
rect 215401 75905 215435 75939
rect 215435 75905 215444 75939
rect 215392 75896 215444 75905
rect 218152 75939 218204 75948
rect 218152 75905 218161 75939
rect 218161 75905 218195 75939
rect 218195 75905 218204 75939
rect 218152 75896 218204 75905
rect 224960 75896 225012 75948
rect 226616 75896 226668 75948
rect 350172 75939 350224 75948
rect 350172 75905 350181 75939
rect 350181 75905 350215 75939
rect 350215 75905 350224 75939
rect 350172 75896 350224 75905
rect 386144 75896 386196 75948
rect 386328 75896 386380 75948
rect 328092 75828 328144 75880
rect 408132 75871 408184 75880
rect 408132 75837 408141 75871
rect 408141 75837 408175 75871
rect 408175 75837 408184 75871
rect 408132 75828 408184 75837
rect 103612 75148 103664 75200
rect 486976 75148 487028 75200
rect 563152 75148 563204 75200
rect 95792 74468 95844 74520
rect 410892 74511 410944 74520
rect 410892 74477 410901 74511
rect 410901 74477 410935 74511
rect 410935 74477 410944 74511
rect 410892 74468 410944 74477
rect 42708 73788 42760 73840
rect 106924 73788 106976 73840
rect 342076 73788 342128 73840
rect 361580 73788 361632 73840
rect 491208 73788 491260 73840
rect 569960 73788 570012 73840
rect 415124 73108 415176 73160
rect 415400 73108 415452 73160
rect 46848 72428 46900 72480
rect 114652 72428 114704 72480
rect 164424 72428 164476 72480
rect 332416 72428 332468 72480
rect 332600 72428 332652 72480
rect 449716 72428 449768 72480
rect 510620 72428 510672 72480
rect 252468 71544 252520 71596
rect 252652 71544 252704 71596
rect 321192 71068 321244 71120
rect 321376 71068 321428 71120
rect 57888 71000 57940 71052
rect 122932 71000 122984 71052
rect 451004 71000 451056 71052
rect 513380 71000 513432 71052
rect 161664 70456 161716 70508
rect 212724 70499 212776 70508
rect 212724 70465 212733 70499
rect 212733 70465 212767 70499
rect 212767 70465 212776 70499
rect 212724 70456 212776 70465
rect 158812 70388 158864 70440
rect 124220 70320 124272 70372
rect 124404 70320 124456 70372
rect 142252 70320 142304 70372
rect 158904 70252 158956 70304
rect 169944 70388 169996 70440
rect 175464 70388 175516 70440
rect 208492 70388 208544 70440
rect 248604 70431 248656 70440
rect 248604 70397 248613 70431
rect 248613 70397 248647 70431
rect 248647 70397 248656 70431
rect 248604 70388 248656 70397
rect 170036 70252 170088 70304
rect 175556 70252 175608 70304
rect 277584 70388 277636 70440
rect 277492 70320 277544 70372
rect 208584 70252 208636 70304
rect 161664 70184 161716 70236
rect 410984 69980 411036 70032
rect 176844 69844 176896 69896
rect 176844 69708 176896 69760
rect 62028 69640 62080 69692
rect 125692 69640 125744 69692
rect 459468 69640 459520 69692
rect 524420 69640 524472 69692
rect 68928 68280 68980 68332
rect 130016 68280 130068 68332
rect 464896 68280 464948 68332
rect 531320 68280 531372 68332
rect 85764 67779 85816 67788
rect 85764 67745 85773 67779
rect 85773 67745 85807 67779
rect 85807 67745 85816 67779
rect 85764 67736 85816 67745
rect 178132 67668 178184 67720
rect 178408 67668 178460 67720
rect 31668 67643 31720 67652
rect 31668 67609 31677 67643
rect 31677 67609 31711 67643
rect 31711 67609 31720 67643
rect 31668 67600 31720 67609
rect 110512 67600 110564 67652
rect 110604 67600 110656 67652
rect 136824 67600 136876 67652
rect 154764 67643 154816 67652
rect 154764 67609 154773 67643
rect 154773 67609 154807 67643
rect 154807 67609 154816 67643
rect 154764 67600 154816 67609
rect 164332 67643 164384 67652
rect 164332 67609 164341 67643
rect 164341 67609 164375 67643
rect 164375 67609 164384 67643
rect 164332 67600 164384 67609
rect 212724 67643 212776 67652
rect 212724 67609 212733 67643
rect 212733 67609 212767 67643
rect 212767 67609 212776 67643
rect 212724 67600 212776 67609
rect 226616 67668 226668 67720
rect 248604 67643 248656 67652
rect 248604 67609 248613 67643
rect 248613 67609 248647 67643
rect 248647 67609 248656 67643
rect 248604 67600 248656 67609
rect 255412 67600 255464 67652
rect 255504 67600 255556 67652
rect 280344 67600 280396 67652
rect 280436 67600 280488 67652
rect 284392 67600 284444 67652
rect 284484 67600 284536 67652
rect 350172 67600 350224 67652
rect 350356 67600 350408 67652
rect 428924 67600 428976 67652
rect 440056 67600 440108 67652
rect 468944 67643 468996 67652
rect 468944 67609 468953 67643
rect 468953 67609 468987 67643
rect 468987 67609 468996 67643
rect 468944 67600 468996 67609
rect 160192 67575 160244 67584
rect 160192 67541 160201 67575
rect 160201 67541 160235 67575
rect 160235 67541 160244 67575
rect 160192 67532 160244 67541
rect 169852 67532 169904 67584
rect 170036 67532 170088 67584
rect 226524 67532 226576 67584
rect 251364 67532 251416 67584
rect 283104 67575 283156 67584
rect 283104 67541 283113 67575
rect 283113 67541 283147 67575
rect 283147 67541 283156 67575
rect 283104 67532 283156 67541
rect 251456 67464 251508 67516
rect 15108 66852 15160 66904
rect 92572 66852 92624 66904
rect 462228 66852 462280 66904
rect 528652 66852 528704 66904
rect 310060 66376 310112 66428
rect 310244 66376 310296 66428
rect 85764 66283 85816 66292
rect 85764 66249 85773 66283
rect 85773 66249 85807 66283
rect 85807 66249 85816 66283
rect 85764 66240 85816 66249
rect 183744 66283 183796 66292
rect 183744 66249 183753 66283
rect 183753 66249 183787 66283
rect 183787 66249 183796 66283
rect 183744 66240 183796 66249
rect 258172 66240 258224 66292
rect 258264 66240 258316 66292
rect 328000 66283 328052 66292
rect 328000 66249 328009 66283
rect 328009 66249 328043 66283
rect 328043 66249 328052 66283
rect 328000 66240 328052 66249
rect 408224 66240 408276 66292
rect 87144 66215 87196 66224
rect 87144 66181 87153 66215
rect 87153 66181 87187 66215
rect 87187 66181 87196 66215
rect 87144 66172 87196 66181
rect 88432 66172 88484 66224
rect 111800 66172 111852 66224
rect 178132 66172 178184 66224
rect 212724 66215 212776 66224
rect 212724 66181 212733 66215
rect 212733 66181 212767 66215
rect 212767 66181 212776 66215
rect 212724 66172 212776 66181
rect 229284 66172 229336 66224
rect 230664 66172 230716 66224
rect 230756 66172 230808 66224
rect 287336 66172 287388 66224
rect 332324 66215 332376 66224
rect 332324 66181 332333 66215
rect 332333 66181 332367 66215
rect 332367 66181 332376 66215
rect 332324 66172 332376 66181
rect 350356 66172 350408 66224
rect 356980 66215 357032 66224
rect 356980 66181 356989 66215
rect 356989 66181 357023 66215
rect 357023 66181 357032 66215
rect 356980 66172 357032 66181
rect 328000 66147 328052 66156
rect 328000 66113 328009 66147
rect 328009 66113 328043 66147
rect 328043 66113 328052 66147
rect 328000 66104 328052 66113
rect 24768 65492 24820 65544
rect 99472 65492 99524 65544
rect 456708 65492 456760 65544
rect 520372 65492 520424 65544
rect 95516 64923 95568 64932
rect 95516 64889 95525 64923
rect 95525 64889 95559 64923
rect 95559 64889 95568 64923
rect 95516 64880 95568 64889
rect 3332 64812 3384 64864
rect 79600 64812 79652 64864
rect 321100 64855 321152 64864
rect 321100 64821 321109 64855
rect 321109 64821 321143 64855
rect 321143 64821 321152 64855
rect 321100 64812 321152 64821
rect 519544 64812 519596 64864
rect 579804 64812 579856 64864
rect 226524 63928 226576 63980
rect 350356 63860 350408 63912
rect 422024 63563 422076 63572
rect 422024 63529 422033 63563
rect 422033 63529 422067 63563
rect 422067 63529 422076 63563
rect 422024 63520 422076 63529
rect 310060 63452 310112 63504
rect 410984 63452 411036 63504
rect 411076 63452 411128 63504
rect 215392 62772 215444 62824
rect 215576 62772 215628 62824
rect 218152 62772 218204 62824
rect 218336 62772 218388 62824
rect 453948 62772 454000 62824
rect 517520 62772 517572 62824
rect 390008 62092 390060 62144
rect 390100 62092 390152 62144
rect 446956 61344 447008 61396
rect 506480 61344 506532 61396
rect 277492 60868 277544 60920
rect 124404 60843 124456 60852
rect 124404 60809 124413 60843
rect 124413 60809 124447 60843
rect 124447 60809 124456 60843
rect 124404 60800 124456 60809
rect 176844 60800 176896 60852
rect 266636 60800 266688 60852
rect 157524 60732 157576 60784
rect 172796 60732 172848 60784
rect 176752 60732 176804 60784
rect 248696 60732 248748 60784
rect 266544 60732 266596 60784
rect 147864 60664 147916 60716
rect 157340 60664 157392 60716
rect 172888 60664 172940 60716
rect 175372 60664 175424 60716
rect 175556 60664 175608 60716
rect 277584 60664 277636 60716
rect 147956 60596 148008 60648
rect 248696 60596 248748 60648
rect 91008 59984 91060 60036
rect 146392 59984 146444 60036
rect 441528 59984 441580 60036
rect 499580 59984 499632 60036
rect 224868 59848 224920 59900
rect 225052 59848 225104 59900
rect 310244 59211 310296 59220
rect 310244 59177 310253 59211
rect 310253 59177 310287 59211
rect 310287 59177 310296 59211
rect 310244 59168 310296 59177
rect 82728 58624 82780 58676
rect 140872 58624 140924 58676
rect 395896 58624 395948 58676
rect 434720 58624 434772 58676
rect 435916 58624 435968 58676
rect 492680 58624 492732 58676
rect 124312 57944 124364 57996
rect 160192 57987 160244 57996
rect 160192 57953 160201 57987
rect 160201 57953 160235 57987
rect 160235 57953 160244 57987
rect 160192 57944 160244 57953
rect 183744 57944 183796 57996
rect 252468 57944 252520 57996
rect 252652 57944 252704 57996
rect 271972 57944 272024 57996
rect 272064 57944 272116 57996
rect 283104 57987 283156 57996
rect 283104 57953 283113 57987
rect 283113 57953 283147 57987
rect 283147 57953 283156 57987
rect 283104 57944 283156 57953
rect 439872 57944 439924 57996
rect 439964 57944 440016 57996
rect 31668 57919 31720 57928
rect 31668 57885 31677 57919
rect 31677 57885 31711 57919
rect 31711 57885 31720 57919
rect 31668 57876 31720 57885
rect 110696 57919 110748 57928
rect 110696 57885 110705 57919
rect 110705 57885 110739 57919
rect 110739 57885 110748 57919
rect 110696 57876 110748 57885
rect 136916 57876 136968 57928
rect 172888 57919 172940 57928
rect 172888 57885 172897 57919
rect 172897 57885 172931 57919
rect 172931 57885 172940 57919
rect 172888 57876 172940 57885
rect 260840 57919 260892 57928
rect 260840 57885 260849 57919
rect 260849 57885 260883 57919
rect 260883 57885 260892 57919
rect 260840 57876 260892 57885
rect 266544 57876 266596 57928
rect 422300 57876 422352 57928
rect 422392 57876 422444 57928
rect 426256 57919 426308 57928
rect 426256 57885 426265 57919
rect 426265 57885 426299 57919
rect 426299 57885 426308 57919
rect 426256 57876 426308 57885
rect 183744 57808 183796 57860
rect 439872 57851 439924 57860
rect 439872 57817 439881 57851
rect 439881 57817 439915 57851
rect 439915 57817 439924 57851
rect 439872 57808 439924 57817
rect 75828 57196 75880 57248
rect 135260 57196 135312 57248
rect 161388 57196 161440 57248
rect 197452 57196 197504 57248
rect 393136 57196 393188 57248
rect 433248 57196 433300 57248
rect 488540 57196 488592 57248
rect 87144 56627 87196 56636
rect 87144 56593 87153 56627
rect 87153 56593 87187 56627
rect 87187 56593 87196 56627
rect 87144 56584 87196 56593
rect 88340 56627 88392 56636
rect 88340 56593 88349 56627
rect 88349 56593 88383 56627
rect 88383 56593 88392 56627
rect 88340 56584 88392 56593
rect 111892 56627 111944 56636
rect 111892 56593 111901 56627
rect 111901 56593 111935 56627
rect 111935 56593 111944 56627
rect 111892 56584 111944 56593
rect 178408 56627 178460 56636
rect 178408 56593 178417 56627
rect 178417 56593 178451 56627
rect 178451 56593 178460 56627
rect 178408 56584 178460 56593
rect 208492 56584 208544 56636
rect 208676 56584 208728 56636
rect 287244 56627 287296 56636
rect 287244 56593 287253 56627
rect 287253 56593 287287 56627
rect 287287 56593 287296 56627
rect 287244 56584 287296 56593
rect 328000 56627 328052 56636
rect 328000 56593 328009 56627
rect 328009 56593 328043 56627
rect 328043 56593 328052 56627
rect 328000 56584 328052 56593
rect 332416 56584 332468 56636
rect 357072 56584 357124 56636
rect 431960 56584 432012 56636
rect 85764 56559 85816 56568
rect 85764 56525 85773 56559
rect 85773 56525 85807 56559
rect 85807 56525 85816 56559
rect 85764 56516 85816 56525
rect 258172 56491 258224 56500
rect 258172 56457 258181 56491
rect 258181 56457 258215 56491
rect 258215 56457 258224 56491
rect 258172 56448 258224 56457
rect 386144 56015 386196 56024
rect 386144 55981 386153 56015
rect 386153 55981 386187 56015
rect 386187 55981 386196 56015
rect 386144 55972 386196 55981
rect 125508 55836 125560 55888
rect 169852 55836 169904 55888
rect 431868 55836 431920 55888
rect 485780 55836 485832 55888
rect 95332 55224 95384 55276
rect 95424 55224 95476 55276
rect 321192 55224 321244 55276
rect 55128 54476 55180 54528
rect 120080 54476 120132 54528
rect 121368 54476 121420 54528
rect 168472 54476 168524 54528
rect 391204 54476 391256 54528
rect 429200 54476 429252 54528
rect 431224 54476 431276 54528
rect 480260 54476 480312 54528
rect 212816 53796 212868 53848
rect 421932 53796 421984 53848
rect 422024 53796 422076 53848
rect 424876 53116 424928 53168
rect 477592 53116 477644 53168
rect 38476 53048 38528 53100
rect 109040 53048 109092 53100
rect 114468 53048 114520 53100
rect 162860 53048 162912 53100
rect 471796 53048 471848 53100
rect 542360 53048 542412 53100
rect 390192 52436 390244 52488
rect 390284 52436 390336 52488
rect 429016 51824 429068 51876
rect 421932 51756 421984 51808
rect 473360 51756 473412 51808
rect 35808 51688 35860 51740
rect 106464 51688 106516 51740
rect 110328 51688 110380 51740
rect 160192 51688 160244 51740
rect 384856 51688 384908 51740
rect 420920 51688 420972 51740
rect 469128 51688 469180 51740
rect 538220 51688 538272 51740
rect 223672 51144 223724 51196
rect 124312 51119 124364 51128
rect 124312 51085 124321 51119
rect 124321 51085 124355 51119
rect 124355 51085 124364 51119
rect 124312 51076 124364 51085
rect 175556 51076 175608 51128
rect 183744 51076 183796 51128
rect 3424 51008 3476 51060
rect 79508 51008 79560 51060
rect 113180 51008 113232 51060
rect 113364 51008 113416 51060
rect 121460 51008 121512 51060
rect 121644 51008 121696 51060
rect 175372 51008 175424 51060
rect 321192 51076 321244 51128
rect 223672 51008 223724 51060
rect 321100 51008 321152 51060
rect 183744 50940 183796 50992
rect 419448 50396 419500 50448
rect 469220 50396 469272 50448
rect 107568 50328 107620 50380
rect 157340 50328 157392 50380
rect 467748 50328 467800 50380
rect 535460 50328 535512 50380
rect 10416 48968 10468 49020
rect 87144 48968 87196 49020
rect 124128 48968 124180 49020
rect 169760 48968 169812 49020
rect 382096 48968 382148 49020
rect 416780 48968 416832 49020
rect 417976 48968 418028 49020
rect 466460 48968 466512 49020
rect 484308 48968 484360 49020
rect 558920 48968 558972 49020
rect 415400 48900 415452 48952
rect 252652 48424 252704 48476
rect 252560 48356 252612 48408
rect 332416 48356 332468 48408
rect 31668 48331 31720 48340
rect 31668 48297 31677 48331
rect 31677 48297 31711 48331
rect 31711 48297 31720 48331
rect 31668 48288 31720 48297
rect 88340 48288 88392 48340
rect 88432 48288 88484 48340
rect 93952 48288 94004 48340
rect 94044 48288 94096 48340
rect 110788 48288 110840 48340
rect 124312 48331 124364 48340
rect 124312 48297 124321 48331
rect 124321 48297 124355 48331
rect 124355 48297 124364 48331
rect 124312 48288 124364 48297
rect 136824 48331 136876 48340
rect 136824 48297 136833 48331
rect 136833 48297 136867 48331
rect 136867 48297 136876 48331
rect 136824 48288 136876 48297
rect 176660 48288 176712 48340
rect 176936 48288 176988 48340
rect 178132 48288 178184 48340
rect 178408 48288 178460 48340
rect 215484 48288 215536 48340
rect 215576 48288 215628 48340
rect 218244 48288 218296 48340
rect 218336 48288 218388 48340
rect 226616 48331 226668 48340
rect 226616 48297 226625 48331
rect 226625 48297 226659 48331
rect 226659 48297 226668 48331
rect 226616 48288 226668 48297
rect 229376 48331 229428 48340
rect 229376 48297 229385 48331
rect 229385 48297 229419 48331
rect 229419 48297 229428 48331
rect 229376 48288 229428 48297
rect 241704 48288 241756 48340
rect 241796 48288 241848 48340
rect 121644 48263 121696 48272
rect 121644 48229 121653 48263
rect 121653 48229 121687 48263
rect 121687 48229 121696 48263
rect 121644 48220 121696 48229
rect 205732 48220 205784 48272
rect 205824 48220 205876 48272
rect 206928 48220 206980 48272
rect 207112 48220 207164 48272
rect 208584 48220 208636 48272
rect 224960 48220 225012 48272
rect 225052 48220 225104 48272
rect 260840 48331 260892 48340
rect 260840 48297 260849 48331
rect 260849 48297 260883 48331
rect 260883 48297 260892 48331
rect 266452 48331 266504 48340
rect 260840 48288 260892 48297
rect 266452 48297 266461 48331
rect 266461 48297 266495 48331
rect 266495 48297 266504 48331
rect 266452 48288 266504 48297
rect 271972 48288 272024 48340
rect 272064 48288 272116 48340
rect 386328 48288 386380 48340
rect 426348 48288 426400 48340
rect 428832 48331 428884 48340
rect 428832 48297 428841 48331
rect 428841 48297 428875 48331
rect 428875 48297 428884 48331
rect 428832 48288 428884 48297
rect 439964 48288 440016 48340
rect 287244 48263 287296 48272
rect 287244 48229 287253 48263
rect 287253 48229 287287 48263
rect 287287 48229 287296 48263
rect 287244 48220 287296 48229
rect 390284 48220 390336 48272
rect 252560 48152 252612 48204
rect 260840 48195 260892 48204
rect 260840 48161 260849 48195
rect 260849 48161 260883 48195
rect 260883 48161 260892 48195
rect 260840 48152 260892 48161
rect 30288 47540 30340 47592
rect 102140 47540 102192 47592
rect 103428 47540 103480 47592
rect 154764 47540 154816 47592
rect 158628 47540 158680 47592
rect 194692 47540 194744 47592
rect 379244 47540 379296 47592
rect 414020 47540 414072 47592
rect 433984 47540 434036 47592
rect 487160 47540 487212 47592
rect 85764 47039 85816 47048
rect 85764 47005 85773 47039
rect 85773 47005 85807 47039
rect 85807 47005 85816 47039
rect 85764 46996 85816 47005
rect 327908 46996 327960 47048
rect 328000 46996 328052 47048
rect 172612 46928 172664 46980
rect 252468 46971 252520 46980
rect 252468 46937 252477 46971
rect 252477 46937 252511 46971
rect 252511 46937 252520 46971
rect 252468 46928 252520 46937
rect 258172 46971 258224 46980
rect 258172 46937 258181 46971
rect 258181 46937 258215 46971
rect 258215 46937 258224 46971
rect 258172 46928 258224 46937
rect 332324 46971 332376 46980
rect 332324 46937 332333 46971
rect 332333 46937 332367 46971
rect 332367 46937 332376 46971
rect 332324 46928 332376 46937
rect 85764 46860 85816 46912
rect 86040 46860 86092 46912
rect 224960 46903 225012 46912
rect 224960 46869 224969 46903
rect 224969 46869 225003 46903
rect 225003 46869 225012 46903
rect 224960 46860 225012 46869
rect 248972 46903 249024 46912
rect 248972 46869 248981 46903
rect 248981 46869 249015 46903
rect 249015 46869 249024 46903
rect 248972 46860 249024 46869
rect 431960 46903 432012 46912
rect 431960 46869 431969 46903
rect 431969 46869 432003 46903
rect 432003 46869 432012 46903
rect 431960 46860 432012 46869
rect 332324 46792 332376 46844
rect 332416 46792 332468 46844
rect 20628 46180 20680 46232
rect 95424 46180 95476 46232
rect 96528 46180 96580 46232
rect 150532 46180 150584 46232
rect 154488 46180 154540 46232
rect 191840 46180 191892 46232
rect 412548 46180 412600 46232
rect 459652 46180 459704 46232
rect 473268 46180 473320 46232
rect 545120 46180 545172 46232
rect 408132 45568 408184 45620
rect 408316 45568 408368 45620
rect 310060 45500 310112 45552
rect 328000 45500 328052 45552
rect 328092 45500 328144 45552
rect 410984 45500 411036 45552
rect 410984 45364 411036 45416
rect 89628 44820 89680 44872
rect 144920 44820 144972 44872
rect 151728 44820 151780 44872
rect 189080 44820 189132 44872
rect 378048 44820 378100 44872
rect 409880 44820 409932 44872
rect 451924 44820 451976 44872
rect 512000 44820 512052 44872
rect 350356 44208 350408 44260
rect 350540 44208 350592 44260
rect 212816 44115 212868 44124
rect 212816 44081 212825 44115
rect 212825 44081 212859 44115
rect 212859 44081 212868 44115
rect 212816 44072 212868 44081
rect 350356 44115 350408 44124
rect 350356 44081 350365 44115
rect 350365 44081 350399 44115
rect 350399 44081 350408 44115
rect 350356 44072 350408 44081
rect 271972 43460 272024 43512
rect 272248 43460 272300 43512
rect 90916 43392 90968 43444
rect 146300 43392 146352 43444
rect 147588 43392 147640 43444
rect 186412 43392 186464 43444
rect 409788 43392 409840 43444
rect 455420 43392 455472 43444
rect 466368 43392 466420 43444
rect 534080 43392 534132 43444
rect 85488 42032 85540 42084
rect 142344 42032 142396 42084
rect 143448 42032 143500 42084
rect 183744 42032 183796 42084
rect 375196 42032 375248 42084
rect 407120 42032 407172 42084
rect 448428 42032 448480 42084
rect 509240 42032 509292 42084
rect 88432 41420 88484 41472
rect 113364 41420 113416 41472
rect 147956 41463 148008 41472
rect 147956 41429 147965 41463
rect 147965 41429 147999 41463
rect 147999 41429 148008 41463
rect 147956 41420 148008 41429
rect 172612 41420 172664 41472
rect 356980 41420 357032 41472
rect 88340 41352 88392 41404
rect 113364 41284 113416 41336
rect 172704 41284 172756 41336
rect 386328 41420 386380 41472
rect 439964 41420 440016 41472
rect 386236 41352 386288 41404
rect 426164 41352 426216 41404
rect 426348 41352 426400 41404
rect 504456 41352 504508 41404
rect 580172 41352 580224 41404
rect 357072 41284 357124 41336
rect 81348 40672 81400 40724
rect 139492 40672 139544 40724
rect 140688 40672 140740 40724
rect 182272 40672 182324 40724
rect 310244 40715 310296 40724
rect 310244 40681 310253 40715
rect 310253 40681 310287 40715
rect 310287 40681 310296 40715
rect 310244 40672 310296 40681
rect 406936 40672 406988 40724
rect 451280 40672 451332 40724
rect 287244 39831 287296 39840
rect 287244 39797 287253 39831
rect 287253 39797 287287 39831
rect 287287 39797 287296 39831
rect 287244 39788 287296 39797
rect 64696 39312 64748 39364
rect 128452 39312 128504 39364
rect 136548 39312 136600 39364
rect 179512 39312 179564 39364
rect 402796 39312 402848 39364
rect 444380 39312 444432 39364
rect 445668 39312 445720 39364
rect 505100 39312 505152 39364
rect 178224 38768 178276 38820
rect 219624 38768 219676 38820
rect 153384 38700 153436 38752
rect 153476 38700 153528 38752
rect 176936 38700 176988 38752
rect 223672 38700 223724 38752
rect 260840 38743 260892 38752
rect 260840 38709 260849 38743
rect 260849 38709 260883 38743
rect 260883 38709 260892 38743
rect 260840 38700 260892 38709
rect 110696 38632 110748 38684
rect 110788 38632 110840 38684
rect 121736 38632 121788 38684
rect 147956 38675 148008 38684
rect 147956 38641 147965 38675
rect 147965 38641 147999 38675
rect 147999 38641 148008 38675
rect 147956 38632 148008 38641
rect 176844 38632 176896 38684
rect 178224 38632 178276 38684
rect 208492 38675 208544 38684
rect 208492 38641 208501 38675
rect 208501 38641 208535 38675
rect 208535 38641 208544 38675
rect 208492 38632 208544 38641
rect 211344 38632 211396 38684
rect 211528 38632 211580 38684
rect 219624 38632 219676 38684
rect 230756 38632 230808 38684
rect 230848 38632 230900 38684
rect 252468 38632 252520 38684
rect 252652 38632 252704 38684
rect 266452 38632 266504 38684
rect 266544 38632 266596 38684
rect 390192 38675 390244 38684
rect 390192 38641 390201 38675
rect 390201 38641 390235 38675
rect 390235 38641 390244 38675
rect 390192 38632 390244 38641
rect 439872 38675 439924 38684
rect 439872 38641 439881 38675
rect 439881 38641 439915 38675
rect 439915 38641 439924 38675
rect 439872 38632 439924 38641
rect 31668 38607 31720 38616
rect 31668 38573 31677 38607
rect 31677 38573 31711 38607
rect 31711 38573 31720 38607
rect 31668 38564 31720 38573
rect 158812 38607 158864 38616
rect 158812 38573 158821 38607
rect 158821 38573 158855 38607
rect 158855 38573 158864 38607
rect 158812 38564 158864 38573
rect 207020 38607 207072 38616
rect 207020 38573 207029 38607
rect 207029 38573 207063 38607
rect 207063 38573 207072 38607
rect 207020 38564 207072 38573
rect 226616 38607 226668 38616
rect 226616 38573 226625 38607
rect 226625 38573 226659 38607
rect 226659 38573 226668 38607
rect 226616 38564 226668 38573
rect 229376 38607 229428 38616
rect 229376 38573 229385 38607
rect 229385 38573 229419 38607
rect 229419 38573 229428 38607
rect 229376 38564 229428 38573
rect 258172 38564 258224 38616
rect 258264 38564 258316 38616
rect 271788 38564 271840 38616
rect 271972 38564 272024 38616
rect 284484 38607 284536 38616
rect 284484 38573 284493 38607
rect 284493 38573 284527 38607
rect 284527 38573 284536 38607
rect 284484 38564 284536 38573
rect 386236 38607 386288 38616
rect 386236 38573 386245 38607
rect 386245 38573 386279 38607
rect 386279 38573 386288 38607
rect 386236 38564 386288 38573
rect 422300 38564 422352 38616
rect 422392 38564 422444 38616
rect 50988 37884 51040 37936
rect 117320 37884 117372 37936
rect 119988 37884 120040 37936
rect 167000 37884 167052 37936
rect 168288 37884 168340 37936
rect 201592 37884 201644 37936
rect 372528 37884 372580 37936
rect 402980 37884 403032 37936
rect 442816 37884 442868 37936
rect 502340 37884 502392 37936
rect 223580 37315 223632 37324
rect 223580 37281 223589 37315
rect 223589 37281 223623 37315
rect 223623 37281 223632 37315
rect 223580 37272 223632 37281
rect 224960 37315 225012 37324
rect 224960 37281 224969 37315
rect 224969 37281 225003 37315
rect 225003 37281 225012 37315
rect 224960 37272 225012 37281
rect 248972 37315 249024 37324
rect 248972 37281 248981 37315
rect 248981 37281 249015 37315
rect 249015 37281 249024 37315
rect 248972 37272 249024 37281
rect 431960 37315 432012 37324
rect 431960 37281 431969 37315
rect 431969 37281 432003 37315
rect 432003 37281 432012 37315
rect 431960 37272 432012 37281
rect 321192 37204 321244 37256
rect 357072 37247 357124 37256
rect 357072 37213 357081 37247
rect 357081 37213 357115 37247
rect 357115 37213 357124 37247
rect 357072 37204 357124 37213
rect 369768 36592 369820 36644
rect 400220 36592 400272 36644
rect 10968 36524 11020 36576
rect 88340 36524 88392 36576
rect 117228 36524 117280 36576
rect 164332 36524 164384 36576
rect 165528 36524 165580 36576
rect 200304 36524 200356 36576
rect 399484 36524 399536 36576
rect 438860 36524 438912 36576
rect 439872 36524 439924 36576
rect 498200 36524 498252 36576
rect 415308 35955 415360 35964
rect 415308 35921 415317 35955
rect 415317 35921 415351 35955
rect 415351 35921 415360 35955
rect 415308 35912 415360 35921
rect 3424 35844 3476 35896
rect 10324 35844 10376 35896
rect 82636 35164 82688 35216
rect 139400 35164 139452 35216
rect 160008 35164 160060 35216
rect 195980 35164 196032 35216
rect 394608 35164 394660 35216
rect 433340 35164 433392 35216
rect 437388 35164 437440 35216
rect 494060 35164 494112 35216
rect 176752 34663 176804 34672
rect 176752 34629 176761 34663
rect 176761 34629 176795 34663
rect 176795 34629 176804 34663
rect 176752 34620 176804 34629
rect 78588 33736 78640 33788
rect 136916 33736 136968 33788
rect 157248 33736 157300 33788
rect 193312 33736 193364 33788
rect 391848 33736 391900 33788
rect 430580 33736 430632 33788
rect 436008 33736 436060 33788
rect 491300 33736 491352 33788
rect 493968 33736 494020 33788
rect 572720 33736 572772 33788
rect 366916 32444 366968 32496
rect 396080 32444 396132 32496
rect 60648 32376 60700 32428
rect 124220 32376 124272 32428
rect 153108 32376 153160 32428
rect 190552 32376 190604 32428
rect 390192 32376 390244 32428
rect 427820 32376 427872 32428
rect 430488 32376 430540 32428
rect 484400 32376 484452 32428
rect 489736 32376 489788 32428
rect 565820 32376 565872 32428
rect 429016 31875 429068 31884
rect 429016 31841 429025 31875
rect 429025 31841 429059 31875
rect 429059 31841 429068 31875
rect 429016 31832 429068 31841
rect 153476 31807 153528 31816
rect 153476 31773 153485 31807
rect 153485 31773 153519 31807
rect 153519 31773 153528 31807
rect 153476 31764 153528 31773
rect 219624 31764 219676 31816
rect 224960 31764 225012 31816
rect 310244 31764 310296 31816
rect 332416 31764 332468 31816
rect 310152 31696 310204 31748
rect 328092 31696 328144 31748
rect 332324 31696 332376 31748
rect 357072 31739 357124 31748
rect 357072 31705 357081 31739
rect 357081 31705 357115 31739
rect 357115 31705 357124 31739
rect 357072 31696 357124 31705
rect 219716 31628 219768 31680
rect 224960 31628 225012 31680
rect 350356 31671 350408 31680
rect 350356 31637 350365 31671
rect 350365 31637 350399 31671
rect 350399 31637 350408 31671
rect 350356 31628 350408 31637
rect 56416 31016 56468 31068
rect 121736 31016 121788 31068
rect 150348 31016 150400 31068
rect 187792 31016 187844 31068
rect 388996 31016 389048 31068
rect 426440 31016 426492 31068
rect 427084 31016 427136 31068
rect 478880 31016 478932 31068
rect 481548 31016 481600 31068
rect 554872 31016 554924 31068
rect 504364 30268 504416 30320
rect 580172 30268 580224 30320
rect 84108 29588 84160 29640
rect 140780 29588 140832 29640
rect 146208 29588 146260 29640
rect 186320 29588 186372 29640
rect 188988 29588 189040 29640
rect 216680 29588 216732 29640
rect 423680 29588 423732 29640
rect 445024 29588 445076 29640
rect 503720 29588 503772 29640
rect 153384 29044 153436 29096
rect 172704 29044 172756 29096
rect 284484 29087 284536 29096
rect 284484 29053 284493 29087
rect 284493 29053 284527 29087
rect 284527 29053 284536 29087
rect 284484 29044 284536 29053
rect 31668 29019 31720 29028
rect 31668 28985 31677 29019
rect 31677 28985 31711 29019
rect 31711 28985 31720 29019
rect 31668 28976 31720 28985
rect 111800 28976 111852 29028
rect 112076 28976 112128 29028
rect 158996 28976 159048 29028
rect 172612 28976 172664 29028
rect 207112 28976 207164 29028
rect 226616 29019 226668 29028
rect 226616 28985 226625 29019
rect 226625 28985 226659 29019
rect 226659 28985 226668 29019
rect 226616 28976 226668 28985
rect 229376 29019 229428 29028
rect 229376 28985 229385 29019
rect 229385 28985 229419 29019
rect 229419 28985 229428 29019
rect 229376 28976 229428 28985
rect 248696 28976 248748 29028
rect 248972 28976 249024 29028
rect 161664 28951 161716 28960
rect 161664 28917 161673 28951
rect 161673 28917 161707 28951
rect 161707 28917 161716 28951
rect 161664 28908 161716 28917
rect 171140 28951 171192 28960
rect 171140 28917 171149 28951
rect 171149 28917 171183 28951
rect 171183 28917 171192 28951
rect 171140 28908 171192 28917
rect 224960 28951 225012 28960
rect 224960 28917 224969 28951
rect 224969 28917 225003 28951
rect 225003 28917 225012 28951
rect 224960 28908 225012 28917
rect 271972 28951 272024 28960
rect 271972 28917 271981 28951
rect 271981 28917 272015 28951
rect 272015 28917 272024 28951
rect 271972 28908 272024 28917
rect 284484 28951 284536 28960
rect 284484 28917 284493 28951
rect 284493 28917 284527 28951
rect 284527 28917 284536 28951
rect 284484 28908 284536 28917
rect 287244 28951 287296 28960
rect 287244 28917 287253 28951
rect 287253 28917 287287 28951
rect 287287 28917 287296 28951
rect 287244 28908 287296 28917
rect 212816 28883 212868 28892
rect 212816 28849 212825 28883
rect 212825 28849 212859 28883
rect 212859 28849 212868 28883
rect 212816 28840 212868 28849
rect 424968 28296 425020 28348
rect 476120 28296 476172 28348
rect 45468 28228 45520 28280
rect 113364 28228 113416 28280
rect 142068 28228 142120 28280
rect 178684 28228 178736 28280
rect 182088 28228 182140 28280
rect 211344 28228 211396 28280
rect 384948 28228 385000 28280
rect 419540 28228 419592 28280
rect 476028 28228 476080 28280
rect 547880 28228 547932 28280
rect 429016 27727 429068 27736
rect 429016 27693 429025 27727
rect 429025 27693 429059 27727
rect 429059 27693 429068 27727
rect 429016 27684 429068 27693
rect 176936 27616 176988 27668
rect 321100 27659 321152 27668
rect 321100 27625 321109 27659
rect 321109 27625 321143 27659
rect 321143 27625 321152 27659
rect 321100 27616 321152 27625
rect 153292 27591 153344 27600
rect 153292 27557 153301 27591
rect 153301 27557 153335 27591
rect 153335 27557 153344 27591
rect 153292 27548 153344 27557
rect 255412 27591 255464 27600
rect 255412 27557 255421 27591
rect 255421 27557 255455 27591
rect 255455 27557 255464 27591
rect 255412 27548 255464 27557
rect 357164 27591 357216 27600
rect 357164 27557 357173 27591
rect 357173 27557 357207 27591
rect 357207 27557 357216 27591
rect 357164 27548 357216 27557
rect 408224 27591 408276 27600
rect 408224 27557 408233 27591
rect 408233 27557 408267 27591
rect 408267 27557 408276 27591
rect 408224 27548 408276 27557
rect 422300 27591 422352 27600
rect 422300 27557 422309 27591
rect 422309 27557 422343 27591
rect 422343 27557 422352 27591
rect 422300 27548 422352 27557
rect 428740 27548 428792 27600
rect 429016 27548 429068 27600
rect 431960 27591 432012 27600
rect 431960 27557 431969 27591
rect 431969 27557 432003 27591
rect 432003 27557 432012 27591
rect 431960 27548 432012 27557
rect 310060 27480 310112 27532
rect 70308 26868 70360 26920
rect 131120 26868 131172 26920
rect 132408 26868 132460 26920
rect 175464 26868 175516 26920
rect 177948 26868 178000 26920
rect 208492 26868 208544 26920
rect 382188 26868 382240 26920
rect 416872 26868 416924 26920
rect 422208 26868 422260 26920
rect 471980 26868 472032 26920
rect 488448 26868 488500 26920
rect 564440 26868 564492 26920
rect 327908 26367 327960 26376
rect 327908 26333 327917 26367
rect 327917 26333 327951 26367
rect 327951 26333 327960 26367
rect 327908 26324 327960 26333
rect 212816 26188 212868 26240
rect 327908 26188 327960 26240
rect 41328 25508 41380 25560
rect 110696 25508 110748 25560
rect 129648 25508 129700 25560
rect 173900 25508 173952 25560
rect 175188 25508 175240 25560
rect 205732 25508 205784 25560
rect 373908 25508 373960 25560
rect 405740 25508 405792 25560
rect 420184 25508 420236 25560
rect 467932 25508 467984 25560
rect 471888 25508 471940 25560
rect 540980 25508 541032 25560
rect 23388 24080 23440 24132
rect 98000 24080 98052 24132
rect 106188 24080 106240 24132
rect 156604 24080 156656 24132
rect 168196 24080 168248 24132
rect 200764 24080 200816 24132
rect 202696 24080 202748 24132
rect 226616 24080 226668 24132
rect 368296 24080 368348 24132
rect 398840 24080 398892 24132
rect 416688 24080 416740 24132
rect 465080 24080 465132 24132
rect 470508 24080 470560 24132
rect 539600 24080 539652 24132
rect 30196 22720 30248 22772
rect 103520 22720 103572 22772
rect 108948 22720 109000 22772
rect 159088 22720 159140 22772
rect 164148 22720 164200 22772
rect 198740 22720 198792 22772
rect 200028 22720 200080 22772
rect 223580 22720 223632 22772
rect 353116 22720 353168 22772
rect 376760 22720 376812 22772
rect 377404 22720 377456 22772
rect 408500 22720 408552 22772
rect 416044 22720 416096 22772
rect 460940 22720 460992 22772
rect 469864 22720 469916 22772
rect 536932 22720 536984 22772
rect 254124 22244 254176 22296
rect 229376 22219 229428 22228
rect 229376 22185 229385 22219
rect 229385 22185 229419 22219
rect 229419 22185 229428 22219
rect 229376 22176 229428 22185
rect 85948 22108 86000 22160
rect 165804 22108 165856 22160
rect 176936 22108 176988 22160
rect 230756 22108 230808 22160
rect 254124 22108 254176 22160
rect 321100 22151 321152 22160
rect 321100 22117 321109 22151
rect 321109 22117 321143 22151
rect 321143 22117 321152 22151
rect 321100 22108 321152 22117
rect 332324 22108 332376 22160
rect 3148 22040 3200 22092
rect 79416 22040 79468 22092
rect 85764 22040 85816 22092
rect 111892 22040 111944 22092
rect 112076 22040 112128 22092
rect 165712 22040 165764 22092
rect 176752 22040 176804 22092
rect 332324 21972 332376 22024
rect 328092 21947 328144 21956
rect 328092 21913 328101 21947
rect 328101 21913 328135 21947
rect 328135 21913 328144 21947
rect 328092 21904 328144 21913
rect 128268 21428 128320 21480
rect 172612 21428 172664 21480
rect 86868 21360 86920 21412
rect 143540 21360 143592 21412
rect 171048 21360 171100 21412
rect 204352 21360 204404 21412
rect 206928 21360 206980 21412
rect 348976 21360 349028 21412
rect 369860 21360 369912 21412
rect 371148 21360 371200 21412
rect 401600 21360 401652 21412
rect 410984 21360 411036 21412
rect 458180 21360 458232 21412
rect 463608 21360 463660 21412
rect 529940 21360 529992 21412
rect 19248 19932 19300 19984
rect 94136 19932 94188 19984
rect 102048 19932 102100 19984
rect 154580 19932 154632 19984
rect 159916 19932 159968 19984
rect 194600 19932 194652 19984
rect 195888 19932 195940 19984
rect 222292 19932 222344 19984
rect 370504 19932 370556 19984
rect 387800 19932 387852 19984
rect 409144 19932 409196 19984
rect 454040 19932 454092 19984
rect 458088 19932 458140 19984
rect 523040 19932 523092 19984
rect 224960 19431 225012 19440
rect 224960 19397 224969 19431
rect 224969 19397 225003 19431
rect 225003 19397 225012 19431
rect 224960 19388 225012 19397
rect 161848 19320 161900 19372
rect 171324 19320 171376 19372
rect 207020 19320 207072 19372
rect 207112 19320 207164 19372
rect 230664 19363 230716 19372
rect 230664 19329 230673 19363
rect 230673 19329 230707 19363
rect 230707 19329 230716 19363
rect 230664 19320 230716 19329
rect 271972 19363 272024 19372
rect 271972 19329 271981 19363
rect 271981 19329 272015 19363
rect 272015 19329 272024 19363
rect 271972 19320 272024 19329
rect 284484 19363 284536 19372
rect 284484 19329 284493 19363
rect 284493 19329 284527 19363
rect 284527 19329 284536 19363
rect 284484 19320 284536 19329
rect 287336 19320 287388 19372
rect 31484 19252 31536 19304
rect 31668 19252 31720 19304
rect 112076 19295 112128 19304
rect 112076 19261 112085 19295
rect 112085 19261 112119 19295
rect 112119 19261 112128 19295
rect 112076 19252 112128 19261
rect 212908 19295 212960 19304
rect 212908 19261 212917 19295
rect 212917 19261 212951 19295
rect 212951 19261 212960 19295
rect 212908 19252 212960 19261
rect 224960 19295 225012 19304
rect 224960 19261 224969 19295
rect 224969 19261 225003 19295
rect 225003 19261 225012 19295
rect 224960 19252 225012 19261
rect 248604 19295 248656 19304
rect 248604 19261 248613 19295
rect 248613 19261 248647 19295
rect 248647 19261 248656 19295
rect 248604 19252 248656 19261
rect 260840 19295 260892 19304
rect 260840 19261 260849 19295
rect 260849 19261 260883 19295
rect 260883 19261 260892 19295
rect 260840 19252 260892 19261
rect 193128 18640 193180 18692
rect 214564 18640 214616 18692
rect 13636 18572 13688 18624
rect 91100 18572 91152 18624
rect 99196 18572 99248 18624
rect 151820 18572 151872 18624
rect 155868 18572 155920 18624
rect 193220 18572 193272 18624
rect 217968 18572 218020 18624
rect 237472 18572 237524 18624
rect 346216 18572 346268 18624
rect 365720 18572 365772 18624
rect 367008 18572 367060 18624
rect 407028 18572 407080 18624
rect 451372 18572 451424 18624
rect 478788 18572 478840 18624
rect 550640 18572 550692 18624
rect 153384 17960 153436 18012
rect 255412 18003 255464 18012
rect 255412 17969 255421 18003
rect 255421 17969 255455 18003
rect 255455 17969 255464 18003
rect 255412 17960 255464 17969
rect 321100 18003 321152 18012
rect 321100 17969 321109 18003
rect 321109 17969 321143 18003
rect 321143 17969 321152 18003
rect 321100 17960 321152 17969
rect 357256 17960 357308 18012
rect 408408 17960 408460 18012
rect 431960 18003 432012 18012
rect 431960 17969 431969 18003
rect 431969 17969 432003 18003
rect 432003 17969 432012 18003
rect 431960 17960 432012 17969
rect 505744 17892 505796 17944
rect 579804 17892 579856 17944
rect 184848 17280 184900 17332
rect 213920 17280 213972 17332
rect 9036 17212 9088 17264
rect 84200 17212 84252 17264
rect 95148 17212 95200 17264
rect 149060 17212 149112 17264
rect 151636 17212 151688 17264
rect 190460 17212 190512 17264
rect 234620 17212 234672 17264
rect 340788 17212 340840 17264
rect 358820 17212 358872 17264
rect 364156 17212 364208 17264
rect 390560 17212 390612 17264
rect 404176 17212 404228 17264
rect 447140 17212 447192 17264
rect 447784 17212 447836 17264
rect 502432 17212 502484 17264
rect 408408 16847 408460 16856
rect 408408 16813 408417 16847
rect 408417 16813 408451 16847
rect 408451 16813 408460 16847
rect 408408 16804 408460 16813
rect 350264 16600 350316 16652
rect 350356 16600 350408 16652
rect 77208 15852 77260 15904
rect 131764 15852 131816 15904
rect 148968 15852 149020 15904
rect 185584 15852 185636 15904
rect 198648 15852 198700 15904
rect 207664 15852 207716 15904
rect 211068 15852 211120 15904
rect 231860 15852 231912 15904
rect 335176 15852 335228 15904
rect 351920 15852 351972 15904
rect 355968 15852 356020 15904
rect 380900 15852 380952 15904
rect 401508 15852 401560 15904
rect 443092 15852 443144 15904
rect 464988 15852 465040 15904
rect 532700 15852 532752 15904
rect 117136 14492 117188 14544
rect 157984 14492 158036 14544
rect 66168 14424 66220 14476
rect 120724 14424 120776 14476
rect 144828 14424 144880 14476
rect 184940 14424 184992 14476
rect 191748 14424 191800 14476
rect 218244 14424 218296 14476
rect 240232 14424 240284 14476
rect 344284 14424 344336 14476
rect 357440 14424 357492 14476
rect 358728 14424 358780 14476
rect 383660 14424 383712 14476
rect 398748 14424 398800 14476
rect 440240 14424 440292 14476
rect 460848 14424 460900 14476
rect 525800 14424 525852 14476
rect 375288 13132 375340 13184
rect 408592 13132 408644 13184
rect 63408 13064 63460 13116
rect 125600 13064 125652 13116
rect 141976 13064 142028 13116
rect 182180 13064 182232 13116
rect 187608 13064 187660 13116
rect 215484 13064 215536 13116
rect 219348 13064 219400 13116
rect 238760 13064 238812 13116
rect 332324 13064 332376 13116
rect 347780 13064 347832 13116
rect 350264 13064 350316 13116
rect 374092 13064 374144 13116
rect 404268 13064 404320 13116
rect 448520 13064 448572 13116
rect 452568 13064 452620 13116
rect 514760 13064 514812 13116
rect 176752 12495 176804 12504
rect 176752 12461 176761 12495
rect 176761 12461 176795 12495
rect 176795 12461 176804 12495
rect 176752 12452 176804 12461
rect 251364 12452 251416 12504
rect 398840 12452 398892 12504
rect 402980 12452 403032 12504
rect 251272 12384 251324 12436
rect 396080 12384 396132 12436
rect 396632 12384 396684 12436
rect 310336 12316 310388 12368
rect 397552 12316 397604 12368
rect 397828 12316 397880 12368
rect 401600 12384 401652 12436
rect 402520 12384 402572 12436
rect 399024 12316 399076 12368
rect 404360 12384 404412 12436
rect 404912 12384 404964 12436
rect 409880 12384 409932 12436
rect 410892 12384 410944 12436
rect 411352 12384 411404 12436
rect 412088 12384 412140 12436
rect 412640 12384 412692 12436
rect 413284 12384 413336 12436
rect 414020 12384 414072 12436
rect 414480 12384 414532 12436
rect 419540 12384 419592 12436
rect 420368 12384 420420 12436
rect 420920 12384 420972 12436
rect 421564 12384 421616 12436
rect 426440 12384 426492 12436
rect 427544 12384 427596 12436
rect 427820 12384 427872 12436
rect 428740 12384 428792 12436
rect 429200 12384 429252 12436
rect 429936 12384 429988 12436
rect 430580 12384 430632 12436
rect 431132 12384 431184 12436
rect 434720 12384 434772 12436
rect 435824 12384 435876 12436
rect 403716 12316 403768 12368
rect 112076 11883 112128 11892
rect 112076 11849 112085 11883
rect 112085 11849 112119 11883
rect 112119 11849 112128 11883
rect 112076 11840 112128 11849
rect 59268 11704 59320 11756
rect 122840 11704 122892 11756
rect 137928 11704 137980 11756
rect 179420 11704 179472 11756
rect 183744 11704 183796 11756
rect 212908 11704 212960 11756
rect 215852 11704 215904 11756
rect 236092 11704 236144 11756
rect 331036 11704 331088 11756
rect 345020 11704 345072 11756
rect 347044 11704 347096 11756
rect 362960 11704 363012 11756
rect 365628 11704 365680 11756
rect 394240 11704 394292 11756
rect 395988 11704 396040 11756
rect 437020 11704 437072 11756
rect 449808 11704 449860 11756
rect 512092 11704 512144 11756
rect 48228 10276 48280 10328
rect 115940 10276 115992 10328
rect 133788 10276 133840 10328
rect 180156 10276 180208 10328
rect 211160 10276 211212 10328
rect 212264 10276 212316 10328
rect 233332 10276 233384 10328
rect 233700 10276 233752 10328
rect 329748 10276 329800 10328
rect 343640 10276 343692 10328
rect 362868 10276 362920 10328
rect 390652 10276 390704 10328
rect 393228 10276 393280 10328
rect 433524 10276 433576 10328
rect 447048 10276 447100 10328
rect 507860 10276 507912 10328
rect 328092 9732 328144 9784
rect 213460 9707 213512 9716
rect 213460 9673 213469 9707
rect 213469 9673 213503 9707
rect 213503 9673 213512 9707
rect 213460 9664 213512 9673
rect 220544 9707 220596 9716
rect 220544 9673 220553 9707
rect 220553 9673 220587 9707
rect 220587 9673 220596 9707
rect 220544 9664 220596 9673
rect 225052 9664 225104 9716
rect 261024 9664 261076 9716
rect 395436 9707 395488 9716
rect 395436 9673 395445 9707
rect 395445 9673 395479 9707
rect 395479 9673 395488 9707
rect 395436 9664 395488 9673
rect 408408 9707 408460 9716
rect 408408 9673 408417 9707
rect 408417 9673 408451 9707
rect 408451 9673 408460 9707
rect 408408 9664 408460 9673
rect 422760 9664 422812 9716
rect 31668 9596 31720 9648
rect 85764 9639 85816 9648
rect 85764 9605 85773 9639
rect 85773 9605 85807 9639
rect 85807 9605 85816 9639
rect 85764 9596 85816 9605
rect 151636 9596 151688 9648
rect 271972 9639 272024 9648
rect 271972 9605 271981 9639
rect 271981 9605 272015 9639
rect 272015 9605 272024 9639
rect 271972 9596 272024 9605
rect 283656 9596 283708 9648
rect 284484 9596 284536 9648
rect 328092 9596 328144 9648
rect 357440 9596 357492 9648
rect 358820 9596 358872 9648
rect 397828 9596 397880 9648
rect 399024 9596 399076 9648
rect 403716 9596 403768 9648
rect 406108 9639 406160 9648
rect 406108 9605 406117 9639
rect 406117 9605 406151 9639
rect 406151 9605 406160 9639
rect 406108 9596 406160 9605
rect 407304 9639 407356 9648
rect 407304 9605 407313 9639
rect 407313 9605 407347 9639
rect 407347 9605 407356 9639
rect 407304 9596 407356 9605
rect 414480 9639 414532 9648
rect 414480 9605 414489 9639
rect 414489 9605 414523 9639
rect 414523 9605 414532 9639
rect 414480 9596 414532 9605
rect 428924 9639 428976 9648
rect 428924 9605 428933 9639
rect 428933 9605 428967 9639
rect 428967 9605 428976 9639
rect 428924 9596 428976 9605
rect 431132 9639 431184 9648
rect 431132 9605 431141 9639
rect 431141 9605 431175 9639
rect 431175 9605 431184 9639
rect 431132 9596 431184 9605
rect 432328 9639 432380 9648
rect 432328 9605 432337 9639
rect 432337 9605 432371 9639
rect 432371 9605 432380 9639
rect 432328 9596 432380 9605
rect 321100 9571 321152 9580
rect 321100 9537 321109 9571
rect 321109 9537 321143 9571
rect 321143 9537 321152 9571
rect 321100 9528 321152 9537
rect 397828 9460 397880 9512
rect 399024 9460 399076 9512
rect 403716 9460 403768 9512
rect 130200 8984 130252 9036
rect 175280 8984 175332 9036
rect 2872 8916 2924 8968
rect 77944 8916 77996 8968
rect 79048 8916 79100 8968
rect 138020 8916 138072 8968
rect 176568 8916 176620 8968
rect 208400 8916 208452 8968
rect 208676 8916 208728 8968
rect 230756 8916 230808 8968
rect 237196 8916 237248 8968
rect 251272 8916 251324 8968
rect 338764 8916 338816 8968
rect 356152 8916 356204 8968
rect 360016 8916 360068 8968
rect 387064 8916 387116 8968
rect 389088 8916 389140 8968
rect 426348 8916 426400 8968
rect 440148 8916 440200 8968
rect 497740 8916 497792 8968
rect 499488 8916 499540 8968
rect 581000 8916 581052 8968
rect 337384 8508 337436 8560
rect 340696 8508 340748 8560
rect 4068 8236 4120 8288
rect 79324 8236 79376 8288
rect 169392 7624 169444 7676
rect 202880 7624 202932 7676
rect 390560 7624 390612 7676
rect 391848 7624 391900 7676
rect 408500 7624 408552 7676
rect 409696 7624 409748 7676
rect 71872 7556 71924 7608
rect 132500 7556 132552 7608
rect 134892 7556 134944 7608
rect 178224 7556 178276 7608
rect 205088 7556 205140 7608
rect 229100 7556 229152 7608
rect 230112 7556 230164 7608
rect 247132 7556 247184 7608
rect 324136 7556 324188 7608
rect 337108 7556 337160 7608
rect 344928 7556 344980 7608
rect 365812 7556 365864 7608
rect 380808 7556 380860 7608
rect 415676 7556 415728 7608
rect 416780 7556 416832 7608
rect 417976 7556 418028 7608
rect 438124 7556 438176 7608
rect 494152 7556 494204 7608
rect 496728 7556 496780 7608
rect 577412 7556 577464 7608
rect 132592 6196 132644 6248
rect 142804 6196 142856 6248
rect 194416 6196 194468 6248
rect 220820 6196 220872 6248
rect 7656 6128 7708 6180
rect 75184 6128 75236 6180
rect 112352 6128 112404 6180
rect 161848 6128 161900 6180
rect 162308 6128 162360 6180
rect 197360 6128 197412 6180
rect 222936 6128 222988 6180
rect 239404 6128 239456 6180
rect 240784 6128 240836 6180
rect 254124 6128 254176 6180
rect 333244 6128 333296 6180
rect 347872 6128 347924 6180
rect 357164 6128 357216 6180
rect 383476 6128 383528 6180
rect 383568 6128 383620 6180
rect 419172 6128 419224 6180
rect 434628 6128 434680 6180
rect 490564 6128 490616 6180
rect 502984 6128 503036 6180
rect 561956 6128 562008 6180
rect 333612 5992 333664 6044
rect 433340 5992 433392 6044
rect 434628 5992 434680 6044
rect 1676 5516 1728 5568
rect 8944 5516 8996 5568
rect 326344 5448 326396 5500
rect 330024 5448 330076 5500
rect 165896 4836 165948 4888
rect 167644 4836 167696 4888
rect 201500 4836 201552 4888
rect 226340 4836 226392 4888
rect 310244 4836 310296 4888
rect 318064 4836 318116 4888
rect 376024 4836 376076 4888
rect 401324 4836 401376 4888
rect 1400 4768 1452 4820
rect 81440 4768 81492 4820
rect 99288 4768 99340 4820
rect 124864 4768 124916 4820
rect 126612 4768 126664 4820
rect 172520 4768 172572 4820
rect 172980 4768 173032 4820
rect 203524 4768 203576 4820
rect 226524 4768 226576 4820
rect 244372 4768 244424 4820
rect 244464 4768 244516 4820
rect 256700 4768 256752 4820
rect 335268 4768 335320 4820
rect 351368 4768 351420 4820
rect 353208 4768 353260 4820
rect 376392 4768 376444 4820
rect 387708 4768 387760 4820
rect 425152 4768 425204 4820
rect 483480 4768 483532 4820
rect 507124 4768 507176 4820
rect 544108 4768 544160 4820
rect 545764 4768 545816 4820
rect 579804 4768 579856 4820
rect 317236 4700 317288 4752
rect 326436 4700 326488 4752
rect 483664 4156 483716 4208
rect 486976 4156 487028 4208
rect 502432 4156 502484 4208
rect 503628 4156 503680 4208
rect 536932 4156 536984 4208
rect 538128 4156 538180 4208
rect 8852 4088 8904 4140
rect 10416 4088 10468 4140
rect 12440 4088 12492 4140
rect 13728 4088 13780 4140
rect 17224 4088 17276 4140
rect 17868 4088 17920 4140
rect 18328 4088 18380 4140
rect 19248 4088 19300 4140
rect 19524 4088 19576 4140
rect 20628 4088 20680 4140
rect 24308 4088 24360 4140
rect 24768 4088 24820 4140
rect 27896 4088 27948 4140
rect 28908 4088 28960 4140
rect 33876 4088 33928 4140
rect 34428 4088 34480 4140
rect 37372 4088 37424 4140
rect 38568 4088 38620 4140
rect 42156 4088 42208 4140
rect 42708 4088 42760 4140
rect 44548 4088 44600 4140
rect 45468 4088 45520 4140
rect 46940 4088 46992 4140
rect 4068 4020 4120 4072
rect 9036 4020 9088 4072
rect 43352 4020 43404 4072
rect 112076 4020 112128 4072
rect 113548 4088 113600 4140
rect 114468 4088 114520 4140
rect 115940 4088 115992 4140
rect 117228 4088 117280 4140
rect 149244 4088 149296 4140
rect 150348 4088 150400 4140
rect 153936 4088 153988 4140
rect 154488 4088 154540 4140
rect 158720 4088 158772 4140
rect 159916 4088 159968 4140
rect 163504 4088 163556 4140
rect 164148 4088 164200 4140
rect 114560 4020 114612 4072
rect 125416 4020 125468 4072
rect 167092 4088 167144 4140
rect 168196 4088 168248 4140
rect 170588 4088 170640 4140
rect 171048 4088 171100 4140
rect 174176 4088 174228 4140
rect 175188 4088 175240 4140
rect 236000 4088 236052 4140
rect 251180 4088 251232 4140
rect 252744 4088 252796 4140
rect 262220 4088 262272 4140
rect 271696 4088 271748 4140
rect 276020 4088 276072 4140
rect 277676 4088 277728 4140
rect 280344 4088 280396 4140
rect 284760 4088 284812 4140
rect 285680 4088 285732 4140
rect 288532 4088 288584 4140
rect 289544 4088 289596 4140
rect 289912 4088 289964 4140
rect 290740 4088 290792 4140
rect 291292 4088 291344 4140
rect 291936 4088 291988 4140
rect 295248 4088 295300 4140
rect 296720 4088 296772 4140
rect 303528 4088 303580 4140
rect 307392 4088 307444 4140
rect 402888 4088 402940 4140
rect 446588 4088 446640 4140
rect 474648 4088 474700 4140
rect 546500 4088 546552 4140
rect 36176 3952 36228 4004
rect 107660 3952 107712 4004
rect 121828 3952 121880 4004
rect 168380 4020 168432 4072
rect 200396 4020 200448 4072
rect 225052 4020 225104 4072
rect 227812 4020 227864 4072
rect 244280 4020 244332 4072
rect 249156 4020 249208 4072
rect 259460 4020 259512 4072
rect 275284 4020 275336 4072
rect 278688 4020 278740 4072
rect 278872 4020 278924 4072
rect 281540 4020 281592 4072
rect 282460 4020 282512 4072
rect 284300 4020 284352 4072
rect 296628 4020 296680 4072
rect 297916 4020 297968 4072
rect 306288 4020 306340 4072
rect 310980 4020 311032 4072
rect 314568 4020 314620 4072
rect 322848 4020 322900 4072
rect 408408 4020 408460 4072
rect 453672 4020 453724 4072
rect 477408 4020 477460 4072
rect 550088 4020 550140 4072
rect 203892 3952 203944 4004
rect 227720 3952 227772 4004
rect 231308 3952 231360 4004
rect 247040 3952 247092 4004
rect 247960 3952 248012 4004
rect 259552 3952 259604 4004
rect 304908 3952 304960 4004
rect 309784 3952 309836 4004
rect 313096 3952 313148 4004
rect 320456 3952 320508 4004
rect 321468 3952 321520 4004
rect 332416 3952 332468 4004
rect 346308 3952 346360 4004
rect 368020 3952 368072 4004
rect 405648 3952 405700 4004
rect 450176 3952 450228 4004
rect 480168 3952 480220 4004
rect 553584 3952 553636 4004
rect 39764 3884 39816 3936
rect 110420 3884 110472 3936
rect 118240 3884 118292 3936
rect 29092 3816 29144 3868
rect 30288 3816 30340 3868
rect 32680 3816 32732 3868
rect 25504 3748 25556 3800
rect 99380 3748 99432 3800
rect 114744 3816 114796 3868
rect 164240 3884 164292 3936
rect 171324 3884 171376 3936
rect 193220 3884 193272 3936
rect 219532 3884 219584 3936
rect 225328 3884 225380 3936
rect 242900 3884 242952 3936
rect 243176 3884 243228 3936
rect 255412 3884 255464 3936
rect 259828 3884 259880 3936
rect 267740 3884 267792 3936
rect 303436 3884 303488 3936
rect 308588 3884 308640 3936
rect 311808 3884 311860 3936
rect 319260 3884 319312 3936
rect 324228 3884 324280 3936
rect 335912 3884 335964 3936
rect 343548 3884 343600 3936
rect 364524 3884 364576 3936
rect 157524 3816 157576 3868
rect 158628 3816 158680 3868
rect 196808 3816 196860 3868
rect 222200 3816 222252 3868
rect 228916 3816 228968 3868
rect 245660 3816 245712 3868
rect 246764 3816 246816 3868
rect 258356 3816 258408 3868
rect 262220 3816 262272 3868
rect 269304 3816 269356 3868
rect 328368 3816 328420 3868
rect 341892 3816 341944 3868
rect 349068 3816 349120 3868
rect 371608 3884 371660 3936
rect 411168 3884 411220 3936
rect 457260 3884 457312 3936
rect 482928 3884 482980 3936
rect 557172 3884 557224 3936
rect 365720 3816 365772 3868
rect 366916 3816 366968 3868
rect 413928 3816 413980 3868
rect 460848 3816 460900 3868
rect 485688 3816 485740 3868
rect 560760 3816 560812 3868
rect 104900 3748 104952 3800
rect 111156 3748 111208 3800
rect 161480 3748 161532 3800
rect 189632 3748 189684 3800
rect 218060 3748 218112 3800
rect 241980 3748 242032 3800
rect 255320 3748 255372 3800
rect 256240 3748 256292 3800
rect 264980 3748 265032 3800
rect 276480 3748 276532 3800
rect 280160 3748 280212 3800
rect 317328 3748 317380 3800
rect 327632 3748 327684 3800
rect 328092 3748 328144 3800
rect 343088 3748 343140 3800
rect 351828 3748 351880 3800
rect 375196 3748 375248 3800
rect 415124 3748 415176 3800
rect 464436 3748 464488 3800
rect 487068 3748 487120 3800
rect 564348 3748 564400 3800
rect 20720 3680 20772 3732
rect 96620 3680 96672 3732
rect 107476 3680 107528 3732
rect 158812 3680 158864 3732
rect 186044 3680 186096 3732
rect 215300 3680 215352 3732
rect 218152 3680 218204 3732
rect 237380 3680 237432 3732
rect 239588 3680 239640 3732
rect 252652 3680 252704 3732
rect 257436 3680 257488 3732
rect 266360 3680 266412 3732
rect 269304 3680 269356 3732
rect 274640 3680 274692 3732
rect 318708 3680 318760 3732
rect 328828 3680 328880 3732
rect 331128 3680 331180 3732
rect 346676 3680 346728 3732
rect 354588 3680 354640 3732
rect 378784 3680 378836 3732
rect 420828 3680 420880 3732
rect 471520 3680 471572 3732
rect 489828 3680 489880 3732
rect 567844 3680 567896 3732
rect 16028 3612 16080 3664
rect 92480 3612 92532 3664
rect 103980 3612 104032 3664
rect 155960 3612 156012 3664
rect 165804 3612 165856 3664
rect 182548 3612 182600 3664
rect 212540 3612 212592 3664
rect 221740 3612 221792 3664
rect 240140 3612 240192 3664
rect 245568 3612 245620 3664
rect 258080 3612 258132 3664
rect 268108 3612 268160 3664
rect 273260 3612 273312 3664
rect 320088 3612 320140 3664
rect 331220 3612 331272 3664
rect 333888 3612 333940 3664
rect 350264 3612 350316 3664
rect 357348 3612 357400 3664
rect 360108 3612 360160 3664
rect 385868 3612 385920 3664
rect 418068 3612 418120 3664
rect 467840 3612 467892 3664
rect 492588 3612 492640 3664
rect 571340 3612 571392 3664
rect 10048 3544 10100 3596
rect 10968 3544 11020 3596
rect 11244 3544 11296 3596
rect 89720 3544 89772 3596
rect 100484 3544 100536 3596
rect 6460 3476 6512 3528
rect 5264 3340 5316 3392
rect 45744 3408 45796 3460
rect 46848 3408 46900 3460
rect 50528 3408 50580 3460
rect 50988 3408 51040 3460
rect 51632 3408 51684 3460
rect 52368 3408 52420 3460
rect 52828 3408 52880 3460
rect 53748 3408 53800 3460
rect 54024 3408 54076 3460
rect 55128 3408 55180 3460
rect 68284 3408 68336 3460
rect 68928 3408 68980 3460
rect 69480 3408 69532 3460
rect 70308 3408 70360 3460
rect 70676 3408 70728 3460
rect 71688 3408 71740 3460
rect 76656 3476 76708 3528
rect 77208 3476 77260 3528
rect 77852 3476 77904 3528
rect 78588 3476 78640 3528
rect 81440 3476 81492 3528
rect 82636 3476 82688 3528
rect 84936 3476 84988 3528
rect 85488 3476 85540 3528
rect 86132 3476 86184 3528
rect 86868 3476 86920 3528
rect 88524 3476 88576 3528
rect 89628 3476 89680 3528
rect 94504 3476 94556 3528
rect 95148 3476 95200 3528
rect 95700 3476 95752 3528
rect 96528 3476 96580 3528
rect 98092 3476 98144 3528
rect 99196 3476 99248 3528
rect 101588 3476 101640 3528
rect 102048 3476 102100 3528
rect 150348 3544 150400 3596
rect 175372 3544 175424 3596
rect 207112 3544 207164 3596
rect 207480 3544 207532 3596
rect 230480 3544 230532 3596
rect 232504 3544 232556 3596
rect 248420 3544 248472 3596
rect 251456 3544 251508 3596
rect 262312 3544 262364 3596
rect 263416 3544 263468 3596
rect 58808 3340 58860 3392
rect 59268 3340 59320 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 62396 3340 62448 3392
rect 63408 3340 63460 3392
rect 93308 3408 93360 3460
rect 145656 3476 145708 3528
rect 146208 3476 146260 3528
rect 146852 3476 146904 3528
rect 147588 3476 147640 3528
rect 150440 3476 150492 3528
rect 151728 3476 151780 3528
rect 164700 3476 164752 3528
rect 165528 3476 165580 3528
rect 178960 3476 179012 3528
rect 209964 3476 210016 3528
rect 63592 3272 63644 3324
rect 64788 3272 64840 3324
rect 55220 3204 55272 3256
rect 56508 3204 56560 3256
rect 96896 3340 96948 3392
rect 105176 3340 105228 3392
rect 106188 3340 106240 3392
rect 106372 3340 106424 3392
rect 107568 3340 107620 3392
rect 119436 3340 119488 3392
rect 119988 3340 120040 3392
rect 120632 3340 120684 3392
rect 121368 3340 121420 3392
rect 123024 3340 123076 3392
rect 124128 3340 124180 3392
rect 124220 3340 124272 3392
rect 125508 3340 125560 3392
rect 127808 3340 127860 3392
rect 128268 3340 128320 3392
rect 129004 3340 129056 3392
rect 129648 3340 129700 3392
rect 131396 3340 131448 3392
rect 132408 3340 132460 3392
rect 136088 3340 136140 3392
rect 136548 3340 136600 3392
rect 137284 3340 137336 3392
rect 137928 3340 137980 3392
rect 138480 3340 138532 3392
rect 139308 3340 139360 3392
rect 139676 3340 139728 3392
rect 140688 3340 140740 3392
rect 140872 3340 140924 3392
rect 141976 3340 142028 3392
rect 153476 3408 153528 3460
rect 171784 3408 171836 3460
rect 204444 3408 204496 3460
rect 209872 3408 209924 3460
rect 211068 3408 211120 3460
rect 148048 3340 148100 3392
rect 188436 3340 188488 3392
rect 188988 3340 189040 3392
rect 190828 3340 190880 3392
rect 191748 3340 191800 3392
rect 192024 3340 192076 3392
rect 193128 3340 193180 3392
rect 198004 3340 198056 3392
rect 198648 3340 198700 3392
rect 199200 3340 199252 3392
rect 200028 3340 200080 3392
rect 233424 3408 233476 3460
rect 236184 3476 236236 3528
rect 238392 3476 238444 3528
rect 252560 3476 252612 3528
rect 253848 3476 253900 3528
rect 263600 3476 263652 3528
rect 264612 3544 264664 3596
rect 270500 3544 270552 3596
rect 285956 3544 286008 3596
rect 287060 3544 287112 3596
rect 313188 3544 313240 3596
rect 321652 3544 321704 3596
rect 322940 3544 322992 3596
rect 334716 3544 334768 3596
rect 336556 3544 336608 3596
rect 347780 3544 347832 3596
rect 349068 3544 349120 3596
rect 382372 3544 382424 3596
rect 426072 3544 426124 3596
rect 478696 3544 478748 3596
rect 495164 3544 495216 3596
rect 571432 3544 571484 3596
rect 572628 3544 572680 3596
rect 270592 3476 270644 3528
rect 272892 3476 272944 3528
rect 277400 3476 277452 3528
rect 300768 3476 300820 3528
rect 303804 3476 303856 3528
rect 306196 3476 306248 3528
rect 312176 3476 312228 3528
rect 315948 3476 316000 3528
rect 325240 3476 325292 3528
rect 325516 3476 325568 3528
rect 338304 3476 338356 3528
rect 339408 3476 339460 3528
rect 357348 3476 357400 3528
rect 364248 3476 364300 3528
rect 393044 3476 393096 3528
rect 423588 3476 423640 3528
rect 475108 3476 475160 3528
rect 494060 3476 494112 3528
rect 495348 3476 495400 3528
rect 498108 3476 498160 3528
rect 578608 3476 578660 3528
rect 234804 3408 234856 3460
rect 249800 3408 249852 3460
rect 255044 3408 255096 3460
rect 265072 3408 265124 3460
rect 267004 3408 267056 3460
rect 273352 3408 273404 3460
rect 280068 3408 280120 3460
rect 282920 3408 282972 3460
rect 292488 3408 292540 3460
rect 293132 3408 293184 3460
rect 314476 3408 314528 3460
rect 324044 3408 324096 3460
rect 325608 3408 325660 3460
rect 339500 3408 339552 3460
rect 342168 3408 342220 3460
rect 360936 3408 360988 3460
rect 361488 3408 361540 3460
rect 389456 3408 389508 3460
rect 429108 3408 429160 3460
rect 482284 3408 482336 3460
rect 500868 3408 500920 3460
rect 582196 3408 582248 3460
rect 217048 3340 217100 3392
rect 217968 3340 218020 3392
rect 224132 3340 224184 3392
rect 241612 3340 241664 3392
rect 250352 3340 250404 3392
rect 261024 3340 261076 3392
rect 270500 3340 270552 3392
rect 276112 3340 276164 3392
rect 299296 3340 299348 3392
rect 302608 3340 302660 3392
rect 353760 3340 353812 3392
rect 451280 3340 451332 3392
rect 452476 3340 452528 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 512000 3340 512052 3392
rect 513196 3340 513248 3392
rect 528560 3340 528612 3392
rect 529848 3340 529900 3392
rect 575020 3340 575072 3392
rect 102784 3272 102836 3324
rect 103428 3272 103480 3324
rect 211068 3272 211120 3324
rect 214656 3272 214708 3324
rect 258632 3272 258684 3324
rect 266544 3272 266596 3324
rect 302056 3272 302108 3324
rect 306196 3272 306248 3324
rect 307668 3272 307720 3324
rect 314568 3272 314620 3324
rect 574744 3272 574796 3324
rect 576216 3272 576268 3324
rect 85672 3204 85724 3256
rect 181352 3204 181404 3256
rect 182088 3204 182140 3256
rect 80244 3136 80296 3188
rect 81348 3136 81400 3188
rect 148048 3136 148100 3188
rect 148968 3136 149020 3188
rect 155132 3136 155184 3188
rect 155868 3136 155920 3188
rect 265808 3136 265860 3188
rect 293868 3136 293920 3188
rect 294328 3136 294380 3188
rect 302148 3136 302200 3188
rect 305000 3136 305052 3188
rect 26700 3068 26752 3120
rect 27528 3068 27580 3120
rect 298008 3068 298060 3120
rect 300308 3068 300360 3120
rect 34980 3000 35032 3052
rect 35808 3000 35860 3052
rect 89720 3000 89772 3052
rect 91008 3000 91060 3052
rect 261024 3000 261076 3052
rect 269120 3000 269172 3052
rect 274088 3000 274140 3052
rect 277584 3000 277636 3052
rect 281264 3000 281316 3052
rect 283104 3000 283156 3052
rect 299388 3000 299440 3052
rect 301412 3000 301464 3052
rect 309048 3000 309100 3052
rect 315764 3000 315816 3052
rect 307576 2932 307628 2984
rect 313372 2932 313424 2984
rect 87328 2864 87380 2916
rect 88248 2864 88300 2916
rect 156328 2864 156380 2916
rect 157248 2864 157300 2916
rect 296536 2864 296588 2916
rect 299112 2864 299164 2916
rect 572 2796 624 2848
rect 1400 2796 1452 2848
rect 14832 2796 14884 2848
rect 15108 2796 15160 2848
rect 23112 2796 23164 2848
rect 23388 2796 23440 2848
rect 40960 2796 41012 2848
rect 41328 2796 41380 2848
rect 83832 2796 83884 2848
rect 84108 2796 84160 2848
rect 177948 2796 178000 2848
rect 310428 2660 310480 2712
rect 316960 2660 317012 2712
rect 206284 1096 206336 1148
rect 206928 1096 206980 1148
rect 31484 595 31536 604
rect 31484 561 31493 595
rect 31493 561 31527 595
rect 31527 561 31536 595
rect 31484 552 31536 561
rect 109960 552 110012 604
rect 110328 552 110380 604
rect 151544 595 151596 604
rect 151544 561 151553 595
rect 151553 561 151587 595
rect 151587 561 151596 595
rect 151544 552 151596 561
rect 161112 552 161164 604
rect 161388 552 161440 604
rect 177764 595 177816 604
rect 177764 561 177773 595
rect 177773 561 177807 595
rect 177807 561 177816 595
rect 177764 552 177816 561
rect 287152 552 287204 604
rect 287336 552 287388 604
rect 351920 552 351972 604
rect 352564 552 352616 604
rect 358544 595 358596 604
rect 358544 561 358553 595
rect 358553 561 358587 595
rect 358587 561 358596 595
rect 358544 552 358596 561
rect 359740 595 359792 604
rect 359740 561 359749 595
rect 359749 561 359783 595
rect 359783 561 359792 595
rect 359740 552 359792 561
rect 406108 595 406160 604
rect 406108 561 406117 595
rect 406117 561 406151 595
rect 406151 561 406160 595
rect 406108 552 406160 561
rect 407304 595 407356 604
rect 407304 561 407313 595
rect 407313 561 407347 595
rect 407347 561 407356 595
rect 407304 552 407356 561
rect 414480 595 414532 604
rect 414480 561 414489 595
rect 414489 561 414523 595
rect 414523 561 414532 595
rect 414480 552 414532 561
rect 431132 595 431184 604
rect 431132 561 431141 595
rect 431141 561 431175 595
rect 431175 561 431184 595
rect 431132 552 431184 561
rect 432328 595 432380 604
rect 432328 561 432337 595
rect 432337 561 432371 595
rect 432371 561 432380 595
rect 432328 552 432380 561
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 8128 679046 8156 685850
rect 8944 681760 8996 681766
rect 8944 681702 8996 681708
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3238 624880 3294 624889
rect 3238 624815 3294 624824
rect 3252 623830 3280 624815
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 3436 585138 3464 667927
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 3514 610464 3570 610473
rect 3514 610399 3570 610408
rect 3424 585132 3476 585138
rect 3424 585074 3476 585080
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 514758 3464 553007
rect 3528 550594 3556 610399
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 603770 8064 605798
rect 8024 603764 8076 603770
rect 8024 603706 8076 603712
rect 8956 596154 8984 681702
rect 14464 652792 14516 652798
rect 14464 652734 14516 652740
rect 10324 623824 10376 623830
rect 10324 623766 10376 623772
rect 8944 596148 8996 596154
rect 8944 596090 8996 596096
rect 9036 594856 9088 594862
rect 9036 594798 9088 594804
rect 9048 567866 9076 594798
rect 9036 567860 9088 567866
rect 9036 567802 9088 567808
rect 8944 567248 8996 567254
rect 8944 567190 8996 567196
rect 3516 550588 3568 550594
rect 3516 550530 3568 550536
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3424 514752 3476 514758
rect 3424 514694 3476 514700
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 3436 492658 3464 509895
rect 3528 503674 3556 538591
rect 8956 527134 8984 567190
rect 10336 561678 10364 623766
rect 14476 574054 14504 652734
rect 24780 603838 24808 699654
rect 41340 603906 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 73068 627972 73120 627978
rect 73068 627914 73120 627920
rect 73080 603974 73108 627914
rect 89640 604042 89668 699654
rect 106200 604110 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 137756 604178 137784 605798
rect 137744 604172 137796 604178
rect 137744 604114 137796 604120
rect 106188 604104 106240 604110
rect 106188 604046 106240 604052
rect 89628 604036 89680 604042
rect 89628 603978 89680 603984
rect 73068 603968 73120 603974
rect 73068 603910 73120 603916
rect 41328 603900 41380 603906
rect 41328 603842 41380 603848
rect 24768 603832 24820 603838
rect 24768 603774 24820 603780
rect 154316 603770 154344 605798
rect 169944 603900 169996 603906
rect 169944 603842 169996 603848
rect 156420 603832 156472 603838
rect 156420 603774 156472 603780
rect 142896 603764 142948 603770
rect 142896 603706 142948 603712
rect 154304 603764 154356 603770
rect 154304 603706 154356 603712
rect 142908 601868 142936 603706
rect 156432 601868 156460 603774
rect 169956 601868 169984 603842
rect 171060 603838 171088 700198
rect 197084 604036 197136 604042
rect 197084 603978 197136 603984
rect 183468 603968 183520 603974
rect 183468 603910 183520 603916
rect 171048 603832 171100 603838
rect 171048 603774 171100 603780
rect 183480 601868 183508 603910
rect 197096 601868 197124 603978
rect 202800 603906 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219348 627972 219400 627978
rect 219348 627914 219400 627920
rect 210608 604104 210660 604110
rect 210608 604046 210660 604052
rect 202788 603900 202840 603906
rect 202788 603842 202840 603848
rect 210620 601868 210648 604046
rect 219360 603974 219388 627914
rect 224132 604172 224184 604178
rect 224132 604114 224184 604120
rect 219348 603968 219400 603974
rect 219348 603910 219400 603916
rect 224144 601868 224172 604114
rect 235920 604042 235948 699654
rect 235908 604036 235960 604042
rect 235908 603978 235960 603984
rect 264796 603900 264848 603906
rect 264796 603842 264848 603848
rect 251272 603832 251324 603838
rect 251272 603774 251324 603780
rect 237656 603764 237708 603770
rect 237656 603706 237708 603712
rect 237668 601868 237696 603706
rect 251284 601868 251312 603774
rect 264808 601868 264836 603842
rect 267660 603770 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654158 284064 663734
rect 284024 654152 284076 654158
rect 284024 654094 284076 654100
rect 284208 654152 284260 654158
rect 284208 654094 284260 654100
rect 284220 644450 284248 654094
rect 284036 644422 284248 644450
rect 284036 634846 284064 644422
rect 284024 634840 284076 634846
rect 284024 634782 284076 634788
rect 284208 634840 284260 634846
rect 284208 634782 284260 634788
rect 284220 625138 284248 634782
rect 284036 625110 284248 625138
rect 284036 615534 284064 625110
rect 284024 615528 284076 615534
rect 284024 615470 284076 615476
rect 284208 615528 284260 615534
rect 284208 615470 284260 615476
rect 284220 605826 284248 615470
rect 284036 605798 284248 605826
rect 278320 603968 278372 603974
rect 278320 603910 278372 603916
rect 267648 603764 267700 603770
rect 267648 603706 267700 603712
rect 278332 601868 278360 603910
rect 284036 603838 284064 605798
rect 291844 604036 291896 604042
rect 291844 603978 291896 603984
rect 284024 603832 284076 603838
rect 284024 603774 284076 603780
rect 291856 601868 291884 603978
rect 300780 603906 300808 699654
rect 332520 620922 332548 703520
rect 348804 703474 348832 703520
rect 348712 703446 348832 703474
rect 348712 695502 348740 703446
rect 364996 699718 365024 703520
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 365628 699712 365680 699718
rect 365628 699654 365680 699660
rect 348700 695496 348752 695502
rect 348700 695438 348752 695444
rect 348792 685908 348844 685914
rect 348792 685850 348844 685856
rect 348804 678994 348832 685850
rect 348712 678966 348832 678994
rect 348712 676190 348740 678966
rect 348700 676184 348752 676190
rect 348700 676126 348752 676132
rect 348792 666596 348844 666602
rect 348792 666538 348844 666544
rect 348804 659682 348832 666538
rect 348804 659666 348924 659682
rect 348804 659660 348936 659666
rect 348804 659654 348884 659660
rect 348884 659602 348936 659608
rect 349068 659660 349120 659666
rect 349068 659602 349120 659608
rect 349080 656878 349108 659602
rect 349068 656872 349120 656878
rect 349068 656814 349120 656820
rect 348976 647284 349028 647290
rect 348976 647226 349028 647232
rect 348988 640422 349016 647226
rect 348976 640416 349028 640422
rect 348976 640358 349028 640364
rect 348792 640280 348844 640286
rect 348792 640222 348844 640228
rect 348804 637566 348832 640222
rect 348792 637560 348844 637566
rect 348792 637502 348844 637508
rect 349068 627972 349120 627978
rect 349068 627914 349120 627920
rect 332428 620894 332548 620922
rect 332428 611402 332456 620894
rect 332336 611374 332456 611402
rect 300768 603900 300820 603906
rect 300768 603842 300820 603848
rect 318984 603832 319036 603838
rect 318984 603774 319036 603780
rect 305460 603764 305512 603770
rect 305460 603706 305512 603712
rect 305472 601868 305500 603706
rect 318996 601868 319024 603774
rect 332336 603770 332364 611374
rect 332508 603900 332560 603906
rect 332508 603842 332560 603848
rect 332324 603764 332376 603770
rect 332324 603706 332376 603712
rect 332520 601868 332548 603842
rect 349080 603770 349108 627914
rect 346032 603764 346084 603770
rect 346032 603706 346084 603712
rect 349068 603764 349120 603770
rect 349068 603706 349120 603712
rect 359648 603764 359700 603770
rect 359648 603706 359700 603712
rect 346044 601868 346072 603706
rect 359660 601868 359688 603706
rect 365640 603294 365668 699654
rect 397472 603770 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 413756 698290 413784 703446
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 429856 684486 429884 703520
rect 429200 684480 429252 684486
rect 429200 684422 429252 684428
rect 429844 684480 429896 684486
rect 429844 684422 429896 684428
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 429212 683126 429240 684422
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 429200 683120 429252 683126
rect 429200 683062 429252 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 413112 659682 413140 666538
rect 429672 659682 429700 666538
rect 412928 659654 413140 659682
rect 429488 659654 429700 659682
rect 412928 647290 412956 659654
rect 429488 647290 429516 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 412836 640422 412864 647226
rect 429396 640422 429424 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 412928 630698 412956 640358
rect 429488 630698 429516 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 412744 630578 412772 630634
rect 429304 630578 429332 630634
rect 412744 630550 412864 630578
rect 429304 630550 429424 630578
rect 412836 621058 412864 630550
rect 429396 621058 429424 630550
rect 412836 621030 412956 621058
rect 429396 621030 429516 621058
rect 412928 611386 412956 621030
rect 429488 611386 429516 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 412744 603770 412772 611322
rect 427360 603900 427412 603906
rect 427360 603842 427412 603848
rect 386696 603764 386748 603770
rect 386696 603706 386748 603712
rect 397460 603764 397512 603770
rect 397460 603706 397512 603712
rect 400220 603764 400272 603770
rect 400220 603706 400272 603712
rect 412732 603764 412784 603770
rect 412732 603706 412784 603712
rect 413836 603764 413888 603770
rect 413836 603706 413888 603712
rect 365628 603288 365680 603294
rect 365628 603230 365680 603236
rect 373172 603288 373224 603294
rect 373172 603230 373224 603236
rect 373184 601868 373212 603230
rect 386708 601868 386736 603706
rect 400232 601868 400260 603706
rect 413848 601868 413876 603706
rect 427372 601868 427400 603842
rect 429304 603770 429332 611322
rect 462332 603906 462360 703520
rect 478524 703474 478552 703520
rect 494808 703474 494836 703520
rect 478524 703446 478644 703474
rect 494808 703446 494928 703474
rect 478616 692850 478644 703446
rect 494900 692850 494928 703446
rect 504364 696992 504416 696998
rect 504364 696934 504416 696940
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 477512 683074 477540 692786
rect 494072 683074 494100 692786
rect 477512 683046 477724 683074
rect 494072 683046 494284 683074
rect 477696 673538 477724 683046
rect 494256 673538 494284 683046
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 494060 673532 494112 673538
rect 494060 673474 494112 673480
rect 494244 673532 494296 673538
rect 494244 673474 494296 673480
rect 477512 663762 477540 673474
rect 494072 663762 494100 673474
rect 477512 663734 477724 663762
rect 494072 663734 494284 663762
rect 477696 654158 477724 663734
rect 494256 654158 494284 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 477512 644450 477540 654094
rect 494072 644450 494100 654094
rect 477512 644422 477724 644450
rect 494072 644422 494284 644450
rect 477696 634846 477724 644422
rect 494256 634846 494284 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 477512 625138 477540 634782
rect 494072 625138 494100 634782
rect 477512 625110 477724 625138
rect 494072 625110 494284 625138
rect 477696 615534 477724 625110
rect 494256 615534 494284 625110
rect 477500 615528 477552 615534
rect 477500 615470 477552 615476
rect 477684 615528 477736 615534
rect 477684 615470 477736 615476
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 477512 605826 477540 615470
rect 494072 605826 494100 615470
rect 477512 605798 477724 605826
rect 494072 605798 494284 605826
rect 462320 603900 462372 603906
rect 462320 603842 462372 603848
rect 468024 603900 468076 603906
rect 468024 603842 468076 603848
rect 440884 603832 440936 603838
rect 440884 603774 440936 603780
rect 429292 603764 429344 603770
rect 429292 603706 429344 603712
rect 440896 601868 440924 603774
rect 454408 603764 454460 603770
rect 454408 603706 454460 603712
rect 454420 601868 454448 603706
rect 468036 601868 468064 603842
rect 477696 603838 477724 605798
rect 477684 603832 477736 603838
rect 477684 603774 477736 603780
rect 481548 603832 481600 603838
rect 481548 603774 481600 603780
rect 481560 601868 481588 603774
rect 494256 603770 494284 605798
rect 494244 603764 494296 603770
rect 494244 603706 494296 603712
rect 495072 603764 495124 603770
rect 495072 603706 495124 603712
rect 495084 601868 495112 603706
rect 78680 596148 78732 596154
rect 78680 596090 78732 596096
rect 78692 596057 78720 596090
rect 78678 596048 78734 596057
rect 78678 595983 78734 595992
rect 504376 585585 504404 696934
rect 514024 673532 514076 673538
rect 514024 673474 514076 673480
rect 504362 585576 504418 585585
rect 504362 585511 504418 585520
rect 78680 585132 78732 585138
rect 78680 585074 78732 585080
rect 78692 584497 78720 585074
rect 78678 584488 78734 584497
rect 78678 584423 78734 584432
rect 514036 581670 514064 673474
rect 525064 650072 525116 650078
rect 525064 650014 525116 650020
rect 519544 626612 519596 626618
rect 519544 626554 519596 626560
rect 504364 581664 504416 581670
rect 504364 581606 504416 581612
rect 514024 581664 514076 581670
rect 514024 581606 514076 581612
rect 14464 574048 14516 574054
rect 14464 573990 14516 573996
rect 78680 574048 78732 574054
rect 78680 573990 78732 573996
rect 78692 572801 78720 573990
rect 78678 572792 78734 572801
rect 78678 572727 78734 572736
rect 79324 567860 79376 567866
rect 79324 567802 79376 567808
rect 10324 561672 10376 561678
rect 10324 561614 10376 561620
rect 78680 561672 78732 561678
rect 78680 561614 78732 561620
rect 78692 561241 78720 561614
rect 78678 561232 78734 561241
rect 78678 561167 78734 561176
rect 78680 550588 78732 550594
rect 78680 550530 78732 550536
rect 78692 549545 78720 550530
rect 78678 549536 78734 549545
rect 78678 549471 78734 549480
rect 79336 537985 79364 567802
rect 504376 563825 504404 581606
rect 514024 579692 514076 579698
rect 514024 579634 514076 579640
rect 505008 575476 505060 575482
rect 505008 575418 505060 575424
rect 505020 574705 505048 575418
rect 505006 574696 505062 574705
rect 505006 574631 505062 574640
rect 504362 563816 504418 563825
rect 504362 563751 504418 563760
rect 509884 556232 509936 556238
rect 509884 556174 509936 556180
rect 503812 553376 503864 553382
rect 503812 553318 503864 553324
rect 503824 552945 503852 553318
rect 503810 552936 503866 552945
rect 503810 552871 503866 552880
rect 505744 545148 505796 545154
rect 505744 545090 505796 545096
rect 505008 542360 505060 542366
rect 505008 542302 505060 542308
rect 505020 542065 505048 542302
rect 505006 542056 505062 542065
rect 505006 541991 505062 542000
rect 79322 537976 79378 537985
rect 79322 537911 79378 537920
rect 504364 537532 504416 537538
rect 504364 537474 504416 537480
rect 504376 531185 504404 537474
rect 504362 531176 504418 531185
rect 504362 531111 504418 531120
rect 8944 527128 8996 527134
rect 8944 527070 8996 527076
rect 78680 527128 78732 527134
rect 78680 527070 78732 527076
rect 78692 526289 78720 527070
rect 78678 526280 78734 526289
rect 78678 526215 78734 526224
rect 504640 521620 504692 521626
rect 504640 521562 504692 521568
rect 504652 520305 504680 521562
rect 504638 520296 504694 520305
rect 504638 520231 504694 520240
rect 78680 514752 78732 514758
rect 78678 514720 78680 514729
rect 78732 514720 78734 514729
rect 78678 514655 78734 514664
rect 505008 510604 505060 510610
rect 505008 510546 505060 510552
rect 505020 509425 505048 510546
rect 505006 509416 505062 509425
rect 505006 509351 505062 509360
rect 504364 508564 504416 508570
rect 504364 508506 504416 508512
rect 3516 503668 3568 503674
rect 3516 503610 3568 503616
rect 78680 503668 78732 503674
rect 78680 503610 78732 503616
rect 78692 503033 78720 503610
rect 78678 503024 78734 503033
rect 78678 502959 78734 502968
rect 3514 495544 3570 495553
rect 3514 495479 3570 495488
rect 3424 492652 3476 492658
rect 3424 492594 3476 492600
rect 3422 481128 3478 481137
rect 3422 481063 3478 481072
rect 3436 469198 3464 481063
rect 3528 480214 3556 495479
rect 78680 492652 78732 492658
rect 78680 492594 78732 492600
rect 78692 491473 78720 492594
rect 78678 491464 78734 491473
rect 78678 491399 78734 491408
rect 3516 480208 3568 480214
rect 3516 480150 3568 480156
rect 78680 480208 78732 480214
rect 78680 480150 78732 480156
rect 78692 479777 78720 480150
rect 78678 479768 78734 479777
rect 78678 479703 78734 479712
rect 503720 477284 503772 477290
rect 503720 477226 503772 477232
rect 503732 476921 503760 477226
rect 503718 476912 503774 476921
rect 503718 476847 503774 476856
rect 3424 469192 3476 469198
rect 3424 469134 3476 469140
rect 78680 469192 78732 469198
rect 78680 469134 78732 469140
rect 78692 468217 78720 469134
rect 78678 468208 78734 468217
rect 78678 468143 78734 468152
rect 78678 456512 78734 456521
rect 78678 456447 78734 456456
rect 78692 452606 78720 456447
rect 504376 455161 504404 508506
rect 505008 499520 505060 499526
rect 505008 499462 505060 499468
rect 505020 498545 505048 499462
rect 505006 498536 505062 498545
rect 505006 498471 505062 498480
rect 505006 487656 505062 487665
rect 505006 487591 505062 487600
rect 505020 487490 505048 487591
rect 505008 487484 505060 487490
rect 505008 487426 505060 487432
rect 505756 477290 505784 545090
rect 509896 487490 509924 556174
rect 514036 499526 514064 579634
rect 519556 537538 519584 626554
rect 520924 592068 520976 592074
rect 520924 592010 520976 592016
rect 519544 537532 519596 537538
rect 519544 537474 519596 537480
rect 519544 532772 519596 532778
rect 519544 532714 519596 532720
rect 514024 499520 514076 499526
rect 514024 499462 514076 499468
rect 509884 487484 509936 487490
rect 509884 487426 509936 487432
rect 514024 485852 514076 485858
rect 514024 485794 514076 485800
rect 505744 477284 505796 477290
rect 505744 477226 505796 477232
rect 505008 466404 505060 466410
rect 505008 466346 505060 466352
rect 505020 466041 505048 466346
rect 505006 466032 505062 466041
rect 505006 465967 505062 465976
rect 505744 462392 505796 462398
rect 505744 462334 505796 462340
rect 504362 455152 504418 455161
rect 504362 455087 504418 455096
rect 3424 452600 3476 452606
rect 3424 452542 3476 452548
rect 78680 452600 78732 452606
rect 78680 452542 78732 452548
rect 3436 452441 3464 452542
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 79322 444952 79378 444961
rect 79322 444887 79378 444896
rect 79336 438870 79364 444887
rect 505008 444372 505060 444378
rect 505008 444314 505060 444320
rect 505020 444281 505048 444314
rect 505006 444272 505062 444281
rect 505006 444207 505062 444216
rect 504364 438932 504416 438938
rect 504364 438874 504416 438880
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 79324 438864 79376 438870
rect 79324 438806 79376 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 79322 433256 79378 433265
rect 79322 433191 79378 433200
rect 79336 425066 79364 433191
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 79324 425060 79376 425066
rect 79324 425002 79376 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 503720 423496 503772 423502
rect 503720 423438 503772 423444
rect 503732 422521 503760 423438
rect 503718 422512 503774 422521
rect 503718 422447 503774 422456
rect 79414 421696 79470 421705
rect 79414 421631 79470 421640
rect 79322 398440 79378 398449
rect 79322 398375 79378 398384
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 79336 367062 79364 398375
rect 79428 396030 79456 421631
rect 79506 410000 79562 410009
rect 79506 409935 79562 409944
rect 79416 396024 79468 396030
rect 79416 395966 79468 395972
rect 79414 386744 79470 386753
rect 79414 386679 79470 386688
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 79324 367056 79376 367062
rect 79324 366998 79376 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 79322 363488 79378 363497
rect 79322 363423 79378 363432
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 78678 316976 78734 316985
rect 78678 316911 78734 316920
rect 78692 316062 78720 316911
rect 8944 316056 8996 316062
rect 8944 315998 8996 316004
rect 78680 316056 78732 316062
rect 78680 315998 78732 316004
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 3148 266348 3200 266354
rect 3148 266290 3200 266296
rect 3160 265713 3188 266290
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 8956 252482 8984 315998
rect 79336 309126 79364 363423
rect 79428 338094 79456 386679
rect 79520 380866 79548 409935
rect 504376 400761 504404 438874
rect 504640 434716 504692 434722
rect 504640 434658 504692 434664
rect 504652 433401 504680 434658
rect 504638 433392 504694 433401
rect 504638 433327 504694 433336
rect 505756 423502 505784 462334
rect 514036 434722 514064 485794
rect 519556 466410 519584 532714
rect 520936 510610 520964 592010
rect 525076 553382 525104 650014
rect 527192 603906 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 694142 542768 698226
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 692782 542584 694078
rect 542544 692776 542596 692782
rect 542544 692718 542596 692724
rect 542728 692776 542780 692782
rect 542728 692718 542780 692724
rect 542740 683233 542768 692718
rect 559668 684486 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 558920 684480 558972 684486
rect 558920 684422 558972 684428
rect 559656 684480 559708 684486
rect 559656 684422 559708 684428
rect 542358 683224 542414 683233
rect 542358 683159 542414 683168
rect 542726 683224 542782 683233
rect 542726 683159 542782 683168
rect 542372 683126 542400 683159
rect 558932 683126 558960 684422
rect 542360 683120 542412 683126
rect 542360 683062 542412 683068
rect 558920 683120 558972 683126
rect 558920 683062 558972 683068
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 542832 659682 542860 666538
rect 559392 659682 559420 666538
rect 542648 659654 542860 659682
rect 559208 659654 559420 659682
rect 542648 647290 542676 659654
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 542556 640422 542584 647226
rect 559116 640422 559144 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 542648 630698 542676 640358
rect 559208 630698 559236 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 542464 630578 542492 630634
rect 559024 630578 559052 630634
rect 542464 630550 542584 630578
rect 559024 630550 559144 630578
rect 542556 621058 542584 630550
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 559116 621030 559236 621058
rect 542648 611386 542676 621030
rect 559208 611386 559236 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 527180 603900 527232 603906
rect 527180 603842 527232 603848
rect 542464 603838 542492 611322
rect 542452 603832 542504 603838
rect 542452 603774 542504 603780
rect 559024 603770 559052 611322
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 559012 603764 559064 603770
rect 559012 603706 559064 603712
rect 580184 603158 580212 604143
rect 560944 603152 560996 603158
rect 560944 603094 560996 603100
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 525064 553376 525116 553382
rect 525064 553318 525116 553324
rect 560956 521626 560984 603094
rect 579894 592512 579950 592521
rect 579894 592447 579950 592456
rect 579908 592074 579936 592447
rect 579896 592068 579948 592074
rect 579896 592010 579948 592016
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580276 575482 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580264 575476 580316 575482
rect 580264 575418 580316 575424
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580368 542366 580396 639367
rect 580356 542360 580408 542366
rect 580356 542302 580408 542308
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 560944 521620 560996 521626
rect 560944 521562 560996 521568
rect 520924 510604 520976 510610
rect 520924 510546 520976 510552
rect 579986 510368 580042 510377
rect 579986 510303 580042 510312
rect 580000 509658 580028 510303
rect 578240 509652 578292 509658
rect 578240 509594 578292 509600
rect 579988 509652 580040 509658
rect 579988 509594 580040 509600
rect 578252 508570 578280 509594
rect 578240 508564 578292 508570
rect 578240 508506 578292 508512
rect 580262 498672 580318 498681
rect 580262 498607 580318 498616
rect 579894 486840 579950 486849
rect 579894 486775 579950 486784
rect 579908 485858 579936 486775
rect 579896 485852 579948 485858
rect 579896 485794 579948 485800
rect 519544 466404 519596 466410
rect 519544 466346 519596 466352
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580276 444378 580304 498607
rect 580354 451752 580410 451761
rect 580354 451687 580410 451696
rect 580264 444372 580316 444378
rect 580264 444314 580316 444320
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 514024 434716 514076 434722
rect 514024 434658 514076 434664
rect 505744 423496 505796 423502
rect 505744 423438 505796 423444
rect 580368 412622 580396 451687
rect 580446 416528 580502 416537
rect 580446 416463 580502 416472
rect 505008 412616 505060 412622
rect 505008 412558 505060 412564
rect 580356 412616 580408 412622
rect 580356 412558 580408 412564
rect 505020 411641 505048 412558
rect 505006 411632 505062 411641
rect 505006 411567 505062 411576
rect 580262 404832 580318 404841
rect 580262 404767 580318 404776
rect 504362 400752 504418 400761
rect 504362 400687 504418 400696
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 579908 392018 579936 392935
rect 514024 392012 514076 392018
rect 514024 391954 514076 391960
rect 579896 392012 579948 392018
rect 579896 391954 579948 391960
rect 505008 390516 505060 390522
rect 505008 390458 505060 390464
rect 505020 389881 505048 390458
rect 505006 389872 505062 389881
rect 505006 389807 505062 389816
rect 79508 380860 79560 380866
rect 79508 380802 79560 380808
rect 503904 379500 503956 379506
rect 503904 379442 503956 379448
rect 503916 379001 503944 379442
rect 503902 378992 503958 379001
rect 503902 378927 503958 378936
rect 79690 375184 79746 375193
rect 79690 375119 79746 375128
rect 79598 351928 79654 351937
rect 79598 351863 79654 351872
rect 79506 340232 79562 340241
rect 79506 340167 79562 340176
rect 79416 338088 79468 338094
rect 79416 338030 79468 338036
rect 79414 328672 79470 328681
rect 79414 328607 79470 328616
rect 79324 309120 79376 309126
rect 79324 309062 79376 309068
rect 79322 305416 79378 305425
rect 79322 305351 79378 305360
rect 78678 282160 78734 282169
rect 78678 282095 78734 282104
rect 78692 281586 78720 282095
rect 17224 281580 17276 281586
rect 17224 281522 17276 281528
rect 78680 281580 78732 281586
rect 78680 281522 78732 281528
rect 3240 252476 3292 252482
rect 3240 252418 3292 252424
rect 8944 252476 8996 252482
rect 8944 252418 8996 252424
rect 3252 251297 3280 252418
rect 3238 251288 3294 251297
rect 3238 251223 3294 251232
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 14464 223644 14516 223650
rect 14464 223586 14516 223592
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 8944 211200 8996 211206
rect 8944 211142 8996 211148
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 8956 122806 8984 211142
rect 10324 142180 10376 142186
rect 10324 142122 10376 142128
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 8944 122800 8996 122806
rect 8944 122742 8996 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 8944 100020 8996 100026
rect 8944 99962 8996 99968
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3424 80028 3476 80034
rect 3424 79970 3476 79976
rect 3436 78985 3464 79970
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1412 2854 1440 4762
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 584 480 612 2790
rect 1688 480 1716 5510
rect 2884 480 2912 8910
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7177 4108 8230
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 480 4108 4014
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5276 480 5304 3334
rect 6472 480 6500 3470
rect 7668 480 7696 6122
rect 8956 5574 8984 99962
rect 10336 35902 10364 142122
rect 14476 136610 14504 223586
rect 17236 208350 17264 281522
rect 78678 247208 78734 247217
rect 78678 247143 78734 247152
rect 78692 247110 78720 247143
rect 28264 247104 28316 247110
rect 28264 247046 28316 247052
rect 78680 247104 78732 247110
rect 78680 247046 78732 247052
rect 17224 208344 17276 208350
rect 17224 208286 17276 208292
rect 19984 189100 20036 189106
rect 19984 189042 20036 189048
rect 17224 176724 17276 176730
rect 17224 176666 17276 176672
rect 14464 136604 14516 136610
rect 14464 136546 14516 136552
rect 13728 94512 13780 94518
rect 13728 94454 13780 94460
rect 10416 49020 10468 49026
rect 10416 48962 10468 48968
rect 10324 35896 10376 35902
rect 10324 35838 10376 35844
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 480 8892 4082
rect 9048 4078 9076 17206
rect 10428 4146 10456 48962
rect 10968 36576 11020 36582
rect 10968 36518 11020 36524
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 10980 3602 11008 36518
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10060 480 10088 3538
rect 11256 480 11284 3538
rect 12452 480 12480 4082
rect 13648 480 13676 18566
rect 13740 4146 13768 94454
rect 17236 80034 17264 176666
rect 19996 93838 20024 189042
rect 28276 165578 28304 247046
rect 79336 237386 79364 305351
rect 79428 266354 79456 328607
rect 79520 280158 79548 340167
rect 79612 295322 79640 351863
rect 79704 324290 79732 375119
rect 514036 368490 514064 391954
rect 580276 379506 580304 404767
rect 580460 390522 580488 416463
rect 580448 390516 580500 390522
rect 580448 390458 580500 390464
rect 580264 379500 580316 379506
rect 580264 379442 580316 379448
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 505008 368484 505060 368490
rect 505008 368426 505060 368432
rect 514024 368484 514076 368490
rect 514024 368426 514076 368432
rect 505020 368121 505048 368426
rect 505006 368112 505062 368121
rect 505006 368047 505062 368056
rect 580276 357406 580304 369543
rect 580354 357912 580410 357921
rect 580354 357847 580410 357856
rect 505008 357400 505060 357406
rect 505006 357368 505008 357377
rect 580264 357400 580316 357406
rect 505060 357368 505062 357377
rect 580264 357342 580316 357348
rect 505006 357303 505062 357312
rect 580368 347750 580396 357847
rect 505008 347744 505060 347750
rect 505008 347686 505060 347692
rect 580356 347744 580408 347750
rect 580356 347686 580408 347692
rect 505020 346497 505048 347686
rect 505006 346488 505062 346497
rect 505006 346423 505062 346432
rect 580262 346080 580318 346089
rect 580262 346015 580318 346024
rect 580276 336734 580304 346015
rect 504548 336728 504600 336734
rect 504548 336670 504600 336676
rect 580264 336728 580316 336734
rect 580264 336670 580316 336676
rect 504560 335617 504588 336670
rect 504546 335608 504602 335617
rect 504546 335543 504602 335552
rect 505006 324728 505062 324737
rect 505006 324663 505062 324672
rect 79692 324284 79744 324290
rect 79692 324226 79744 324232
rect 505020 322930 505048 324663
rect 505008 322924 505060 322930
rect 505008 322866 505060 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 504086 313848 504142 313857
rect 504086 313783 504142 313792
rect 504100 311846 504128 313783
rect 504088 311840 504140 311846
rect 504088 311782 504140 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 504546 302968 504602 302977
rect 504546 302903 504602 302912
rect 504560 299470 504588 302903
rect 504548 299464 504600 299470
rect 504548 299406 504600 299412
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 79600 295316 79652 295322
rect 79600 295258 79652 295264
rect 79598 293720 79654 293729
rect 79598 293655 79654 293664
rect 79508 280152 79560 280158
rect 79508 280094 79560 280100
rect 79506 270464 79562 270473
rect 79506 270399 79562 270408
rect 79416 266348 79468 266354
rect 79416 266290 79468 266296
rect 79414 258904 79470 258913
rect 79414 258839 79470 258848
rect 79324 237380 79376 237386
rect 79324 237322 79376 237328
rect 79322 235648 79378 235657
rect 79322 235583 79378 235592
rect 78678 223952 78734 223961
rect 78678 223887 78734 223896
rect 78692 223650 78720 223887
rect 78680 223644 78732 223650
rect 78680 223586 78732 223592
rect 78678 212392 78734 212401
rect 78678 212327 78734 212336
rect 78692 211206 78720 212327
rect 78680 211200 78732 211206
rect 78680 211142 78732 211148
rect 78678 189136 78734 189145
rect 78678 189071 78680 189080
rect 78732 189071 78734 189080
rect 78680 189042 78732 189048
rect 78678 177440 78734 177449
rect 78678 177375 78734 177384
rect 78692 176730 78720 177375
rect 78680 176724 78732 176730
rect 78680 176666 78732 176672
rect 28264 165572 28316 165578
rect 28264 165514 28316 165520
rect 79336 151774 79364 235583
rect 79428 180810 79456 258839
rect 79520 194546 79548 270399
rect 79612 223582 79640 293655
rect 504362 292088 504418 292097
rect 504362 292023 504418 292032
rect 504376 276010 504404 292023
rect 504454 281208 504510 281217
rect 504454 281143 504510 281152
rect 504364 276004 504416 276010
rect 504364 275946 504416 275952
rect 504362 270328 504418 270337
rect 504362 270263 504418 270272
rect 504376 252550 504404 270263
rect 504468 264926 504496 281143
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 504456 264920 504508 264926
rect 504456 264862 504508 264868
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 504546 259448 504602 259457
rect 504546 259383 504602 259392
rect 504364 252544 504416 252550
rect 504364 252486 504416 252492
rect 504454 248568 504510 248577
rect 504454 248503 504510 248512
rect 504362 237688 504418 237697
rect 504362 237623 504418 237632
rect 79600 223576 79652 223582
rect 79600 223518 79652 223524
rect 504376 205630 504404 237623
rect 504468 218006 504496 248503
rect 504560 229090 504588 259383
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 504548 229084 504600 229090
rect 504548 229026 504600 229032
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 504638 226944 504694 226953
rect 504638 226879 504694 226888
rect 504456 218000 504508 218006
rect 504456 217942 504508 217948
rect 504546 216064 504602 216073
rect 504546 215999 504602 216008
rect 504364 205624 504416 205630
rect 504364 205566 504416 205572
rect 504454 205184 504510 205193
rect 504454 205119 504510 205128
rect 79690 200696 79746 200705
rect 79690 200631 79746 200640
rect 79508 194540 79560 194546
rect 79508 194482 79560 194488
rect 79416 180804 79468 180810
rect 79416 180746 79468 180752
rect 79598 165880 79654 165889
rect 79598 165815 79654 165824
rect 79506 154184 79562 154193
rect 79506 154119 79562 154128
rect 79324 151768 79376 151774
rect 79324 151710 79376 151716
rect 78678 142624 78734 142633
rect 78678 142559 78734 142568
rect 78692 142186 78720 142559
rect 78680 142180 78732 142186
rect 78680 142122 78732 142128
rect 79414 130928 79470 130937
rect 79414 130863 79470 130872
rect 79322 119368 79378 119377
rect 79322 119303 79378 119312
rect 75184 100088 75236 100094
rect 75184 100030 75236 100036
rect 52368 98660 52420 98666
rect 52368 98602 52420 98608
rect 19984 93832 20036 93838
rect 19984 93774 20036 93780
rect 22008 93152 22060 93158
rect 22008 93094 22060 93100
rect 17224 80028 17276 80034
rect 17224 79970 17276 79976
rect 17868 79348 17920 79354
rect 17868 79290 17920 79296
rect 15108 66904 15160 66910
rect 15108 66846 15160 66852
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 15120 2854 15148 66846
rect 17880 4146 17908 79290
rect 20628 46232 20680 46238
rect 20628 46174 20680 46180
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19260 4146 19288 19926
rect 20640 4146 20668 46174
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14844 480 14872 2790
rect 16040 480 16068 3606
rect 17236 480 17264 4082
rect 18340 480 18368 4082
rect 19536 480 19564 4082
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20732 480 20760 3674
rect 22020 2802 22048 93094
rect 27528 90364 27580 90370
rect 27528 90306 27580 90312
rect 24768 65544 24820 65550
rect 24768 65486 24820 65492
rect 23388 24132 23440 24138
rect 23388 24074 23440 24080
rect 23400 2854 23428 24074
rect 24780 4146 24808 65486
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 21928 2774 22048 2802
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 21928 480 21956 2774
rect 23124 480 23152 2790
rect 24320 480 24348 4082
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 25516 480 25544 3742
rect 27540 3126 27568 90306
rect 34428 89004 34480 89010
rect 34428 88946 34480 88952
rect 28908 76560 28960 76566
rect 28908 76502 28960 76508
rect 28920 4146 28948 76502
rect 31668 67652 31720 67658
rect 31668 67594 31720 67600
rect 31680 57934 31708 67594
rect 31668 57928 31720 57934
rect 31668 57870 31720 57876
rect 31668 48340 31720 48346
rect 31668 48282 31720 48288
rect 30288 47592 30340 47598
rect 30288 47534 30340 47540
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 26712 480 26740 3062
rect 27908 480 27936 4082
rect 29092 3868 29144 3874
rect 29092 3810 29144 3816
rect 29104 480 29132 3810
rect 30208 3618 30236 22714
rect 30300 3874 30328 47534
rect 31680 38622 31708 48282
rect 31668 38616 31720 38622
rect 31668 38558 31720 38564
rect 31668 29028 31720 29034
rect 31668 28970 31720 28976
rect 31680 19310 31708 28970
rect 31484 19304 31536 19310
rect 31484 19246 31536 19252
rect 31668 19304 31720 19310
rect 31668 19246 31720 19252
rect 31496 9761 31524 19246
rect 31482 9752 31538 9761
rect 31482 9687 31538 9696
rect 31666 9752 31722 9761
rect 31666 9687 31722 9696
rect 31680 9654 31708 9687
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 34440 4146 34468 88946
rect 38568 87644 38620 87650
rect 38568 87586 38620 87592
rect 38476 53100 38528 53106
rect 38476 53042 38528 53048
rect 35808 51740 35860 51746
rect 35808 51682 35860 51688
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 34428 4140 34480 4146
rect 34428 4082 34480 4088
rect 30288 3868 30340 3874
rect 30288 3810 30340 3816
rect 32680 3868 32732 3874
rect 32680 3810 32732 3816
rect 30208 3590 30328 3618
rect 30300 480 30328 3590
rect 31484 604 31536 610
rect 31484 546 31536 552
rect 31496 480 31524 546
rect 32692 480 32720 3810
rect 33888 480 33916 4082
rect 35820 3058 35848 51682
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 36176 4004 36228 4010
rect 36176 3946 36228 3952
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 35808 3052 35860 3058
rect 35808 2994 35860 3000
rect 34992 480 35020 2994
rect 36188 480 36216 3946
rect 37384 480 37412 4082
rect 38488 4026 38516 53042
rect 38580 4146 38608 87586
rect 49608 86284 49660 86290
rect 49608 86226 49660 86232
rect 42708 73840 42760 73846
rect 42708 73782 42760 73788
rect 41328 25560 41380 25566
rect 41328 25502 41380 25508
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38488 3998 38608 4026
rect 38580 480 38608 3998
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 39776 480 39804 3878
rect 41340 2854 41368 25502
rect 42720 4146 42748 73782
rect 46848 72480 46900 72486
rect 46848 72422 46900 72428
rect 45468 28280 45520 28286
rect 45468 28222 45520 28228
rect 45480 4146 45508 28222
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 44548 4140 44600 4146
rect 44548 4082 44600 4088
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 40960 2848 41012 2854
rect 40960 2790 41012 2796
rect 41328 2848 41380 2854
rect 41328 2790 41380 2796
rect 40972 480 41000 2790
rect 42168 480 42196 4082
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 43364 480 43392 4014
rect 44560 480 44588 4082
rect 46860 3466 46888 72422
rect 48228 10328 48280 10334
rect 48228 10270 48280 10276
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 45744 3460 45796 3466
rect 45744 3402 45796 3408
rect 46848 3460 46900 3466
rect 46848 3402 46900 3408
rect 45756 480 45784 3402
rect 46952 480 46980 4082
rect 48240 3482 48268 10270
rect 48148 3454 48268 3482
rect 48148 480 48176 3454
rect 49620 3346 49648 86226
rect 50988 37936 51040 37942
rect 50988 37878 51040 37884
rect 51000 3466 51028 37878
rect 52380 3466 52408 98602
rect 56508 97300 56560 97306
rect 56508 97242 56560 97248
rect 53748 84856 53800 84862
rect 53748 84798 53800 84804
rect 53760 3466 53788 84798
rect 55128 54528 55180 54534
rect 55128 54470 55180 54476
rect 55140 3466 55168 54470
rect 56416 31068 56468 31074
rect 56416 31010 56468 31016
rect 50528 3460 50580 3466
rect 50528 3402 50580 3408
rect 50988 3460 51040 3466
rect 50988 3402 51040 3408
rect 51632 3460 51684 3466
rect 51632 3402 51684 3408
rect 52368 3460 52420 3466
rect 52368 3402 52420 3408
rect 52828 3460 52880 3466
rect 52828 3402 52880 3408
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 54024 3460 54076 3466
rect 54024 3402 54076 3408
rect 55128 3460 55180 3466
rect 55128 3402 55180 3408
rect 49344 3318 49648 3346
rect 49344 480 49372 3318
rect 50540 480 50568 3402
rect 51644 480 51672 3402
rect 52840 480 52868 3402
rect 54036 480 54064 3402
rect 55220 3256 55272 3262
rect 55220 3198 55272 3204
rect 55232 480 55260 3198
rect 56428 480 56456 31010
rect 56520 3262 56548 97242
rect 73068 95940 73120 95946
rect 73068 95882 73120 95888
rect 64788 83496 64840 83502
rect 64788 83438 64840 83444
rect 57888 71052 57940 71058
rect 57888 70994 57940 71000
rect 57900 3482 57928 70994
rect 62028 69692 62080 69698
rect 62028 69634 62080 69640
rect 60648 32428 60700 32434
rect 60648 32370 60700 32376
rect 59268 11756 59320 11762
rect 59268 11698 59320 11704
rect 57624 3454 57928 3482
rect 56508 3256 56560 3262
rect 56508 3198 56560 3204
rect 57624 480 57652 3454
rect 59280 3398 59308 11698
rect 60660 3398 60688 32370
rect 62040 3398 62068 69634
rect 64696 39364 64748 39370
rect 64696 39306 64748 39312
rect 63408 13116 63460 13122
rect 63408 13058 63460 13064
rect 63420 3398 63448 13058
rect 58808 3392 58860 3398
rect 58808 3334 58860 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 62396 3392 62448 3398
rect 62396 3334 62448 3340
rect 63408 3392 63460 3398
rect 63408 3334 63460 3340
rect 58820 480 58848 3334
rect 60016 480 60044 3334
rect 61212 480 61240 3334
rect 62408 480 62436 3334
rect 63592 3324 63644 3330
rect 63592 3266 63644 3272
rect 63604 480 63632 3266
rect 64708 1578 64736 39306
rect 64800 3330 64828 83438
rect 67548 82136 67600 82142
rect 67548 82078 67600 82084
rect 66168 14476 66220 14482
rect 66168 14418 66220 14424
rect 66180 3482 66208 14418
rect 67560 3482 67588 82078
rect 71688 80708 71740 80714
rect 71688 80650 71740 80656
rect 68928 68332 68980 68338
rect 68928 68274 68980 68280
rect 65996 3454 66208 3482
rect 67192 3454 67588 3482
rect 68940 3466 68968 68274
rect 70308 26920 70360 26926
rect 70308 26862 70360 26868
rect 70320 3466 70348 26862
rect 71700 3466 71728 80650
rect 71872 7608 71924 7614
rect 71872 7550 71924 7556
rect 68284 3460 68336 3466
rect 64788 3324 64840 3330
rect 64788 3266 64840 3272
rect 64708 1550 64828 1578
rect 64800 480 64828 1550
rect 65996 480 66024 3454
rect 67192 480 67220 3454
rect 68284 3402 68336 3408
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 69480 3460 69532 3466
rect 69480 3402 69532 3408
rect 70308 3460 70360 3466
rect 70308 3402 70360 3408
rect 70676 3460 70728 3466
rect 70676 3402 70728 3408
rect 71688 3460 71740 3466
rect 71688 3402 71740 3408
rect 68296 480 68324 3402
rect 69492 480 69520 3402
rect 70688 480 70716 3402
rect 71884 480 71912 7550
rect 73080 480 73108 95882
rect 74448 77988 74500 77994
rect 74448 77930 74500 77936
rect 74460 3482 74488 77930
rect 75196 6186 75224 100030
rect 77944 99408 77996 99414
rect 77944 99350 77996 99356
rect 75828 57248 75880 57254
rect 75828 57190 75880 57196
rect 75184 6180 75236 6186
rect 75184 6122 75236 6128
rect 74276 3454 74488 3482
rect 74276 480 74304 3454
rect 75840 3346 75868 57190
rect 77208 15904 77260 15910
rect 77208 15846 77260 15852
rect 77220 3534 77248 15846
rect 77956 8974 77984 99350
rect 78588 33788 78640 33794
rect 78588 33730 78640 33736
rect 77944 8968 77996 8974
rect 77944 8910 77996 8916
rect 78600 3534 78628 33730
rect 79048 8968 79100 8974
rect 79048 8910 79100 8916
rect 76656 3528 76708 3534
rect 76656 3470 76708 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 77852 3528 77904 3534
rect 77852 3470 77904 3476
rect 78588 3528 78640 3534
rect 78588 3470 78640 3476
rect 75472 3318 75868 3346
rect 75472 480 75500 3318
rect 76668 480 76696 3470
rect 77864 480 77892 3470
rect 79060 480 79088 8910
rect 79336 8294 79364 119303
rect 79428 22098 79456 130863
rect 79520 51066 79548 154119
rect 79612 64870 79640 165815
rect 79704 109002 79732 200631
rect 504362 194304 504418 194313
rect 504362 194239 504418 194248
rect 504376 135250 504404 194239
rect 504468 158710 504496 205119
rect 504560 171086 504588 215999
rect 504652 182170 504680 226879
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 504822 183424 504878 183433
rect 504822 183359 504878 183368
rect 504640 182164 504692 182170
rect 504640 182106 504692 182112
rect 504730 172544 504786 172553
rect 504730 172479 504786 172488
rect 504548 171080 504600 171086
rect 504548 171022 504600 171028
rect 504638 161664 504694 161673
rect 504638 161599 504694 161608
rect 504456 158704 504508 158710
rect 504456 158646 504508 158652
rect 504546 150784 504602 150793
rect 504546 150719 504602 150728
rect 504364 135244 504416 135250
rect 504364 135186 504416 135192
rect 504454 129024 504510 129033
rect 504454 128959 504510 128968
rect 504362 118144 504418 118153
rect 504362 118079 504418 118088
rect 79692 108996 79744 109002
rect 79692 108938 79744 108944
rect 175568 102190 176226 102218
rect 184124 102190 184782 102218
rect 186608 102190 187358 102218
rect 188356 102190 189014 102218
rect 189184 102190 189934 102218
rect 190932 102190 191590 102218
rect 193508 102190 194166 102218
rect 243004 102190 243662 102218
rect 248984 102190 249642 102218
rect 251560 102190 252218 102218
rect 253216 102190 253874 102218
rect 277964 102190 278714 102218
rect 280540 102190 281198 102218
rect 284772 102190 285522 102218
rect 289096 102190 289754 102218
rect 350382 102190 350580 102218
rect 81452 102054 82386 102082
rect 79600 64864 79652 64870
rect 79600 64806 79652 64812
rect 79508 51060 79560 51066
rect 79508 51002 79560 51008
rect 81348 40724 81400 40730
rect 81348 40666 81400 40672
rect 79416 22092 79468 22098
rect 79416 22034 79468 22040
rect 79324 8288 79376 8294
rect 79324 8230 79376 8236
rect 81360 3194 81388 40666
rect 81452 4826 81480 102054
rect 83200 100026 83228 102068
rect 83188 100020 83240 100026
rect 83188 99962 83240 99968
rect 84028 99414 84056 102068
rect 84212 102054 84870 102082
rect 85684 102054 85790 102082
rect 86328 102054 86618 102082
rect 84016 99408 84068 99414
rect 84016 99350 84068 99356
rect 82728 58676 82780 58682
rect 82728 58618 82780 58624
rect 82636 35216 82688 35222
rect 82636 35158 82688 35164
rect 81440 4820 81492 4826
rect 81440 4762 81492 4768
rect 82648 3534 82676 35158
rect 81440 3528 81492 3534
rect 81440 3470 81492 3476
rect 82636 3528 82688 3534
rect 82636 3470 82688 3476
rect 80244 3188 80296 3194
rect 80244 3130 80296 3136
rect 81348 3188 81400 3194
rect 81348 3130 81400 3136
rect 80256 480 80284 3130
rect 81452 480 81480 3470
rect 82740 3210 82768 58618
rect 84108 29640 84160 29646
rect 84108 29582 84160 29588
rect 82648 3182 82768 3210
rect 82648 480 82676 3182
rect 84120 2854 84148 29582
rect 84212 17270 84240 102054
rect 85488 42084 85540 42090
rect 85488 42026 85540 42032
rect 84200 17264 84252 17270
rect 84200 17206 84252 17212
rect 85500 3534 85528 42026
rect 84936 3528 84988 3534
rect 84936 3470 84988 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 83832 2848 83884 2854
rect 83832 2790 83884 2796
rect 84108 2848 84160 2854
rect 84108 2790 84160 2796
rect 83844 480 83872 2790
rect 84948 480 84976 3470
rect 85684 3262 85712 102054
rect 86328 89842 86356 102054
rect 87432 100094 87460 102068
rect 87800 102054 88274 102082
rect 87420 100088 87472 100094
rect 87420 100030 87472 100036
rect 87800 89842 87828 102054
rect 88248 100020 88300 100026
rect 88248 99962 88300 99968
rect 88260 98666 88288 99962
rect 88248 98660 88300 98666
rect 88248 98602 88300 98608
rect 89180 96665 89208 102068
rect 89732 102054 90022 102082
rect 88522 96656 88578 96665
rect 88522 96591 88578 96600
rect 89166 96656 89222 96665
rect 89166 96591 89222 96600
rect 88248 91792 88300 91798
rect 88248 91734 88300 91740
rect 86144 89814 86356 89842
rect 87616 89814 87828 89842
rect 86144 86970 86172 89814
rect 86132 86964 86184 86970
rect 86132 86906 86184 86912
rect 87616 77314 87644 89814
rect 85856 77308 85908 77314
rect 85856 77250 85908 77256
rect 87236 77308 87288 77314
rect 87236 77250 87288 77256
rect 87604 77308 87656 77314
rect 87604 77250 87656 77256
rect 85868 77194 85896 77250
rect 85776 77166 85896 77194
rect 85776 67794 85804 77166
rect 85764 67788 85816 67794
rect 85764 67730 85816 67736
rect 87248 66314 87276 77250
rect 85764 66292 85816 66298
rect 85764 66234 85816 66240
rect 87156 66286 87276 66314
rect 85776 56574 85804 66234
rect 87156 66230 87184 66286
rect 87144 66224 87196 66230
rect 87144 66166 87196 66172
rect 87144 56636 87196 56642
rect 87144 56578 87196 56584
rect 85764 56568 85816 56574
rect 85764 56510 85816 56516
rect 87156 49026 87184 56578
rect 87144 49020 87196 49026
rect 87144 48962 87196 48968
rect 85764 47048 85816 47054
rect 85764 46990 85816 46996
rect 85776 46918 85804 46990
rect 85764 46912 85816 46918
rect 85764 46854 85816 46860
rect 86040 46912 86092 46918
rect 86040 46854 86092 46860
rect 86052 31634 86080 46854
rect 85960 31606 86080 31634
rect 85960 22166 85988 31606
rect 85948 22160 86000 22166
rect 85948 22102 86000 22108
rect 85764 22092 85816 22098
rect 85764 22034 85816 22040
rect 85776 9654 85804 22034
rect 86868 21412 86920 21418
rect 86868 21354 86920 21360
rect 85764 9648 85816 9654
rect 85764 9590 85816 9596
rect 86880 3534 86908 21354
rect 86132 3528 86184 3534
rect 86132 3470 86184 3476
rect 86868 3528 86920 3534
rect 86868 3470 86920 3476
rect 85672 3256 85724 3262
rect 85672 3198 85724 3204
rect 86144 480 86172 3470
rect 88260 2922 88288 91734
rect 88536 86970 88564 96591
rect 88524 86964 88576 86970
rect 88524 86906 88576 86912
rect 88524 77308 88576 77314
rect 88524 77250 88576 77256
rect 88536 66314 88564 77250
rect 88444 66286 88564 66314
rect 88444 66230 88472 66286
rect 88432 66224 88484 66230
rect 88432 66166 88484 66172
rect 88340 56636 88392 56642
rect 88340 56578 88392 56584
rect 88352 48346 88380 56578
rect 88340 48340 88392 48346
rect 88340 48282 88392 48288
rect 88432 48340 88484 48346
rect 88432 48282 88484 48288
rect 88444 41478 88472 48282
rect 89628 44872 89680 44878
rect 89628 44814 89680 44820
rect 88432 41472 88484 41478
rect 88432 41414 88484 41420
rect 88340 41404 88392 41410
rect 88340 41346 88392 41352
rect 88352 36582 88380 41346
rect 88340 36576 88392 36582
rect 88340 36518 88392 36524
rect 89640 3534 89668 44814
rect 89732 3602 89760 102054
rect 90836 94518 90864 102068
rect 91112 102054 91770 102082
rect 90824 94512 90876 94518
rect 90824 94454 90876 94460
rect 91008 60036 91060 60042
rect 91008 59978 91060 59984
rect 90916 43444 90968 43450
rect 90916 43386 90968 43392
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 88524 3528 88576 3534
rect 88524 3470 88576 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 87328 2916 87380 2922
rect 87328 2858 87380 2864
rect 88248 2916 88300 2922
rect 88248 2858 88300 2864
rect 87340 480 87368 2858
rect 88536 480 88564 3470
rect 89720 3052 89772 3058
rect 89720 2994 89772 3000
rect 89732 480 89760 2994
rect 90928 480 90956 43386
rect 91020 3058 91048 59978
rect 91112 18630 91140 102054
rect 91744 99408 91796 99414
rect 91744 99350 91796 99356
rect 91756 79354 91784 99350
rect 92480 94580 92532 94586
rect 92480 94522 92532 94528
rect 91744 79348 91796 79354
rect 91744 79290 91796 79296
rect 92388 79348 92440 79354
rect 92388 79290 92440 79296
rect 91100 18624 91152 18630
rect 91100 18566 91152 18572
rect 92400 3346 92428 79290
rect 92492 3670 92520 94522
rect 92584 66910 92612 102068
rect 93136 102054 93426 102082
rect 93136 94586 93164 102054
rect 94240 99414 94268 102068
rect 94516 102054 95174 102082
rect 95620 102054 96002 102082
rect 96632 102054 96830 102082
rect 97184 102054 97750 102082
rect 98012 102054 98578 102082
rect 94228 99408 94280 99414
rect 94228 99350 94280 99356
rect 93124 94580 93176 94586
rect 93124 94522 93176 94528
rect 94516 94466 94544 102054
rect 93964 94438 94544 94466
rect 93964 80186 93992 94438
rect 95620 87038 95648 102054
rect 95608 87032 95660 87038
rect 95608 86974 95660 86980
rect 95700 86896 95752 86902
rect 95700 86838 95752 86844
rect 93872 80158 93992 80186
rect 93872 80050 93900 80158
rect 93872 80022 93992 80050
rect 93964 79914 93992 80022
rect 93964 79886 94084 79914
rect 92572 66904 92624 66910
rect 92572 66846 92624 66852
rect 94056 48346 94084 79886
rect 95712 77466 95740 86838
rect 95712 77438 95832 77466
rect 95804 74526 95832 77438
rect 95792 74520 95844 74526
rect 95792 74462 95844 74468
rect 95516 64932 95568 64938
rect 95516 64874 95568 64880
rect 95528 60874 95556 64874
rect 95436 60846 95556 60874
rect 95436 55282 95464 60846
rect 95332 55276 95384 55282
rect 95332 55218 95384 55224
rect 95424 55276 95476 55282
rect 95424 55218 95476 55224
rect 95344 51082 95372 55218
rect 95344 51054 95464 51082
rect 93952 48340 94004 48346
rect 93952 48282 94004 48288
rect 94044 48340 94096 48346
rect 94044 48282 94096 48288
rect 93964 41426 93992 48282
rect 95436 46238 95464 51054
rect 95424 46232 95476 46238
rect 95424 46174 95476 46180
rect 96528 46232 96580 46238
rect 96528 46174 96580 46180
rect 93964 41398 94084 41426
rect 94056 31770 94084 41398
rect 94056 31742 94176 31770
rect 94148 19990 94176 31742
rect 94136 19984 94188 19990
rect 94136 19926 94188 19932
rect 95148 17264 95200 17270
rect 95148 17206 95200 17212
rect 92480 3664 92532 3670
rect 92480 3606 92532 3612
rect 95160 3534 95188 17206
rect 96540 3534 96568 46174
rect 96632 3738 96660 102054
rect 97184 93158 97212 102054
rect 97172 93152 97224 93158
rect 97172 93094 97224 93100
rect 98012 24138 98040 102054
rect 99392 94738 99420 102068
rect 99944 102054 100234 102082
rect 100864 102054 101154 102082
rect 99392 94710 99512 94738
rect 99380 94580 99432 94586
rect 99380 94522 99432 94528
rect 98000 24132 98052 24138
rect 98000 24074 98052 24080
rect 99196 18624 99248 18630
rect 99196 18566 99248 18572
rect 96620 3732 96672 3738
rect 96620 3674 96672 3680
rect 99208 3534 99236 18566
rect 99288 4820 99340 4826
rect 99288 4762 99340 4768
rect 94504 3528 94556 3534
rect 94504 3470 94556 3476
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 95700 3528 95752 3534
rect 95700 3470 95752 3476
rect 96528 3528 96580 3534
rect 96528 3470 96580 3476
rect 98092 3528 98144 3534
rect 98092 3470 98144 3476
rect 99196 3528 99248 3534
rect 99196 3470 99248 3476
rect 93308 3460 93360 3466
rect 93308 3402 93360 3408
rect 92124 3318 92428 3346
rect 91008 3052 91060 3058
rect 91008 2994 91060 3000
rect 92124 480 92152 3318
rect 93320 480 93348 3402
rect 94516 480 94544 3470
rect 95712 480 95740 3470
rect 96896 3392 96948 3398
rect 96896 3334 96948 3340
rect 96908 480 96936 3334
rect 98104 480 98132 3470
rect 99300 480 99328 4762
rect 99392 3806 99420 94522
rect 99484 65550 99512 94710
rect 99944 94586 99972 102054
rect 99932 94580 99984 94586
rect 99932 94522 99984 94528
rect 100864 90370 100892 102054
rect 101968 96665 101996 102068
rect 102152 102054 102810 102082
rect 103532 102054 103638 102082
rect 101586 96656 101642 96665
rect 101586 96591 101642 96600
rect 101954 96656 102010 96665
rect 101954 96591 102010 96600
rect 100852 90364 100904 90370
rect 100852 90306 100904 90312
rect 101600 80186 101628 96591
rect 101508 80158 101628 80186
rect 101508 80102 101536 80158
rect 100760 80096 100812 80102
rect 100760 80038 100812 80044
rect 101496 80096 101548 80102
rect 101496 80038 101548 80044
rect 100772 76566 100800 80038
rect 100760 76560 100812 76566
rect 100760 76502 100812 76508
rect 99472 65544 99524 65550
rect 99472 65486 99524 65492
rect 102152 47598 102180 102054
rect 102140 47592 102192 47598
rect 102140 47534 102192 47540
rect 103428 47592 103480 47598
rect 103428 47534 103480 47540
rect 102048 19984 102100 19990
rect 102048 19926 102100 19932
rect 99380 3800 99432 3806
rect 99380 3742 99432 3748
rect 100484 3596 100536 3602
rect 100484 3538 100536 3544
rect 100496 480 100524 3538
rect 102060 3534 102088 19926
rect 101588 3528 101640 3534
rect 101588 3470 101640 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 101600 480 101628 3470
rect 103440 3330 103468 47534
rect 103532 22778 103560 102054
rect 104544 96665 104572 102068
rect 104912 102054 105386 102082
rect 104070 96656 104126 96665
rect 104070 96591 104126 96600
rect 104530 96656 104586 96665
rect 104530 96591 104586 96600
rect 104084 77314 104112 96591
rect 103612 77308 103664 77314
rect 103612 77250 103664 77256
rect 104072 77308 104124 77314
rect 104072 77250 104124 77256
rect 103624 75206 103652 77250
rect 103612 75200 103664 75206
rect 103612 75142 103664 75148
rect 103520 22772 103572 22778
rect 103520 22714 103572 22720
rect 104912 3806 104940 102054
rect 106200 96665 106228 102068
rect 106924 99408 106976 99414
rect 106924 99350 106976 99356
rect 105542 96656 105598 96665
rect 105542 96591 105598 96600
rect 106186 96656 106242 96665
rect 106186 96591 106242 96600
rect 106646 96656 106702 96665
rect 106646 96591 106702 96600
rect 105556 89010 105584 96591
rect 105544 89004 105596 89010
rect 105544 88946 105596 88952
rect 106660 77314 106688 96591
rect 106280 77308 106332 77314
rect 106280 77250 106332 77256
rect 106648 77308 106700 77314
rect 106648 77250 106700 77256
rect 106292 70394 106320 77250
rect 106936 73846 106964 99350
rect 107120 96665 107148 102068
rect 107672 102054 107962 102082
rect 107106 96656 107162 96665
rect 107106 96591 107162 96600
rect 106924 73840 106976 73846
rect 106924 73782 106976 73788
rect 106292 70366 106504 70394
rect 106476 51746 106504 70366
rect 106464 51740 106516 51746
rect 106464 51682 106516 51688
rect 107568 50380 107620 50386
rect 107568 50322 107620 50328
rect 106188 24132 106240 24138
rect 106188 24074 106240 24080
rect 104900 3800 104952 3806
rect 104900 3742 104952 3748
rect 103980 3664 104032 3670
rect 103980 3606 104032 3612
rect 102784 3324 102836 3330
rect 102784 3266 102836 3272
rect 103428 3324 103480 3330
rect 103428 3266 103480 3272
rect 102796 480 102824 3266
rect 103992 480 104020 3606
rect 106200 3398 106228 24074
rect 107476 3732 107528 3738
rect 107476 3674 107528 3680
rect 105176 3392 105228 3398
rect 105176 3334 105228 3340
rect 106188 3392 106240 3398
rect 106188 3334 106240 3340
rect 106372 3392 106424 3398
rect 106372 3334 106424 3340
rect 105188 480 105216 3334
rect 106384 480 106412 3334
rect 107488 1850 107516 3674
rect 107580 3398 107608 50322
rect 107672 4010 107700 102054
rect 108776 96665 108804 102068
rect 109052 102054 109618 102082
rect 110432 102054 110538 102082
rect 110984 102054 111366 102082
rect 108302 96656 108358 96665
rect 108302 96591 108358 96600
rect 108762 96656 108818 96665
rect 108762 96591 108818 96600
rect 108316 87650 108344 96591
rect 108304 87644 108356 87650
rect 108304 87586 108356 87592
rect 109052 53106 109080 102054
rect 109040 53100 109092 53106
rect 109040 53042 109092 53048
rect 110328 51740 110380 51746
rect 110328 51682 110380 51688
rect 108948 22772 109000 22778
rect 108948 22714 109000 22720
rect 107660 4004 107712 4010
rect 107660 3946 107712 3952
rect 107568 3392 107620 3398
rect 107568 3334 107620 3340
rect 107488 1822 107608 1850
rect 107580 480 107608 1822
rect 108960 626 108988 22714
rect 108776 598 108988 626
rect 110340 610 110368 51682
rect 110432 3942 110460 102054
rect 110984 89842 111012 102054
rect 112180 99414 112208 102068
rect 112640 102054 113114 102082
rect 113468 102054 113942 102082
rect 114664 102054 114770 102082
rect 115216 102054 115598 102082
rect 115952 102054 116518 102082
rect 112168 99408 112220 99414
rect 112168 99350 112220 99356
rect 112640 89842 112668 102054
rect 113468 89842 113496 102054
rect 114560 94580 114612 94586
rect 114560 94522 114612 94528
rect 110800 89814 111012 89842
rect 112272 89814 112668 89842
rect 113376 89814 113496 89842
rect 110800 89706 110828 89814
rect 112272 89706 112300 89814
rect 110616 89678 110828 89706
rect 111996 89678 112300 89706
rect 110616 86970 110644 89678
rect 110604 86964 110656 86970
rect 110604 86906 110656 86912
rect 111996 80186 112024 89678
rect 111996 80158 112116 80186
rect 112088 77314 112116 80158
rect 110512 77308 110564 77314
rect 110512 77250 110564 77256
rect 111800 77308 111852 77314
rect 111800 77250 111852 77256
rect 112076 77308 112128 77314
rect 112076 77250 112128 77256
rect 110524 67658 110552 77250
rect 110512 67652 110564 67658
rect 110512 67594 110564 67600
rect 110604 67652 110656 67658
rect 110604 67594 110656 67600
rect 110616 60602 110644 67594
rect 111812 66230 111840 77250
rect 113376 70394 113404 89814
rect 113192 70366 113404 70394
rect 113192 70258 113220 70366
rect 113192 70230 113312 70258
rect 111800 66224 111852 66230
rect 111800 66166 111852 66172
rect 110616 60574 110736 60602
rect 110708 57934 110736 60574
rect 110696 57928 110748 57934
rect 110696 57870 110748 57876
rect 111892 56636 111944 56642
rect 111892 56578 111944 56584
rect 111904 51082 111932 56578
rect 113284 51082 113312 70230
rect 114468 53100 114520 53106
rect 114468 53042 114520 53048
rect 111812 51054 111932 51082
rect 113192 51066 113312 51082
rect 113180 51060 113312 51066
rect 110788 48340 110840 48346
rect 110788 48282 110840 48288
rect 110800 38690 110828 48282
rect 111812 48226 111840 51054
rect 113232 51054 113312 51060
rect 113364 51060 113416 51066
rect 113180 51002 113232 51008
rect 113364 51002 113416 51008
rect 113192 50971 113220 51002
rect 111812 48198 111932 48226
rect 111904 43330 111932 48198
rect 111812 43302 111932 43330
rect 111812 38729 111840 43302
rect 113376 41478 113404 51002
rect 113364 41472 113416 41478
rect 113364 41414 113416 41420
rect 113364 41336 113416 41342
rect 113364 41278 113416 41284
rect 111798 38720 111854 38729
rect 110696 38684 110748 38690
rect 110696 38626 110748 38632
rect 110788 38684 110840 38690
rect 111798 38655 111854 38664
rect 110788 38626 110840 38632
rect 110708 25566 110736 38626
rect 111798 38584 111854 38593
rect 111798 38519 111854 38528
rect 111812 29034 111840 38519
rect 111800 29028 111852 29034
rect 111800 28970 111852 28976
rect 112076 29028 112128 29034
rect 112076 28970 112128 28976
rect 110696 25560 110748 25566
rect 110696 25502 110748 25508
rect 112088 22114 112116 28970
rect 113376 28286 113404 41278
rect 113364 28280 113416 28286
rect 113364 28222 113416 28228
rect 111904 22098 112116 22114
rect 111892 22092 112128 22098
rect 111944 22086 112076 22092
rect 111892 22034 111944 22040
rect 112076 22034 112128 22040
rect 112088 19310 112116 22034
rect 112076 19304 112128 19310
rect 112076 19246 112128 19252
rect 112076 11892 112128 11898
rect 112076 11834 112128 11840
rect 112088 4078 112116 11834
rect 112352 6180 112404 6186
rect 112352 6122 112404 6128
rect 112076 4072 112128 4078
rect 112076 4014 112128 4020
rect 110420 3936 110472 3942
rect 110420 3878 110472 3884
rect 111156 3800 111208 3806
rect 111156 3742 111208 3748
rect 109960 604 110012 610
rect 108776 480 108804 598
rect 109960 546 110012 552
rect 110328 604 110380 610
rect 110328 546 110380 552
rect 109972 480 110000 546
rect 111168 480 111196 3742
rect 112364 480 112392 6122
rect 114480 4146 114508 53042
rect 113548 4140 113600 4146
rect 113548 4082 113600 4088
rect 114468 4140 114520 4146
rect 114468 4082 114520 4088
rect 113560 480 113588 4082
rect 114572 4078 114600 94522
rect 114664 72486 114692 102054
rect 115216 94586 115244 102054
rect 115204 94580 115256 94586
rect 115204 94522 115256 94528
rect 114652 72480 114704 72486
rect 114652 72422 114704 72428
rect 115952 10334 115980 102054
rect 117332 94738 117360 102068
rect 117792 102054 118174 102082
rect 117332 94710 117452 94738
rect 117320 94580 117372 94586
rect 117320 94522 117372 94528
rect 117332 37942 117360 94522
rect 117424 86290 117452 94710
rect 117792 94586 117820 102054
rect 118988 100026 119016 102068
rect 119632 102054 119922 102082
rect 120092 102054 120750 102082
rect 118976 100020 119028 100026
rect 118976 99962 119028 99968
rect 117780 94580 117832 94586
rect 117780 94522 117832 94528
rect 119632 89842 119660 102054
rect 119540 89814 119660 89842
rect 119540 89758 119568 89814
rect 118792 89752 118844 89758
rect 118792 89694 118844 89700
rect 119528 89752 119580 89758
rect 119528 89694 119580 89700
rect 117412 86284 117464 86290
rect 117412 86226 117464 86232
rect 118804 84862 118832 89694
rect 118792 84856 118844 84862
rect 118792 84798 118844 84804
rect 120092 54534 120120 102054
rect 120724 100020 120776 100026
rect 120724 99962 120776 99968
rect 120080 54528 120132 54534
rect 120080 54470 120132 54476
rect 117320 37936 117372 37942
rect 117320 37878 117372 37884
rect 119988 37936 120040 37942
rect 119988 37878 120040 37884
rect 117228 36576 117280 36582
rect 117228 36518 117280 36524
rect 117136 14544 117188 14550
rect 117136 14486 117188 14492
rect 115940 10328 115992 10334
rect 115940 10270 115992 10276
rect 115940 4140 115992 4146
rect 115940 4082 115992 4088
rect 114560 4072 114612 4078
rect 114560 4014 114612 4020
rect 114744 3868 114796 3874
rect 114744 3810 114796 3816
rect 114756 480 114784 3810
rect 115952 480 115980 4082
rect 117148 480 117176 14486
rect 117240 4146 117268 36518
rect 117228 4140 117280 4146
rect 117228 4082 117280 4088
rect 118240 3936 118292 3942
rect 118240 3878 118292 3884
rect 118252 480 118280 3878
rect 120000 3398 120028 37878
rect 120736 14482 120764 99962
rect 121564 97306 121592 102068
rect 121748 102054 122498 102082
rect 122944 102054 123326 102082
rect 123864 102054 124154 102082
rect 121552 97300 121604 97306
rect 121552 97242 121604 97248
rect 121748 89842 121776 102054
rect 122840 94580 122892 94586
rect 122840 94522 122892 94528
rect 121656 89814 121776 89842
rect 121656 70394 121684 89814
rect 121472 70366 121684 70394
rect 121472 70258 121500 70366
rect 121472 70230 121592 70258
rect 121368 54528 121420 54534
rect 121368 54470 121420 54476
rect 120724 14476 120776 14482
rect 120724 14418 120776 14424
rect 121380 3398 121408 54470
rect 121564 51082 121592 70230
rect 121472 51066 121592 51082
rect 121460 51060 121592 51066
rect 121512 51054 121592 51060
rect 121644 51060 121696 51066
rect 121460 51002 121512 51008
rect 121644 51002 121696 51008
rect 121472 50971 121500 51002
rect 121656 48278 121684 51002
rect 121644 48272 121696 48278
rect 121644 48214 121696 48220
rect 121736 38684 121788 38690
rect 121736 38626 121788 38632
rect 121748 31074 121776 38626
rect 121736 31068 121788 31074
rect 121736 31010 121788 31016
rect 122852 11762 122880 94522
rect 122944 71058 122972 102054
rect 123864 94586 123892 102054
rect 124864 100088 124916 100094
rect 124864 100030 124916 100036
rect 124402 96656 124458 96665
rect 124402 96591 124458 96600
rect 123852 94580 123904 94586
rect 123852 94522 123904 94528
rect 124416 89706 124444 96591
rect 124324 89678 124444 89706
rect 124324 86970 124352 89678
rect 124312 86964 124364 86970
rect 124312 86906 124364 86912
rect 124220 77308 124272 77314
rect 124220 77250 124272 77256
rect 122932 71052 122984 71058
rect 122932 70994 122984 71000
rect 124232 70378 124260 77250
rect 124220 70372 124272 70378
rect 124220 70314 124272 70320
rect 124404 70372 124456 70378
rect 124404 70314 124456 70320
rect 124416 60858 124444 70314
rect 124404 60852 124456 60858
rect 124404 60794 124456 60800
rect 124312 57996 124364 58002
rect 124312 57938 124364 57944
rect 124324 51134 124352 57938
rect 124312 51128 124364 51134
rect 124312 51070 124364 51076
rect 124128 49020 124180 49026
rect 124128 48962 124180 48968
rect 122840 11756 122892 11762
rect 122840 11698 122892 11704
rect 121828 4004 121880 4010
rect 121828 3946 121880 3952
rect 119436 3392 119488 3398
rect 119436 3334 119488 3340
rect 119988 3392 120040 3398
rect 119988 3334 120040 3340
rect 120632 3392 120684 3398
rect 120632 3334 120684 3340
rect 121368 3392 121420 3398
rect 121368 3334 121420 3340
rect 119448 480 119476 3334
rect 120644 480 120672 3334
rect 121840 480 121868 3946
rect 124140 3398 124168 48962
rect 124312 48340 124364 48346
rect 124312 48282 124364 48288
rect 124324 48226 124352 48282
rect 124232 48198 124352 48226
rect 124232 32434 124260 48198
rect 124220 32428 124272 32434
rect 124220 32370 124272 32376
rect 124876 4826 124904 100030
rect 124968 96665 124996 102068
rect 125704 102054 125902 102082
rect 126440 102054 126730 102082
rect 126992 102054 127558 102082
rect 124954 96656 125010 96665
rect 124954 96591 125010 96600
rect 125600 94580 125652 94586
rect 125600 94522 125652 94528
rect 125508 55888 125560 55894
rect 125508 55830 125560 55836
rect 124864 4820 124916 4826
rect 124864 4762 124916 4768
rect 125416 4072 125468 4078
rect 125416 4014 125468 4020
rect 123024 3392 123076 3398
rect 123024 3334 123076 3340
rect 124128 3392 124180 3398
rect 124128 3334 124180 3340
rect 124220 3392 124272 3398
rect 124220 3334 124272 3340
rect 123036 480 123064 3334
rect 124232 480 124260 3334
rect 125428 480 125456 4014
rect 125520 3398 125548 55830
rect 125612 13122 125640 94522
rect 125704 69698 125732 102054
rect 126440 94586 126468 102054
rect 126428 94580 126480 94586
rect 126428 94522 126480 94528
rect 126992 83502 127020 102054
rect 126980 83496 127032 83502
rect 126980 83438 127032 83444
rect 125692 69692 125744 69698
rect 125692 69634 125744 69640
rect 128464 39370 128492 102068
rect 129292 100026 129320 102068
rect 129280 100020 129332 100026
rect 129280 99962 129332 99968
rect 130120 99414 130148 102068
rect 130488 102054 130962 102082
rect 131132 102054 131882 102082
rect 132604 102054 132710 102082
rect 133248 102054 133538 102082
rect 129004 99408 129056 99414
rect 129004 99350 129056 99356
rect 130108 99408 130160 99414
rect 130108 99350 130160 99356
rect 129016 82142 129044 99350
rect 130488 89842 130516 102054
rect 130396 89814 130516 89842
rect 130396 89758 130424 89814
rect 129740 89752 129792 89758
rect 130384 89752 130436 89758
rect 129792 89700 129964 89706
rect 129740 89694 129964 89700
rect 130384 89694 130436 89700
rect 129752 89678 129964 89694
rect 129936 86970 129964 89678
rect 129924 86964 129976 86970
rect 129924 86906 129976 86912
rect 129004 82136 129056 82142
rect 129004 82078 129056 82084
rect 129832 77308 129884 77314
rect 129832 77250 129884 77256
rect 129844 70394 129872 77250
rect 129844 70366 130056 70394
rect 130028 68338 130056 70366
rect 130016 68332 130068 68338
rect 130016 68274 130068 68280
rect 128452 39364 128504 39370
rect 128452 39306 128504 39312
rect 131132 26926 131160 102054
rect 131764 100020 131816 100026
rect 131764 99962 131816 99968
rect 131120 26920 131172 26926
rect 131120 26862 131172 26868
rect 129648 25560 129700 25566
rect 129648 25502 129700 25508
rect 128268 21480 128320 21486
rect 128268 21422 128320 21428
rect 125600 13116 125652 13122
rect 125600 13058 125652 13064
rect 126612 4820 126664 4826
rect 126612 4762 126664 4768
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 126624 480 126652 4762
rect 128280 3398 128308 21422
rect 129660 3398 129688 25502
rect 131776 15910 131804 99962
rect 132500 94580 132552 94586
rect 132500 94522 132552 94528
rect 132408 26920 132460 26926
rect 132408 26862 132460 26868
rect 131764 15904 131816 15910
rect 131764 15846 131816 15852
rect 130200 9036 130252 9042
rect 130200 8978 130252 8984
rect 127808 3392 127860 3398
rect 127808 3334 127860 3340
rect 128268 3392 128320 3398
rect 128268 3334 128320 3340
rect 129004 3392 129056 3398
rect 129004 3334 129056 3340
rect 129648 3392 129700 3398
rect 129648 3334 129700 3340
rect 127820 480 127848 3334
rect 129016 480 129044 3334
rect 130212 480 130240 8978
rect 132420 3398 132448 26862
rect 132512 7614 132540 94522
rect 132604 80714 132632 102054
rect 133248 94586 133276 102054
rect 134352 95946 134380 102068
rect 134340 95940 134392 95946
rect 134340 95882 134392 95888
rect 135272 94738 135300 102068
rect 135824 102054 136114 102082
rect 135272 94710 135392 94738
rect 133236 94580 133288 94586
rect 133236 94522 133288 94528
rect 135260 94580 135312 94586
rect 135260 94522 135312 94528
rect 132592 80708 132644 80714
rect 132592 80650 132644 80656
rect 135272 57254 135300 94522
rect 135364 77994 135392 94710
rect 135824 94586 135852 102054
rect 136928 100026 136956 102068
rect 137296 102054 137862 102082
rect 138032 102054 138690 102082
rect 136916 100020 136968 100026
rect 136916 99962 136968 99968
rect 135812 94580 135864 94586
rect 135812 94522 135864 94528
rect 137296 89842 137324 102054
rect 137112 89814 137324 89842
rect 137112 89706 137140 89814
rect 136836 89678 137140 89706
rect 136836 80186 136864 89678
rect 136836 80158 136956 80186
rect 135352 77988 135404 77994
rect 135352 77930 135404 77936
rect 136928 77466 136956 80158
rect 136836 77438 136956 77466
rect 136836 77330 136864 77438
rect 136744 77302 136864 77330
rect 136744 77246 136772 77302
rect 136732 77240 136784 77246
rect 136732 77182 136784 77188
rect 136824 67652 136876 67658
rect 136824 67594 136876 67600
rect 136836 60738 136864 67594
rect 136836 60710 136956 60738
rect 136928 57934 136956 60710
rect 136916 57928 136968 57934
rect 136916 57870 136968 57876
rect 135260 57248 135312 57254
rect 135260 57190 135312 57196
rect 136824 48340 136876 48346
rect 136824 48282 136876 48288
rect 136836 41426 136864 48282
rect 136836 41398 136956 41426
rect 136548 39364 136600 39370
rect 136548 39306 136600 39312
rect 133788 10328 133840 10334
rect 133788 10270 133840 10276
rect 132500 7608 132552 7614
rect 132500 7550 132552 7556
rect 132592 6248 132644 6254
rect 132592 6190 132644 6196
rect 131396 3392 131448 3398
rect 131396 3334 131448 3340
rect 132408 3392 132460 3398
rect 132408 3334 132460 3340
rect 131408 480 131436 3334
rect 132604 480 132632 6190
rect 133800 480 133828 10270
rect 134892 7608 134944 7614
rect 134892 7550 134944 7556
rect 134904 480 134932 7550
rect 136560 3398 136588 39306
rect 136928 33794 136956 41398
rect 136916 33788 136968 33794
rect 136916 33730 136968 33736
rect 137928 11756 137980 11762
rect 137928 11698 137980 11704
rect 137940 3398 137968 11698
rect 138032 8974 138060 102054
rect 139400 94580 139452 94586
rect 139400 94522 139452 94528
rect 139308 90364 139360 90370
rect 139308 90306 139360 90312
rect 138020 8968 138072 8974
rect 138020 8910 138072 8916
rect 139320 3398 139348 90306
rect 139412 35222 139440 94522
rect 139504 40730 139532 102068
rect 140056 102054 140346 102082
rect 140884 102054 141266 102082
rect 141712 102054 142094 102082
rect 140056 94586 140084 102054
rect 140044 94580 140096 94586
rect 140044 94522 140096 94528
rect 140780 94580 140832 94586
rect 140780 94522 140832 94528
rect 139492 40724 139544 40730
rect 139492 40666 139544 40672
rect 140688 40724 140740 40730
rect 140688 40666 140740 40672
rect 139400 35216 139452 35222
rect 139400 35158 139452 35164
rect 140700 3398 140728 40666
rect 140792 29646 140820 94522
rect 140884 58682 140912 102054
rect 141712 94586 141740 102054
rect 142804 100020 142856 100026
rect 142804 99962 142856 99968
rect 142342 96656 142398 96665
rect 142342 96591 142398 96600
rect 141700 94580 141752 94586
rect 141700 94522 141752 94528
rect 142356 89706 142384 96591
rect 142264 89678 142384 89706
rect 142264 86970 142292 89678
rect 142252 86964 142304 86970
rect 142252 86906 142304 86912
rect 142160 77308 142212 77314
rect 142160 77250 142212 77256
rect 142172 77178 142200 77250
rect 142160 77172 142212 77178
rect 142160 77114 142212 77120
rect 142252 70372 142304 70378
rect 142252 70314 142304 70320
rect 140872 58676 140924 58682
rect 140872 58618 140924 58624
rect 142264 51082 142292 70314
rect 142264 51054 142384 51082
rect 142356 42090 142384 51054
rect 142344 42084 142396 42090
rect 142344 42026 142396 42032
rect 140780 29640 140832 29646
rect 140780 29582 140832 29588
rect 142068 28280 142120 28286
rect 142068 28222 142120 28228
rect 141976 13116 142028 13122
rect 141976 13058 142028 13064
rect 141988 3398 142016 13058
rect 136088 3392 136140 3398
rect 136088 3334 136140 3340
rect 136548 3392 136600 3398
rect 136548 3334 136600 3340
rect 137284 3392 137336 3398
rect 137284 3334 137336 3340
rect 137928 3392 137980 3398
rect 137928 3334 137980 3340
rect 138480 3392 138532 3398
rect 138480 3334 138532 3340
rect 139308 3392 139360 3398
rect 139308 3334 139360 3340
rect 139676 3392 139728 3398
rect 139676 3334 139728 3340
rect 140688 3392 140740 3398
rect 140688 3334 140740 3340
rect 140872 3392 140924 3398
rect 140872 3334 140924 3340
rect 141976 3392 142028 3398
rect 141976 3334 142028 3340
rect 136100 480 136128 3334
rect 137296 480 137324 3334
rect 138492 480 138520 3334
rect 139688 480 139716 3334
rect 140884 480 140912 3334
rect 142080 480 142108 28222
rect 142816 6254 142844 99962
rect 142908 96665 142936 102068
rect 143552 102054 143842 102082
rect 144104 102054 144670 102082
rect 144932 102054 145498 102082
rect 142894 96656 142950 96665
rect 142894 96591 142950 96600
rect 143448 42084 143500 42090
rect 143448 42026 143500 42032
rect 142804 6248 142856 6254
rect 142804 6190 142856 6196
rect 143460 3380 143488 42026
rect 143552 21418 143580 102054
rect 144104 91798 144132 102054
rect 144092 91792 144144 91798
rect 144092 91734 144144 91740
rect 144932 44878 144960 102054
rect 146312 94738 146340 102068
rect 146864 102054 147246 102082
rect 147784 102054 148074 102082
rect 148336 102054 148902 102082
rect 149072 102054 149730 102082
rect 150544 102054 150650 102082
rect 151096 102054 151478 102082
rect 151832 102054 152306 102082
rect 146312 94710 146432 94738
rect 146300 94580 146352 94586
rect 146300 94522 146352 94528
rect 144920 44872 144972 44878
rect 144920 44814 144972 44820
rect 146312 43450 146340 94522
rect 146404 60042 146432 94710
rect 146864 94586 146892 102054
rect 146852 94580 146904 94586
rect 146852 94522 146904 94528
rect 147680 80096 147732 80102
rect 147680 80038 147732 80044
rect 147692 75290 147720 80038
rect 147784 79354 147812 102054
rect 148336 89842 148364 102054
rect 147968 89814 148364 89842
rect 147968 80186 147996 89814
rect 147876 80158 147996 80186
rect 147876 80102 147904 80158
rect 147864 80096 147916 80102
rect 147864 80038 147916 80044
rect 147772 79348 147824 79354
rect 147772 79290 147824 79296
rect 147692 75262 147812 75290
rect 147784 70258 147812 75262
rect 147784 70230 147904 70258
rect 147876 60722 147904 70230
rect 147864 60716 147916 60722
rect 147864 60658 147916 60664
rect 147956 60648 148008 60654
rect 147956 60590 148008 60596
rect 146392 60036 146444 60042
rect 146392 59978 146444 59984
rect 146300 43444 146352 43450
rect 146300 43386 146352 43392
rect 147588 43444 147640 43450
rect 147588 43386 147640 43392
rect 146208 29640 146260 29646
rect 146208 29582 146260 29588
rect 143540 21412 143592 21418
rect 143540 21354 143592 21360
rect 144828 14476 144880 14482
rect 144828 14418 144880 14424
rect 144840 3380 144868 14418
rect 146220 3534 146248 29582
rect 147600 3534 147628 43386
rect 147968 41478 147996 60590
rect 147956 41472 148008 41478
rect 147956 41414 148008 41420
rect 147956 38684 148008 38690
rect 147956 38626 148008 38632
rect 147968 21978 147996 38626
rect 147968 21950 148088 21978
rect 145656 3528 145708 3534
rect 145656 3470 145708 3476
rect 146208 3528 146260 3534
rect 146208 3470 146260 3476
rect 146852 3528 146904 3534
rect 146852 3470 146904 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 143276 3352 143488 3380
rect 144472 3352 144868 3380
rect 143276 480 143304 3352
rect 144472 480 144500 3352
rect 145668 480 145696 3470
rect 146864 480 146892 3470
rect 148060 3398 148088 21950
rect 149072 17270 149100 102054
rect 150440 94580 150492 94586
rect 150440 94522 150492 94528
rect 150348 31068 150400 31074
rect 150348 31010 150400 31016
rect 149060 17264 149112 17270
rect 149060 17206 149112 17212
rect 148968 15904 149020 15910
rect 148968 15846 149020 15852
rect 148048 3392 148100 3398
rect 148048 3334 148100 3340
rect 148980 3194 149008 15846
rect 150360 4146 150388 31010
rect 149244 4140 149296 4146
rect 149244 4082 149296 4088
rect 150348 4140 150400 4146
rect 150348 4082 150400 4088
rect 148048 3188 148100 3194
rect 148048 3130 148100 3136
rect 148968 3188 149020 3194
rect 148968 3130 149020 3136
rect 148060 480 148088 3130
rect 149256 480 149284 4082
rect 150452 3618 150480 94522
rect 150544 46238 150572 102054
rect 151096 94586 151124 102054
rect 151084 94580 151136 94586
rect 151084 94522 151136 94528
rect 150532 46232 150584 46238
rect 150532 46174 150584 46180
rect 151728 44872 151780 44878
rect 151728 44814 151780 44820
rect 151636 17264 151688 17270
rect 151636 17206 151688 17212
rect 151648 9654 151676 17206
rect 151636 9648 151688 9654
rect 151636 9590 151688 9596
rect 150360 3602 150480 3618
rect 150348 3596 150480 3602
rect 150400 3590 150480 3596
rect 150348 3538 150400 3544
rect 151740 3534 151768 44814
rect 151832 18630 151860 102054
rect 153212 100094 153240 102068
rect 153200 100088 153252 100094
rect 153200 100030 153252 100036
rect 154040 96665 154068 102068
rect 154592 102054 154882 102082
rect 155144 102054 155710 102082
rect 155972 102054 156630 102082
rect 153382 96656 153438 96665
rect 153382 96591 153438 96600
rect 154026 96656 154082 96665
rect 154026 96591 154082 96600
rect 153396 38758 153424 96591
rect 154488 46232 154540 46238
rect 154488 46174 154540 46180
rect 153384 38752 153436 38758
rect 153384 38694 153436 38700
rect 153476 38752 153528 38758
rect 153476 38694 153528 38700
rect 153108 32428 153160 32434
rect 153108 32370 153160 32376
rect 151820 18624 151872 18630
rect 151820 18566 151872 18572
rect 150440 3528 150492 3534
rect 150440 3470 150492 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 150452 480 150480 3470
rect 153120 626 153148 32370
rect 153488 31822 153516 38694
rect 153476 31816 153528 31822
rect 153476 31758 153528 31764
rect 153384 29096 153436 29102
rect 153304 29044 153384 29050
rect 153304 29038 153436 29044
rect 153304 29022 153424 29038
rect 153304 27606 153332 29022
rect 153292 27600 153344 27606
rect 153292 27542 153344 27548
rect 153384 18012 153436 18018
rect 153384 17954 153436 17960
rect 153396 9602 153424 17954
rect 153396 9574 153516 9602
rect 153488 3466 153516 9574
rect 154500 4146 154528 46174
rect 154592 19990 154620 102054
rect 155144 89842 155172 102054
rect 154960 89814 155172 89842
rect 154960 80782 154988 89814
rect 154948 80776 155000 80782
rect 154948 80718 155000 80724
rect 154764 67652 154816 67658
rect 154764 67594 154816 67600
rect 154776 47598 154804 67594
rect 154764 47592 154816 47598
rect 154764 47534 154816 47540
rect 154580 19984 154632 19990
rect 154580 19926 154632 19932
rect 155868 18624 155920 18630
rect 155868 18566 155920 18572
rect 153936 4140 153988 4146
rect 153936 4082 153988 4088
rect 154488 4140 154540 4146
rect 154488 4082 154540 4088
rect 153476 3460 153528 3466
rect 153476 3402 153528 3408
rect 151544 604 151596 610
rect 151544 546 151596 552
rect 152752 598 153148 626
rect 151556 480 151584 546
rect 152752 480 152780 598
rect 153948 480 153976 4082
rect 155880 3194 155908 18566
rect 155972 3670 156000 102054
rect 157444 99414 157472 102068
rect 157628 102054 158286 102082
rect 158732 102054 159206 102082
rect 159652 102054 160034 102082
rect 156604 99408 156656 99414
rect 156604 99350 156656 99356
rect 157432 99408 157484 99414
rect 157432 99350 157484 99356
rect 156616 24138 156644 99350
rect 157628 89842 157656 102054
rect 157984 100700 158036 100706
rect 157984 100642 158036 100648
rect 157536 89814 157656 89842
rect 157536 60790 157564 89814
rect 157524 60784 157576 60790
rect 157524 60726 157576 60732
rect 157340 60716 157392 60722
rect 157340 60658 157392 60664
rect 157352 50386 157380 60658
rect 157340 50380 157392 50386
rect 157340 50322 157392 50328
rect 157248 33788 157300 33794
rect 157248 33730 157300 33736
rect 156604 24132 156656 24138
rect 156604 24074 156656 24080
rect 155960 3664 156012 3670
rect 155960 3606 156012 3612
rect 155132 3188 155184 3194
rect 155132 3130 155184 3136
rect 155868 3188 155920 3194
rect 155868 3130 155920 3136
rect 155144 480 155172 3130
rect 157260 2922 157288 33730
rect 157996 14550 158024 100642
rect 158628 47592 158680 47598
rect 158628 47534 158680 47540
rect 157984 14544 158036 14550
rect 157984 14486 158036 14492
rect 158640 3874 158668 47534
rect 158732 4298 158760 102054
rect 159652 89758 159680 102054
rect 160848 99414 160876 102068
rect 161492 102054 161690 102082
rect 162136 102054 162610 102082
rect 162872 102054 163438 102082
rect 160100 99408 160152 99414
rect 160100 99350 160152 99356
rect 160836 99408 160888 99414
rect 160836 99350 160888 99356
rect 160112 89758 160140 99350
rect 158904 89752 158956 89758
rect 158904 89694 158956 89700
rect 159640 89752 159692 89758
rect 159640 89694 159692 89700
rect 160100 89752 160152 89758
rect 160100 89694 160152 89700
rect 158916 80186 158944 89694
rect 160192 89616 160244 89622
rect 160192 89558 160244 89564
rect 160204 85542 160232 89558
rect 160192 85536 160244 85542
rect 160192 85478 160244 85484
rect 158824 80158 158944 80186
rect 158824 70446 158852 80158
rect 160192 75948 160244 75954
rect 160192 75890 160244 75896
rect 158812 70440 158864 70446
rect 158812 70382 158864 70388
rect 158904 70304 158956 70310
rect 158904 70246 158956 70252
rect 158916 41426 158944 70246
rect 160204 67590 160232 75890
rect 160192 67584 160244 67590
rect 160192 67526 160244 67532
rect 160192 57996 160244 58002
rect 160192 57938 160244 57944
rect 160204 51746 160232 57938
rect 161388 57248 161440 57254
rect 161388 57190 161440 57196
rect 160192 51740 160244 51746
rect 160192 51682 160244 51688
rect 158824 41398 158944 41426
rect 158824 38622 158852 41398
rect 158812 38616 158864 38622
rect 158812 38558 158864 38564
rect 160008 35216 160060 35222
rect 160008 35158 160060 35164
rect 158996 29028 159048 29034
rect 158996 28970 159048 28976
rect 159008 28914 159036 28970
rect 159008 28886 159128 28914
rect 159100 22778 159128 28886
rect 159088 22772 159140 22778
rect 159088 22714 159140 22720
rect 159916 19984 159968 19990
rect 159916 19926 159968 19932
rect 158732 4270 158852 4298
rect 158720 4140 158772 4146
rect 158720 4082 158772 4088
rect 157524 3868 157576 3874
rect 157524 3810 157576 3816
rect 158628 3868 158680 3874
rect 158628 3810 158680 3816
rect 156328 2916 156380 2922
rect 156328 2858 156380 2864
rect 157248 2916 157300 2922
rect 157248 2858 157300 2864
rect 156340 480 156368 2858
rect 157536 480 157564 3810
rect 158732 480 158760 4082
rect 158824 3738 158852 4270
rect 159928 4146 159956 19926
rect 159916 4140 159968 4146
rect 159916 4082 159968 4088
rect 160020 4026 160048 35158
rect 159928 3998 160048 4026
rect 158812 3732 158864 3738
rect 158812 3674 158864 3680
rect 159928 480 159956 3998
rect 161400 610 161428 57190
rect 161492 3806 161520 102054
rect 162136 89842 162164 102054
rect 161768 89814 162164 89842
rect 161768 80170 161796 89814
rect 161756 80164 161808 80170
rect 161756 80106 161808 80112
rect 161664 80096 161716 80102
rect 161664 80038 161716 80044
rect 161676 70514 161704 80038
rect 161664 70508 161716 70514
rect 161664 70450 161716 70456
rect 161664 70236 161716 70242
rect 161664 70178 161716 70184
rect 161676 41426 161704 70178
rect 162872 53106 162900 102054
rect 162860 53100 162912 53106
rect 162860 53042 162912 53048
rect 161584 41398 161704 41426
rect 161584 35578 161612 41398
rect 161584 35550 161704 35578
rect 161676 28966 161704 35550
rect 161664 28960 161716 28966
rect 161664 28902 161716 28908
rect 164148 22772 164200 22778
rect 164148 22714 164200 22720
rect 161848 19372 161900 19378
rect 161848 19314 161900 19320
rect 161860 6186 161888 19314
rect 161848 6180 161900 6186
rect 161848 6122 161900 6128
rect 162308 6180 162360 6186
rect 162308 6122 162360 6128
rect 161480 3800 161532 3806
rect 161480 3742 161532 3748
rect 161112 604 161164 610
rect 161112 546 161164 552
rect 161388 604 161440 610
rect 161388 546 161440 552
rect 161124 480 161152 546
rect 162320 480 162348 6122
rect 164160 4146 164188 22714
rect 163504 4140 163556 4146
rect 163504 4082 163556 4088
rect 164148 4140 164200 4146
rect 164148 4082 164200 4088
rect 163516 480 163544 4082
rect 164252 3942 164280 102068
rect 165172 95266 165200 102068
rect 166000 100706 166028 102068
rect 166368 102054 166842 102082
rect 167012 102054 167670 102082
rect 168484 102054 168590 102082
rect 169128 102054 169418 102082
rect 169772 102054 170246 102082
rect 170508 102054 171074 102082
rect 171244 102054 171994 102082
rect 172532 102054 172822 102082
rect 173176 102054 173650 102082
rect 173912 102054 174570 102082
rect 175292 102054 175398 102082
rect 165988 100700 166040 100706
rect 165988 100642 166040 100648
rect 164424 95260 164476 95266
rect 164424 95202 164476 95208
rect 165160 95260 165212 95266
rect 165160 95202 165212 95208
rect 164436 85542 164464 95202
rect 166368 89758 166396 102054
rect 165712 89752 165764 89758
rect 165712 89694 165764 89700
rect 166356 89752 166408 89758
rect 166356 89694 166408 89700
rect 164424 85536 164476 85542
rect 164424 85478 164476 85484
rect 164424 75948 164476 75954
rect 164424 75890 164476 75896
rect 164436 72486 164464 75890
rect 164424 72480 164476 72486
rect 164424 72422 164476 72428
rect 164332 67652 164384 67658
rect 164332 67594 164384 67600
rect 164344 67561 164372 67594
rect 164330 67552 164386 67561
rect 164330 67487 164386 67496
rect 164422 67416 164478 67425
rect 164422 67351 164478 67360
rect 164436 41426 164464 67351
rect 164344 41398 164464 41426
rect 164344 36582 164372 41398
rect 165724 41290 165752 89694
rect 165724 41262 165844 41290
rect 164332 36576 164384 36582
rect 164332 36518 164384 36524
rect 165528 36576 165580 36582
rect 165528 36518 165580 36524
rect 164240 3936 164292 3942
rect 164240 3878 164292 3884
rect 165540 3534 165568 36518
rect 165816 22166 165844 41262
rect 167012 37942 167040 102054
rect 167644 100088 167696 100094
rect 167644 100030 167696 100036
rect 167000 37936 167052 37942
rect 167000 37878 167052 37884
rect 165804 22160 165856 22166
rect 165804 22102 165856 22108
rect 165712 22092 165764 22098
rect 165712 22034 165764 22040
rect 165724 12458 165752 22034
rect 165724 12430 165844 12458
rect 165816 3670 165844 12430
rect 167656 4894 167684 100030
rect 168380 94580 168432 94586
rect 168380 94522 168432 94528
rect 168288 37936 168340 37942
rect 168288 37878 168340 37884
rect 168196 24132 168248 24138
rect 168196 24074 168248 24080
rect 165896 4888 165948 4894
rect 165896 4830 165948 4836
rect 167644 4888 167696 4894
rect 167644 4830 167696 4836
rect 165804 3664 165856 3670
rect 165804 3606 165856 3612
rect 164700 3528 164752 3534
rect 164700 3470 164752 3476
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 164712 480 164740 3470
rect 165908 480 165936 4830
rect 168208 4146 168236 24074
rect 167092 4140 167144 4146
rect 167092 4082 167144 4088
rect 168196 4140 168248 4146
rect 168196 4082 168248 4088
rect 167104 480 167132 4082
rect 168300 4026 168328 37878
rect 168392 4078 168420 94522
rect 168484 54534 168512 102054
rect 169128 94586 169156 102054
rect 169116 94580 169168 94586
rect 169116 94522 169168 94528
rect 168472 54528 168524 54534
rect 168472 54470 168524 54476
rect 169772 49026 169800 102054
rect 170508 89842 170536 102054
rect 171244 89842 171272 102054
rect 170416 89814 170536 89842
rect 171152 89814 171272 89842
rect 170416 89758 170444 89814
rect 169944 89752 169996 89758
rect 169944 89694 169996 89700
rect 170404 89752 170456 89758
rect 170404 89694 170456 89700
rect 169956 85542 169984 89694
rect 169944 85536 169996 85542
rect 169944 85478 169996 85484
rect 169944 75948 169996 75954
rect 169944 75890 169996 75896
rect 169956 70446 169984 75890
rect 169944 70440 169996 70446
rect 169944 70382 169996 70388
rect 170036 70304 170088 70310
rect 170036 70246 170088 70252
rect 170048 67590 170076 70246
rect 169852 67584 169904 67590
rect 169852 67526 169904 67532
rect 170036 67584 170088 67590
rect 170036 67526 170088 67532
rect 169864 55894 169892 67526
rect 169852 55888 169904 55894
rect 169852 55830 169904 55836
rect 169760 49020 169812 49026
rect 169760 48962 169812 48968
rect 171152 28966 171180 89814
rect 171140 28960 171192 28966
rect 171140 28902 171192 28908
rect 171048 21412 171100 21418
rect 171048 21354 171100 21360
rect 169392 7676 169444 7682
rect 169392 7618 169444 7624
rect 168208 3998 168328 4026
rect 168380 4072 168432 4078
rect 168380 4014 168432 4020
rect 168208 480 168236 3998
rect 169404 480 169432 7618
rect 171060 4146 171088 21354
rect 171324 19372 171376 19378
rect 171324 19314 171376 19320
rect 170588 4140 170640 4146
rect 170588 4082 170640 4088
rect 171048 4140 171100 4146
rect 171048 4082 171100 4088
rect 170600 480 170628 4082
rect 171336 3942 171364 19314
rect 172532 4826 172560 102054
rect 173176 96626 173204 102054
rect 173164 96620 173216 96626
rect 173164 96562 173216 96568
rect 172888 89684 172940 89690
rect 172888 89626 172940 89632
rect 172900 80782 172928 89626
rect 172888 80776 172940 80782
rect 172888 80718 172940 80724
rect 172612 75948 172664 75954
rect 172612 75890 172664 75896
rect 172624 70394 172652 75890
rect 172624 70366 172836 70394
rect 172808 60790 172836 70366
rect 172796 60784 172848 60790
rect 172796 60726 172848 60732
rect 172888 60716 172940 60722
rect 172888 60658 172940 60664
rect 172900 57934 172928 60658
rect 172888 57928 172940 57934
rect 172888 57870 172940 57876
rect 172612 46980 172664 46986
rect 172612 46922 172664 46928
rect 172624 41478 172652 46922
rect 172612 41472 172664 41478
rect 172612 41414 172664 41420
rect 172704 41336 172756 41342
rect 172704 41278 172756 41284
rect 172716 29102 172744 41278
rect 172704 29096 172756 29102
rect 172704 29038 172756 29044
rect 172612 29028 172664 29034
rect 172612 28970 172664 28976
rect 172624 21486 172652 28970
rect 173912 25566 173940 102054
rect 173900 25560 173952 25566
rect 173900 25502 173952 25508
rect 175188 25560 175240 25566
rect 175188 25502 175240 25508
rect 172612 21480 172664 21486
rect 172612 21422 172664 21428
rect 172520 4820 172572 4826
rect 172520 4762 172572 4768
rect 172980 4820 173032 4826
rect 172980 4762 173032 4768
rect 171324 3936 171376 3942
rect 171324 3878 171376 3884
rect 171784 3460 171836 3466
rect 171784 3402 171836 3408
rect 171796 480 171824 3402
rect 172992 480 173020 4762
rect 175200 4146 175228 25502
rect 175292 9042 175320 102054
rect 175568 89826 175596 102190
rect 177040 100026 177068 102068
rect 177316 102054 177974 102082
rect 178420 102054 178802 102082
rect 179524 102054 179630 102082
rect 180168 102054 180550 102082
rect 180812 102054 181378 102082
rect 177028 100020 177080 100026
rect 177028 99962 177080 99968
rect 177316 89842 177344 102054
rect 178420 96626 178448 102054
rect 178684 100020 178736 100026
rect 178684 99962 178736 99968
rect 178408 96620 178460 96626
rect 178408 96562 178460 96568
rect 175556 89820 175608 89826
rect 175556 89762 175608 89768
rect 177224 89814 177344 89842
rect 175464 89752 175516 89758
rect 175464 89694 175516 89700
rect 175476 70446 175504 89694
rect 177224 80186 177252 89814
rect 178132 87100 178184 87106
rect 178132 87042 178184 87048
rect 178144 85542 178172 87042
rect 178132 85536 178184 85542
rect 178132 85478 178184 85484
rect 177132 80158 177252 80186
rect 176672 80102 176700 80133
rect 177132 80102 177160 80158
rect 176660 80096 176712 80102
rect 177120 80096 177172 80102
rect 176712 80044 176884 80050
rect 176660 80038 176884 80044
rect 177120 80038 177172 80044
rect 176672 80022 176884 80038
rect 175464 70440 175516 70446
rect 175464 70382 175516 70388
rect 175556 70304 175608 70310
rect 175556 70246 175608 70252
rect 175568 60738 175596 70246
rect 176856 69902 176884 80022
rect 178408 75948 178460 75954
rect 178408 75890 178460 75896
rect 176844 69896 176896 69902
rect 176844 69838 176896 69844
rect 176844 69760 176896 69766
rect 176844 69702 176896 69708
rect 176856 60858 176884 69702
rect 178420 67726 178448 75890
rect 178132 67720 178184 67726
rect 178132 67662 178184 67668
rect 178408 67720 178460 67726
rect 178408 67662 178460 67668
rect 178144 66230 178172 67662
rect 178132 66224 178184 66230
rect 178132 66166 178184 66172
rect 176844 60852 176896 60858
rect 176844 60794 176896 60800
rect 175384 60722 175596 60738
rect 176752 60784 176804 60790
rect 176752 60726 176804 60732
rect 175372 60716 175608 60722
rect 175424 60710 175556 60716
rect 175372 60658 175424 60664
rect 175556 60658 175608 60664
rect 175568 51134 175596 60658
rect 176764 53122 176792 60726
rect 178408 56636 178460 56642
rect 178408 56578 178460 56584
rect 176672 53094 176792 53122
rect 175556 51128 175608 51134
rect 175556 51070 175608 51076
rect 175372 51060 175424 51066
rect 175372 51002 175424 51008
rect 175384 48249 175412 51002
rect 176672 48346 176700 53094
rect 178420 48346 178448 56578
rect 176660 48340 176712 48346
rect 176660 48282 176712 48288
rect 176936 48340 176988 48346
rect 176936 48282 176988 48288
rect 178132 48340 178184 48346
rect 178132 48282 178184 48288
rect 178408 48340 178460 48346
rect 178408 48282 178460 48288
rect 175370 48240 175426 48249
rect 175370 48175 175426 48184
rect 175462 48104 175518 48113
rect 175462 48039 175518 48048
rect 175476 26926 175504 48039
rect 176948 38758 176976 48282
rect 178144 44962 178172 48282
rect 178144 44934 178264 44962
rect 178236 38826 178264 44934
rect 178224 38820 178276 38826
rect 178224 38762 178276 38768
rect 176936 38752 176988 38758
rect 176936 38694 176988 38700
rect 176844 38684 176896 38690
rect 176844 38626 176896 38632
rect 178224 38684 178276 38690
rect 178224 38626 178276 38632
rect 176856 38570 176884 38626
rect 176764 38542 176884 38570
rect 176764 34678 176792 38542
rect 176752 34672 176804 34678
rect 176752 34614 176804 34620
rect 178236 33810 178264 38626
rect 178144 33782 178264 33810
rect 178144 31634 178172 33782
rect 178144 31606 178356 31634
rect 176936 27668 176988 27674
rect 176936 27610 176988 27616
rect 175464 26920 175516 26926
rect 175464 26862 175516 26868
rect 176948 22166 176976 27610
rect 177948 26920 178000 26926
rect 177948 26862 178000 26868
rect 176936 22160 176988 22166
rect 176936 22102 176988 22108
rect 176752 22092 176804 22098
rect 176752 22034 176804 22040
rect 176764 12510 176792 22034
rect 176752 12504 176804 12510
rect 176752 12446 176804 12452
rect 175280 9036 175332 9042
rect 175280 8978 175332 8984
rect 176568 8968 176620 8974
rect 176568 8910 176620 8916
rect 174176 4140 174228 4146
rect 174176 4082 174228 4088
rect 175188 4140 175240 4146
rect 175188 4082 175240 4088
rect 174188 480 174216 4082
rect 175372 3596 175424 3602
rect 175372 3538 175424 3544
rect 175384 480 175412 3538
rect 176580 480 176608 8910
rect 177960 2854 177988 26862
rect 178328 22114 178356 31606
rect 178696 28286 178724 99962
rect 179420 92404 179472 92410
rect 179420 92346 179472 92352
rect 178684 28280 178736 28286
rect 178684 28222 178736 28228
rect 178144 22086 178356 22114
rect 178144 21978 178172 22086
rect 178144 21950 178264 21978
rect 178236 7614 178264 21950
rect 179432 11762 179460 92346
rect 179524 39370 179552 102054
rect 180168 92410 180196 102054
rect 180156 92404 180208 92410
rect 180156 92346 180208 92352
rect 180812 90370 180840 102054
rect 182192 94738 182220 102068
rect 182744 102054 183034 102082
rect 182192 94710 182312 94738
rect 182180 94580 182232 94586
rect 182180 94522 182232 94528
rect 180800 90364 180852 90370
rect 180800 90306 180852 90312
rect 179512 39364 179564 39370
rect 179512 39306 179564 39312
rect 182088 28280 182140 28286
rect 182088 28222 182140 28228
rect 179420 11756 179472 11762
rect 179420 11698 179472 11704
rect 180156 10328 180208 10334
rect 180156 10270 180208 10276
rect 178224 7608 178276 7614
rect 178224 7550 178276 7556
rect 178960 3528 179012 3534
rect 178960 3470 179012 3476
rect 177948 2848 178000 2854
rect 177948 2790 178000 2796
rect 177764 604 177816 610
rect 177764 546 177816 552
rect 177776 480 177804 546
rect 178972 480 179000 3470
rect 180168 480 180196 10270
rect 182100 3262 182128 28222
rect 182192 13122 182220 94522
rect 182284 40730 182312 94710
rect 182744 94586 182772 102054
rect 183940 100026 183968 102068
rect 183928 100020 183980 100026
rect 183928 99962 183980 99968
rect 182732 94580 182784 94586
rect 182732 94522 182784 94528
rect 184124 89842 184152 102190
rect 184032 89814 184152 89842
rect 184952 102054 185610 102082
rect 186332 102054 186438 102082
rect 184032 86970 184060 89814
rect 184020 86964 184072 86970
rect 184020 86906 184072 86912
rect 183744 80028 183796 80034
rect 183744 79970 183796 79976
rect 183756 77246 183784 79970
rect 183744 77240 183796 77246
rect 183744 77182 183796 77188
rect 183744 66292 183796 66298
rect 183744 66234 183796 66240
rect 183756 58002 183784 66234
rect 183744 57996 183796 58002
rect 183744 57938 183796 57944
rect 183744 57860 183796 57866
rect 183744 57802 183796 57808
rect 183756 51134 183784 57802
rect 183744 51128 183796 51134
rect 183744 51070 183796 51076
rect 183744 50992 183796 50998
rect 183744 50934 183796 50940
rect 183756 42090 183784 50934
rect 183744 42084 183796 42090
rect 183744 42026 183796 42032
rect 182272 40724 182324 40730
rect 182272 40666 182324 40672
rect 184848 17332 184900 17338
rect 184848 17274 184900 17280
rect 182180 13116 182232 13122
rect 182180 13058 182232 13064
rect 183744 11756 183796 11762
rect 183744 11698 183796 11704
rect 182548 3664 182600 3670
rect 182548 3606 182600 3612
rect 181352 3256 181404 3262
rect 181352 3198 181404 3204
rect 182088 3256 182140 3262
rect 182088 3198 182140 3204
rect 181364 480 181392 3198
rect 182560 480 182588 3606
rect 183756 480 183784 11698
rect 184860 480 184888 17274
rect 184952 14482 184980 102054
rect 185584 99408 185636 99414
rect 185584 99350 185636 99356
rect 185596 15910 185624 99350
rect 186332 29646 186360 102054
rect 186608 98002 186636 102190
rect 188172 99414 188200 102068
rect 188160 99408 188212 99414
rect 188160 99350 188212 99356
rect 188356 98002 188384 102190
rect 189184 98002 189212 102190
rect 186424 97974 186636 98002
rect 187804 97974 188384 98002
rect 189092 97974 189212 98002
rect 190472 102054 190762 102082
rect 186424 43450 186452 97974
rect 186412 43444 186464 43450
rect 186412 43386 186464 43392
rect 187804 31074 187832 97974
rect 189092 44878 189120 97974
rect 189080 44872 189132 44878
rect 189080 44814 189132 44820
rect 187792 31068 187844 31074
rect 187792 31010 187844 31016
rect 186320 29640 186372 29646
rect 186320 29582 186372 29588
rect 188988 29640 189040 29646
rect 188988 29582 189040 29588
rect 185584 15904 185636 15910
rect 185584 15846 185636 15852
rect 184940 14476 184992 14482
rect 184940 14418 184992 14424
rect 187608 13116 187660 13122
rect 187608 13058 187660 13064
rect 186044 3732 186096 3738
rect 186044 3674 186096 3680
rect 186056 480 186084 3674
rect 187620 3482 187648 13058
rect 187252 3454 187648 3482
rect 187252 480 187280 3454
rect 189000 3398 189028 29582
rect 190472 17270 190500 102054
rect 190932 98002 190960 102190
rect 190564 97974 190960 98002
rect 191852 102054 192418 102082
rect 193232 102054 193338 102082
rect 190564 32434 190592 97974
rect 191852 46238 191880 102054
rect 191840 46232 191892 46238
rect 191840 46174 191892 46180
rect 190552 32428 190604 32434
rect 190552 32370 190604 32376
rect 193128 18692 193180 18698
rect 193128 18634 193180 18640
rect 190460 17264 190512 17270
rect 190460 17206 190512 17212
rect 191748 14476 191800 14482
rect 191748 14418 191800 14424
rect 189632 3800 189684 3806
rect 189632 3742 189684 3748
rect 188436 3392 188488 3398
rect 188436 3334 188488 3340
rect 188988 3392 189040 3398
rect 188988 3334 189040 3340
rect 188448 480 188476 3334
rect 189644 480 189672 3742
rect 191760 3398 191788 14418
rect 193140 3398 193168 18634
rect 193232 18630 193260 102054
rect 193508 98002 193536 102190
rect 193324 97974 193536 98002
rect 194704 102054 194994 102082
rect 195624 102054 195914 102082
rect 196360 102054 196742 102082
rect 197464 102054 197570 102082
rect 198016 102054 198398 102082
rect 198752 102054 199318 102082
rect 200040 102054 200146 102082
rect 194600 97980 194652 97986
rect 193324 33794 193352 97974
rect 194600 97922 194652 97928
rect 193312 33788 193364 33794
rect 193312 33730 193364 33736
rect 194612 19990 194640 97922
rect 194704 47598 194732 102054
rect 195624 97986 195652 102054
rect 195612 97980 195664 97986
rect 195612 97922 195664 97928
rect 196360 89842 196388 102054
rect 197360 94580 197412 94586
rect 197360 94522 197412 94528
rect 196176 89814 196388 89842
rect 196176 89706 196204 89814
rect 196084 89678 196204 89706
rect 196084 86970 196112 89678
rect 196072 86964 196124 86970
rect 196072 86906 196124 86912
rect 195980 77308 196032 77314
rect 195980 77250 196032 77256
rect 194692 47592 194744 47598
rect 194692 47534 194744 47540
rect 195992 35222 196020 77250
rect 195980 35216 196032 35222
rect 195980 35158 196032 35164
rect 194600 19984 194652 19990
rect 194600 19926 194652 19932
rect 195888 19984 195940 19990
rect 195888 19926 195940 19932
rect 193220 18624 193272 18630
rect 193220 18566 193272 18572
rect 194416 6248 194468 6254
rect 194416 6190 194468 6196
rect 193220 3936 193272 3942
rect 193220 3878 193272 3884
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 191748 3392 191800 3398
rect 191748 3334 191800 3340
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 190840 480 190868 3334
rect 192036 480 192064 3334
rect 193232 480 193260 3878
rect 194428 480 194456 6190
rect 195900 3482 195928 19926
rect 197372 6186 197400 94522
rect 197464 57254 197492 102054
rect 198016 94586 198044 102054
rect 198004 94580 198056 94586
rect 198004 94522 198056 94528
rect 197452 57248 197504 57254
rect 197452 57190 197504 57196
rect 198752 22778 198780 102054
rect 200040 96665 200068 102054
rect 200764 100428 200816 100434
rect 200764 100370 200816 100376
rect 200026 96656 200082 96665
rect 200026 96591 200082 96600
rect 200302 96656 200358 96665
rect 200302 96591 200358 96600
rect 200316 86970 200344 96591
rect 200304 86964 200356 86970
rect 200304 86906 200356 86912
rect 200304 77308 200356 77314
rect 200304 77250 200356 77256
rect 200316 36582 200344 77250
rect 200304 36576 200356 36582
rect 200304 36518 200356 36524
rect 200776 24138 200804 100370
rect 200960 100094 200988 102068
rect 201788 100434 201816 102068
rect 202064 102054 202722 102082
rect 202892 102054 203550 102082
rect 201776 100428 201828 100434
rect 201776 100370 201828 100376
rect 200948 100088 201000 100094
rect 200948 100030 201000 100036
rect 202064 94466 202092 102054
rect 201604 94438 202092 94466
rect 201604 37942 201632 94438
rect 201592 37936 201644 37942
rect 201592 37878 201644 37884
rect 200764 24132 200816 24138
rect 200764 24074 200816 24080
rect 202696 24132 202748 24138
rect 202696 24074 202748 24080
rect 198740 22772 198792 22778
rect 198740 22714 198792 22720
rect 200028 22772 200080 22778
rect 200028 22714 200080 22720
rect 198648 15904 198700 15910
rect 198648 15846 198700 15852
rect 197360 6180 197412 6186
rect 197360 6122 197412 6128
rect 196808 3868 196860 3874
rect 196808 3810 196860 3816
rect 195624 3454 195928 3482
rect 195624 480 195652 3454
rect 196820 480 196848 3810
rect 198660 3398 198688 15846
rect 200040 3398 200068 22714
rect 201500 4888 201552 4894
rect 201500 4830 201552 4836
rect 200396 4072 200448 4078
rect 200396 4014 200448 4020
rect 198004 3392 198056 3398
rect 198004 3334 198056 3340
rect 198648 3392 198700 3398
rect 198648 3334 198700 3340
rect 199200 3392 199252 3398
rect 199200 3334 199252 3340
rect 200028 3392 200080 3398
rect 200028 3334 200080 3340
rect 198016 480 198044 3334
rect 199212 480 199240 3334
rect 200408 480 200436 4014
rect 201512 480 201540 4830
rect 202708 480 202736 24074
rect 202892 7682 202920 102054
rect 203524 99408 203576 99414
rect 203524 99350 203576 99356
rect 202880 7676 202932 7682
rect 202880 7618 202932 7624
rect 203536 4826 203564 99350
rect 204364 21418 204392 102068
rect 204548 102054 205298 102082
rect 204548 89842 204576 102054
rect 206112 99414 206140 102068
rect 206100 99408 206152 99414
rect 206100 99350 206152 99356
rect 206940 96665 206968 102068
rect 207664 100020 207716 100026
rect 207664 99962 207716 99968
rect 206558 96656 206614 96665
rect 206558 96591 206614 96600
rect 206926 96656 206982 96665
rect 206926 96591 206982 96600
rect 207294 96656 207350 96665
rect 207294 96591 207350 96600
rect 204456 89814 204576 89842
rect 204352 21412 204404 21418
rect 204352 21354 204404 21360
rect 203524 4820 203576 4826
rect 203524 4762 203576 4768
rect 203892 4004 203944 4010
rect 203892 3946 203944 3952
rect 203904 480 203932 3946
rect 204456 3466 204484 89814
rect 206572 86986 206600 96591
rect 207308 86986 207336 96591
rect 206480 86958 206600 86986
rect 207216 86958 207336 86986
rect 206480 80238 206508 86958
rect 205732 80232 205784 80238
rect 205732 80174 205784 80180
rect 206468 80232 206520 80238
rect 206468 80174 206520 80180
rect 205744 72978 205772 80174
rect 207216 77353 207244 86958
rect 207018 77344 207074 77353
rect 207018 77279 207074 77288
rect 207202 77344 207258 77353
rect 207202 77279 207258 77288
rect 205744 72950 205956 72978
rect 205928 53122 205956 72950
rect 207032 71074 207060 77279
rect 207032 71046 207244 71074
rect 207216 53122 207244 71046
rect 205836 53094 205956 53122
rect 207124 53094 207244 53122
rect 205836 48278 205864 53094
rect 207124 48278 207152 53094
rect 205732 48272 205784 48278
rect 205732 48214 205784 48220
rect 205824 48272 205876 48278
rect 205824 48214 205876 48220
rect 206928 48272 206980 48278
rect 206928 48214 206980 48220
rect 207112 48272 207164 48278
rect 207112 48214 207164 48220
rect 205744 25566 205772 48214
rect 206940 38706 206968 48214
rect 206940 38678 207060 38706
rect 207032 38622 207060 38678
rect 207020 38616 207072 38622
rect 207020 38558 207072 38564
rect 207112 29028 207164 29034
rect 207112 28970 207164 28976
rect 205732 25560 205784 25566
rect 205732 25502 205784 25508
rect 206928 21412 206980 21418
rect 206928 21354 206980 21360
rect 205088 7608 205140 7614
rect 205088 7550 205140 7556
rect 204444 3460 204496 3466
rect 204444 3402 204496 3408
rect 205100 480 205128 7550
rect 206940 1154 206968 21354
rect 207124 19378 207152 28970
rect 207020 19372 207072 19378
rect 207020 19314 207072 19320
rect 207112 19372 207164 19378
rect 207112 19314 207164 19320
rect 207032 9602 207060 19314
rect 207676 15910 207704 99962
rect 207768 96665 207796 102068
rect 208412 102054 208702 102082
rect 207754 96656 207810 96665
rect 207754 96591 207810 96600
rect 207664 15904 207716 15910
rect 207664 15846 207716 15852
rect 207032 9574 207152 9602
rect 207124 3602 207152 9574
rect 208412 8974 208440 102054
rect 209516 96665 209544 102068
rect 209976 102054 210358 102082
rect 211172 102054 211278 102082
rect 208858 96656 208914 96665
rect 208676 96620 208728 96626
rect 208858 96591 208860 96600
rect 208676 96562 208728 96568
rect 208912 96591 208914 96600
rect 209502 96656 209558 96665
rect 209502 96591 209558 96600
rect 208860 96562 208912 96568
rect 208688 86986 208716 96562
rect 208504 86958 208716 86986
rect 208504 70446 208532 86958
rect 208492 70440 208544 70446
rect 208492 70382 208544 70388
rect 208584 70304 208636 70310
rect 208584 70246 208636 70252
rect 208596 60874 208624 70246
rect 208596 60846 208716 60874
rect 208688 56642 208716 60846
rect 208492 56636 208544 56642
rect 208492 56578 208544 56584
rect 208676 56636 208728 56642
rect 208676 56578 208728 56584
rect 208504 53122 208532 56578
rect 208504 53094 208716 53122
rect 208688 50946 208716 53094
rect 208596 50918 208716 50946
rect 208596 48278 208624 50918
rect 208584 48272 208636 48278
rect 208584 48214 208636 48220
rect 208492 38684 208544 38690
rect 208492 38626 208544 38632
rect 208504 26926 208532 38626
rect 208492 26920 208544 26926
rect 208492 26862 208544 26868
rect 208400 8968 208452 8974
rect 208400 8910 208452 8916
rect 208676 8968 208728 8974
rect 208676 8910 208728 8916
rect 207112 3596 207164 3602
rect 207112 3538 207164 3544
rect 207480 3596 207532 3602
rect 207480 3538 207532 3544
rect 206284 1148 206336 1154
rect 206284 1090 206336 1096
rect 206928 1148 206980 1154
rect 206928 1090 206980 1096
rect 206296 480 206324 1090
rect 207492 480 207520 3538
rect 208688 480 208716 8910
rect 209976 3534 210004 102054
rect 211068 15904 211120 15910
rect 211068 15846 211120 15852
rect 209964 3528 210016 3534
rect 209964 3470 210016 3476
rect 211080 3466 211108 15846
rect 211172 10334 211200 102054
rect 212092 96762 212120 102068
rect 212552 102054 212934 102082
rect 211436 96756 211488 96762
rect 211436 96698 211488 96704
rect 212080 96756 212132 96762
rect 212080 96698 212132 96704
rect 211448 80186 211476 96698
rect 211448 80158 211568 80186
rect 211540 80050 211568 80158
rect 211356 80022 211568 80050
rect 211356 53122 211384 80022
rect 211356 53094 211476 53122
rect 211448 41426 211476 53094
rect 211448 41398 211568 41426
rect 211540 38690 211568 41398
rect 211344 38684 211396 38690
rect 211344 38626 211396 38632
rect 211528 38684 211580 38690
rect 211528 38626 211580 38632
rect 211356 28286 211384 38626
rect 211344 28280 211396 28286
rect 211344 28222 211396 28228
rect 211160 10328 211212 10334
rect 211160 10270 211212 10276
rect 212264 10328 212316 10334
rect 212264 10270 212316 10276
rect 209872 3460 209924 3466
rect 209872 3402 209924 3408
rect 211068 3460 211120 3466
rect 211068 3402 211120 3408
rect 209884 480 209912 3402
rect 211068 3324 211120 3330
rect 211068 3266 211120 3272
rect 211080 480 211108 3266
rect 212276 480 212304 10270
rect 212552 3670 212580 102054
rect 213748 96665 213776 102068
rect 213932 102054 214682 102082
rect 215312 102054 215510 102082
rect 213090 96656 213146 96665
rect 213090 96591 213146 96600
rect 213734 96656 213790 96665
rect 213734 96591 213790 96600
rect 213104 82142 213132 96591
rect 212724 82136 212776 82142
rect 212724 82078 212776 82084
rect 213092 82136 213144 82142
rect 213092 82078 213144 82084
rect 212736 70514 212764 82078
rect 212724 70508 212776 70514
rect 212724 70450 212776 70456
rect 212724 67652 212776 67658
rect 212724 67594 212776 67600
rect 212736 66230 212764 67594
rect 212724 66224 212776 66230
rect 212724 66166 212776 66172
rect 212816 53848 212868 53854
rect 212816 53790 212868 53796
rect 212828 44130 212856 53790
rect 212816 44124 212868 44130
rect 212816 44066 212868 44072
rect 212816 28892 212868 28898
rect 212816 28834 212868 28840
rect 212828 26246 212856 28834
rect 212816 26240 212868 26246
rect 212816 26182 212868 26188
rect 212908 19304 212960 19310
rect 212908 19246 212960 19252
rect 212920 11762 212948 19246
rect 213932 17338 213960 102054
rect 214564 99408 214616 99414
rect 214564 99350 214616 99356
rect 214576 18698 214604 99350
rect 214564 18692 214616 18698
rect 214564 18634 214616 18640
rect 213920 17332 213972 17338
rect 213920 17274 213972 17280
rect 212908 11756 212960 11762
rect 212908 11698 212960 11704
rect 213460 9716 213512 9722
rect 213460 9658 213512 9664
rect 212540 3664 212592 3670
rect 212540 3606 212592 3612
rect 213472 480 213500 9658
rect 215312 3738 215340 102054
rect 216324 95266 216352 102068
rect 216692 102054 217166 102082
rect 215576 95260 215628 95266
rect 215576 95202 215628 95208
rect 216312 95260 216364 95266
rect 216312 95202 216364 95208
rect 215588 86986 215616 95202
rect 215496 86958 215616 86986
rect 215496 85542 215524 86958
rect 215484 85536 215536 85542
rect 215484 85478 215536 85484
rect 215392 75948 215444 75954
rect 215392 75890 215444 75896
rect 215404 62830 215432 75890
rect 215392 62824 215444 62830
rect 215392 62766 215444 62772
rect 215576 62824 215628 62830
rect 215576 62766 215628 62772
rect 215588 48346 215616 62766
rect 215484 48340 215536 48346
rect 215484 48282 215536 48288
rect 215576 48340 215628 48346
rect 215576 48282 215628 48288
rect 215496 41562 215524 48282
rect 215496 41534 215616 41562
rect 215588 41392 215616 41534
rect 215496 41364 215616 41392
rect 215496 13122 215524 41364
rect 216692 29646 216720 102054
rect 216680 29640 216732 29646
rect 216680 29582 216732 29588
rect 217968 18624 218020 18630
rect 217968 18566 218020 18572
rect 215484 13116 215536 13122
rect 215484 13058 215536 13064
rect 215852 11756 215904 11762
rect 215852 11698 215904 11704
rect 215300 3732 215352 3738
rect 215300 3674 215352 3680
rect 214656 3324 214708 3330
rect 214656 3266 214708 3272
rect 214668 480 214696 3266
rect 215864 480 215892 11698
rect 217980 3398 218008 18566
rect 218072 3806 218100 102068
rect 218900 96898 218928 102068
rect 219728 99414 219756 102068
rect 220280 102054 220662 102082
rect 220832 102054 221490 102082
rect 219716 99408 219768 99414
rect 219716 99350 219768 99356
rect 218336 96892 218388 96898
rect 218336 96834 218388 96840
rect 218888 96892 218940 96898
rect 218888 96834 218940 96840
rect 218348 87174 218376 96834
rect 220280 94466 220308 102054
rect 219636 94438 220308 94466
rect 218336 87168 218388 87174
rect 218336 87110 218388 87116
rect 218244 87032 218296 87038
rect 218244 86974 218296 86980
rect 218256 85542 218284 86974
rect 218244 85536 218296 85542
rect 218244 85478 218296 85484
rect 218152 75948 218204 75954
rect 218152 75890 218204 75896
rect 218164 62830 218192 75890
rect 218152 62824 218204 62830
rect 218152 62766 218204 62772
rect 218336 62824 218388 62830
rect 218336 62766 218388 62772
rect 218348 48346 218376 62766
rect 219636 60738 219664 94438
rect 219544 60710 219664 60738
rect 219544 60602 219572 60710
rect 219544 60574 219664 60602
rect 218244 48340 218296 48346
rect 218244 48282 218296 48288
rect 218336 48340 218388 48346
rect 218336 48282 218388 48288
rect 218256 14482 218284 48282
rect 219636 38826 219664 60574
rect 219624 38820 219676 38826
rect 219624 38762 219676 38768
rect 219624 38684 219676 38690
rect 219624 38626 219676 38632
rect 219636 31822 219664 38626
rect 219624 31816 219676 31822
rect 219624 31758 219676 31764
rect 219716 31680 219768 31686
rect 219716 31622 219768 31628
rect 219728 22114 219756 31622
rect 219544 22086 219756 22114
rect 218244 14476 218296 14482
rect 218244 14418 218296 14424
rect 219348 13116 219400 13122
rect 219348 13058 219400 13064
rect 218060 3800 218112 3806
rect 218060 3742 218112 3748
rect 218152 3732 218204 3738
rect 218152 3674 218204 3680
rect 217048 3392 217100 3398
rect 217048 3334 217100 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 217060 480 217088 3334
rect 218164 480 218192 3674
rect 219360 480 219388 13058
rect 219544 3942 219572 22086
rect 220544 9716 220596 9722
rect 220544 9658 220596 9664
rect 219532 3936 219584 3942
rect 219532 3878 219584 3884
rect 220556 480 220584 9658
rect 220832 6254 220860 102054
rect 222200 94580 222252 94586
rect 222200 94522 222252 94528
rect 220820 6248 220872 6254
rect 220820 6190 220872 6196
rect 222212 3874 222240 94522
rect 222304 19990 222332 102068
rect 222856 102054 223146 102082
rect 222856 94586 222884 102054
rect 224052 100026 224080 102068
rect 224236 102054 224894 102082
rect 225340 102054 225722 102082
rect 226352 102054 226642 102082
rect 226996 102054 227470 102082
rect 227732 102054 228298 102082
rect 224040 100020 224092 100026
rect 224040 99962 224092 99968
rect 222844 94580 222896 94586
rect 222844 94522 222896 94528
rect 224236 89842 224264 102054
rect 224144 89814 224264 89842
rect 224144 78606 224172 89814
rect 225340 87038 225368 102054
rect 224868 87032 224920 87038
rect 224868 86974 224920 86980
rect 225328 87032 225380 87038
rect 225328 86974 225380 86980
rect 224880 85542 224908 86974
rect 224868 85536 224920 85542
rect 224868 85478 224920 85484
rect 223672 78600 223724 78606
rect 223672 78542 223724 78548
rect 224132 78600 224184 78606
rect 224132 78542 224184 78548
rect 223684 51202 223712 78542
rect 224960 75948 225012 75954
rect 224960 75890 225012 75896
rect 224972 75834 225000 75890
rect 224880 75806 225000 75834
rect 224880 67538 224908 75806
rect 224880 67510 225092 67538
rect 225064 59906 225092 67510
rect 224868 59900 224920 59906
rect 224868 59842 224920 59848
rect 225052 59900 225104 59906
rect 225052 59842 225104 59848
rect 224880 52986 224908 59842
rect 224880 52958 225092 52986
rect 223672 51196 223724 51202
rect 223672 51138 223724 51144
rect 223672 51060 223724 51066
rect 223672 51002 223724 51008
rect 223684 38758 223712 51002
rect 225064 48278 225092 52958
rect 224960 48272 225012 48278
rect 224960 48214 225012 48220
rect 225052 48272 225104 48278
rect 225052 48214 225104 48220
rect 224972 46918 225000 48214
rect 224960 46912 225012 46918
rect 224960 46854 225012 46860
rect 223672 38752 223724 38758
rect 223672 38694 223724 38700
rect 223580 37324 223632 37330
rect 223580 37266 223632 37272
rect 224960 37324 225012 37330
rect 224960 37266 225012 37272
rect 223592 22778 223620 37266
rect 224972 31822 225000 37266
rect 224960 31816 225012 31822
rect 224960 31758 225012 31764
rect 224960 31680 225012 31686
rect 224960 31622 225012 31628
rect 224972 28966 225000 31622
rect 224960 28960 225012 28966
rect 224960 28902 225012 28908
rect 223580 22772 223632 22778
rect 223580 22714 223632 22720
rect 222292 19984 222344 19990
rect 222292 19926 222344 19932
rect 224960 19440 225012 19446
rect 224960 19382 225012 19388
rect 224972 19310 225000 19382
rect 224960 19304 225012 19310
rect 224960 19246 225012 19252
rect 225052 9716 225104 9722
rect 225052 9658 225104 9664
rect 222936 6180 222988 6186
rect 222936 6122 222988 6128
rect 222200 3868 222252 3874
rect 222200 3810 222252 3816
rect 221740 3664 221792 3670
rect 221740 3606 221792 3612
rect 221752 480 221780 3606
rect 222948 480 222976 6122
rect 225064 4078 225092 9658
rect 226352 4894 226380 102054
rect 226996 87009 227024 102054
rect 226522 87000 226578 87009
rect 226522 86935 226578 86944
rect 226982 87000 227038 87009
rect 226982 86935 227038 86944
rect 226536 85542 226564 86935
rect 226524 85536 226576 85542
rect 226524 85478 226576 85484
rect 226616 75948 226668 75954
rect 226616 75890 226668 75896
rect 226628 67726 226656 75890
rect 226616 67720 226668 67726
rect 226616 67662 226668 67668
rect 226524 67584 226576 67590
rect 226524 67526 226576 67532
rect 226536 63986 226564 67526
rect 226524 63980 226576 63986
rect 226524 63922 226576 63928
rect 226616 48340 226668 48346
rect 226616 48282 226668 48288
rect 226628 38622 226656 48282
rect 226616 38616 226668 38622
rect 226616 38558 226668 38564
rect 226616 29028 226668 29034
rect 226616 28970 226668 28976
rect 226628 24138 226656 28970
rect 226616 24132 226668 24138
rect 226616 24074 226668 24080
rect 226340 4888 226392 4894
rect 226340 4830 226392 4836
rect 226524 4820 226576 4826
rect 226524 4762 226576 4768
rect 225052 4072 225104 4078
rect 225052 4014 225104 4020
rect 225328 3936 225380 3942
rect 225328 3878 225380 3884
rect 224132 3392 224184 3398
rect 224132 3334 224184 3340
rect 224144 480 224172 3334
rect 225340 480 225368 3878
rect 226536 480 226564 4762
rect 227732 4010 227760 102054
rect 229006 75848 229062 75857
rect 229006 75783 229062 75792
rect 229020 66337 229048 75783
rect 229006 66328 229062 66337
rect 229006 66263 229062 66272
rect 229112 7614 229140 102068
rect 229664 102054 230046 102082
rect 230492 102054 230874 102082
rect 229664 85610 229692 102054
rect 229284 85604 229336 85610
rect 229284 85546 229336 85552
rect 229652 85604 229704 85610
rect 229652 85546 229704 85552
rect 229296 75857 229324 85546
rect 229282 75848 229338 75857
rect 229282 75783 229338 75792
rect 229282 66328 229338 66337
rect 229282 66263 229338 66272
rect 229296 66230 229324 66263
rect 229284 66224 229336 66230
rect 229284 66166 229336 66172
rect 229376 48340 229428 48346
rect 229376 48282 229428 48288
rect 229388 38622 229416 48282
rect 229376 38616 229428 38622
rect 229376 38558 229428 38564
rect 229376 29028 229428 29034
rect 229376 28970 229428 28976
rect 229388 22234 229416 28970
rect 229376 22228 229428 22234
rect 229376 22170 229428 22176
rect 229100 7608 229152 7614
rect 229100 7550 229152 7556
rect 230112 7608 230164 7614
rect 230112 7550 230164 7556
rect 227812 4072 227864 4078
rect 227812 4014 227864 4020
rect 227720 4004 227772 4010
rect 227720 3946 227772 3952
rect 227824 2122 227852 4014
rect 228916 3868 228968 3874
rect 228916 3810 228968 3816
rect 227732 2094 227852 2122
rect 227732 480 227760 2094
rect 228928 480 228956 3810
rect 230124 480 230152 7550
rect 230492 3602 230520 102054
rect 231688 95266 231716 102068
rect 231872 102054 232622 102082
rect 230848 95260 230900 95266
rect 230848 95202 230900 95208
rect 231676 95260 231728 95266
rect 231676 95202 231728 95208
rect 230860 87038 230888 95202
rect 230848 87032 230900 87038
rect 230848 86974 230900 86980
rect 230848 85604 230900 85610
rect 230848 85546 230900 85552
rect 230860 76702 230888 85546
rect 230848 76696 230900 76702
rect 230848 76638 230900 76644
rect 230848 76560 230900 76566
rect 230848 76502 230900 76508
rect 230860 67697 230888 76502
rect 230662 67688 230718 67697
rect 230662 67623 230718 67632
rect 230846 67688 230902 67697
rect 230846 67623 230902 67632
rect 230676 66230 230704 67623
rect 230664 66224 230716 66230
rect 230664 66166 230716 66172
rect 230756 66224 230808 66230
rect 230756 66166 230808 66172
rect 230768 53122 230796 66166
rect 230768 53094 230888 53122
rect 230860 38690 230888 53094
rect 230756 38684 230808 38690
rect 230756 38626 230808 38632
rect 230848 38684 230900 38690
rect 230848 38626 230900 38632
rect 230768 22166 230796 38626
rect 230756 22160 230808 22166
rect 230756 22102 230808 22108
rect 230664 19372 230716 19378
rect 230664 19314 230716 19320
rect 230676 12458 230704 19314
rect 231872 15910 231900 102054
rect 233332 94580 233384 94586
rect 233332 94522 233384 94528
rect 231860 15904 231912 15910
rect 231860 15846 231912 15852
rect 230676 12430 230796 12458
rect 230768 8974 230796 12430
rect 233344 10334 233372 94522
rect 233332 10328 233384 10334
rect 233332 10270 233384 10276
rect 230756 8968 230808 8974
rect 230756 8910 230808 8916
rect 231308 4004 231360 4010
rect 231308 3946 231360 3952
rect 230480 3596 230532 3602
rect 230480 3538 230532 3544
rect 231320 480 231348 3946
rect 232504 3596 232556 3602
rect 232504 3538 232556 3544
rect 232516 480 232544 3538
rect 233436 3466 233464 102068
rect 233896 102054 234278 102082
rect 234632 102054 235106 102082
rect 236026 102054 236224 102082
rect 233896 94586 233924 102054
rect 233884 94580 233936 94586
rect 233884 94522 233936 94528
rect 234632 17270 234660 102054
rect 236092 94580 236144 94586
rect 236092 94522 236144 94528
rect 234620 17264 234672 17270
rect 234620 17206 234672 17212
rect 236104 11762 236132 94522
rect 236092 11756 236144 11762
rect 236092 11698 236144 11704
rect 233700 10328 233752 10334
rect 233700 10270 233752 10276
rect 233424 3460 233476 3466
rect 233424 3402 233476 3408
rect 233712 480 233740 10270
rect 236000 4140 236052 4146
rect 236000 4082 236052 4088
rect 234804 3460 234856 3466
rect 234804 3402 234856 3408
rect 234816 480 234844 3402
rect 236012 480 236040 4082
rect 236196 3534 236224 102054
rect 236472 102054 236854 102082
rect 237484 102054 237682 102082
rect 238128 102054 238510 102082
rect 238772 102054 239430 102082
rect 236472 94586 236500 102054
rect 236460 94580 236512 94586
rect 236460 94522 236512 94528
rect 237380 94580 237432 94586
rect 237380 94522 237432 94528
rect 237196 8968 237248 8974
rect 237196 8910 237248 8916
rect 236184 3528 236236 3534
rect 236184 3470 236236 3476
rect 237208 480 237236 8910
rect 237392 3738 237420 94522
rect 237484 18630 237512 102054
rect 238128 94586 238156 102054
rect 238116 94580 238168 94586
rect 238116 94522 238168 94528
rect 237472 18624 237524 18630
rect 237472 18566 237524 18572
rect 238772 13122 238800 102054
rect 239404 99408 239456 99414
rect 239404 99350 239456 99356
rect 238760 13116 238812 13122
rect 238760 13058 238812 13064
rect 239416 6186 239444 99350
rect 240140 94580 240192 94586
rect 240140 94522 240192 94528
rect 239404 6180 239456 6186
rect 239404 6122 239456 6128
rect 237380 3732 237432 3738
rect 237380 3674 237432 3680
rect 239588 3732 239640 3738
rect 239588 3674 239640 3680
rect 238392 3528 238444 3534
rect 238392 3470 238444 3476
rect 238404 480 238432 3470
rect 239600 480 239628 3674
rect 240152 3670 240180 94522
rect 240244 14482 240272 102068
rect 240704 102054 241086 102082
rect 240704 94586 240732 102054
rect 241992 99414 242020 102068
rect 242452 102054 242834 102082
rect 241980 99408 242032 99414
rect 241980 99350 242032 99356
rect 240692 94580 240744 94586
rect 240692 94522 240744 94528
rect 242452 94466 242480 102054
rect 241808 94438 242480 94466
rect 241808 84250 241836 94438
rect 243004 89842 243032 102190
rect 244384 102054 244490 102082
rect 245120 102054 245410 102082
rect 245672 102054 246238 102082
rect 244280 92404 244332 92410
rect 244280 92346 244332 92352
rect 242912 89814 243032 89842
rect 241612 84244 241664 84250
rect 241612 84186 241664 84192
rect 241796 84244 241848 84250
rect 241796 84186 241848 84192
rect 241624 80050 241652 84186
rect 241624 80022 241744 80050
rect 241716 70394 241744 80022
rect 241716 70366 241836 70394
rect 241808 48346 241836 70366
rect 241704 48340 241756 48346
rect 241704 48282 241756 48288
rect 241796 48340 241848 48346
rect 241796 48282 241848 48288
rect 241716 41426 241744 48282
rect 241716 41398 241836 41426
rect 241808 31770 241836 41398
rect 241624 31742 241836 31770
rect 241624 31634 241652 31742
rect 241624 31606 241744 31634
rect 240232 14476 240284 14482
rect 240232 14418 240284 14424
rect 241716 12458 241744 31606
rect 241624 12430 241744 12458
rect 240784 6180 240836 6186
rect 240784 6122 240836 6128
rect 240140 3664 240192 3670
rect 240140 3606 240192 3612
rect 240796 480 240824 6122
rect 241624 3398 241652 12430
rect 242912 3942 242940 89814
rect 244292 4078 244320 92346
rect 244384 4826 244412 102054
rect 245120 92410 245148 102054
rect 245108 92404 245160 92410
rect 245108 92346 245160 92352
rect 244372 4820 244424 4826
rect 244372 4762 244424 4768
rect 244464 4820 244516 4826
rect 244464 4762 244516 4768
rect 244280 4072 244332 4078
rect 244280 4014 244332 4020
rect 242900 3936 242952 3942
rect 242900 3878 242952 3884
rect 243176 3936 243228 3942
rect 243176 3878 243228 3884
rect 241980 3800 242032 3806
rect 241980 3742 242032 3748
rect 241612 3392 241664 3398
rect 241612 3334 241664 3340
rect 241992 480 242020 3742
rect 243188 480 243216 3878
rect 244476 2394 244504 4762
rect 245672 3874 245700 102054
rect 247052 94738 247080 102068
rect 247696 102054 247986 102082
rect 248432 102054 248814 102082
rect 247052 94710 247172 94738
rect 247040 94580 247092 94586
rect 247040 94522 247092 94528
rect 247052 4010 247080 94522
rect 247144 7614 247172 94710
rect 247696 94586 247724 102054
rect 247684 94580 247736 94586
rect 247684 94522 247736 94528
rect 247132 7608 247184 7614
rect 247132 7550 247184 7556
rect 247040 4004 247092 4010
rect 247040 3946 247092 3952
rect 247960 4004 248012 4010
rect 247960 3946 248012 3952
rect 245660 3868 245712 3874
rect 245660 3810 245712 3816
rect 246764 3868 246816 3874
rect 246764 3810 246816 3816
rect 245568 3664 245620 3670
rect 245568 3606 245620 3612
rect 244384 2366 244504 2394
rect 244384 480 244412 2366
rect 245580 480 245608 3606
rect 246776 480 246804 3810
rect 247972 480 248000 3946
rect 248432 3602 248460 102054
rect 248984 87038 249012 102190
rect 249812 102054 250470 102082
rect 251192 102054 251390 102082
rect 248880 87032 248932 87038
rect 248880 86974 248932 86980
rect 248972 87032 249024 87038
rect 248972 86974 249024 86980
rect 248892 80170 248920 86974
rect 248880 80164 248932 80170
rect 248880 80106 248932 80112
rect 248604 77308 248656 77314
rect 248604 77250 248656 77256
rect 248616 70446 248644 77250
rect 248604 70440 248656 70446
rect 248604 70382 248656 70388
rect 248604 67652 248656 67658
rect 248604 67594 248656 67600
rect 248616 67538 248644 67594
rect 248616 67510 248736 67538
rect 248708 60790 248736 67510
rect 248696 60784 248748 60790
rect 248696 60726 248748 60732
rect 248696 60648 248748 60654
rect 248696 60590 248748 60596
rect 248708 48249 248736 60590
rect 248694 48240 248750 48249
rect 248694 48175 248750 48184
rect 248970 48240 249026 48249
rect 248970 48175 249026 48184
rect 248984 46918 249012 48175
rect 248972 46912 249024 46918
rect 248972 46854 249024 46860
rect 248972 37324 249024 37330
rect 248972 37266 249024 37272
rect 248984 29034 249012 37266
rect 248696 29028 248748 29034
rect 248696 28970 248748 28976
rect 248972 29028 249024 29034
rect 248972 28970 249024 28976
rect 248708 22114 248736 28970
rect 248616 22086 248736 22114
rect 248616 19310 248644 22086
rect 248604 19304 248656 19310
rect 248604 19246 248656 19252
rect 249156 4072 249208 4078
rect 249156 4014 249208 4020
rect 248420 3596 248472 3602
rect 248420 3538 248472 3544
rect 249168 480 249196 4014
rect 249812 3466 249840 102054
rect 251192 4146 251220 102054
rect 251560 93838 251588 102190
rect 252572 102054 253046 102082
rect 251548 93832 251600 93838
rect 251548 93774 251600 93780
rect 251456 84244 251508 84250
rect 251456 84186 251508 84192
rect 251468 72434 251496 84186
rect 251376 72406 251496 72434
rect 251376 67590 251404 72406
rect 252468 71596 252520 71602
rect 252468 71538 252520 71544
rect 251364 67584 251416 67590
rect 251364 67526 251416 67532
rect 251456 67516 251508 67522
rect 251456 67458 251508 67464
rect 251468 22114 251496 67458
rect 252480 58002 252508 71538
rect 252468 57996 252520 58002
rect 252468 57938 252520 57944
rect 252572 48414 252600 102054
rect 253216 89842 253244 102190
rect 253032 89814 253244 89842
rect 254044 102054 254794 102082
rect 255332 102054 255622 102082
rect 253032 89706 253060 89814
rect 252756 89678 253060 89706
rect 252756 86970 252784 89678
rect 252744 86964 252796 86970
rect 252744 86906 252796 86912
rect 252652 77308 252704 77314
rect 252652 77250 252704 77256
rect 252664 71602 252692 77250
rect 252652 71596 252704 71602
rect 252652 71538 252704 71544
rect 254044 62778 254072 102054
rect 254044 62750 254164 62778
rect 252652 57996 252704 58002
rect 252652 57938 252704 57944
rect 252664 48482 252692 57938
rect 252652 48476 252704 48482
rect 252652 48418 252704 48424
rect 252560 48408 252612 48414
rect 252560 48350 252612 48356
rect 252560 48204 252612 48210
rect 252560 48146 252612 48152
rect 252468 46980 252520 46986
rect 252468 46922 252520 46928
rect 252480 38690 252508 46922
rect 252468 38684 252520 38690
rect 252468 38626 252520 38632
rect 251376 22086 251496 22114
rect 251376 12510 251404 22086
rect 251364 12504 251416 12510
rect 251364 12446 251416 12452
rect 251272 12436 251324 12442
rect 251272 12378 251324 12384
rect 251284 8974 251312 12378
rect 251272 8968 251324 8974
rect 251272 8910 251324 8916
rect 251180 4140 251232 4146
rect 251180 4082 251232 4088
rect 251456 3596 251508 3602
rect 251456 3538 251508 3544
rect 249800 3460 249852 3466
rect 249800 3402 249852 3408
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 250364 480 250392 3334
rect 251468 480 251496 3538
rect 252572 3534 252600 48146
rect 252652 38684 252704 38690
rect 252652 38626 252704 38632
rect 252664 3738 252692 38626
rect 254136 22302 254164 62750
rect 254124 22296 254176 22302
rect 254124 22238 254176 22244
rect 254124 22160 254176 22166
rect 254124 22102 254176 22108
rect 254136 12050 254164 22102
rect 254136 12022 254256 12050
rect 254228 11778 254256 12022
rect 254136 11750 254256 11778
rect 254136 6186 254164 11750
rect 254124 6180 254176 6186
rect 254124 6122 254176 6128
rect 252744 4140 252796 4146
rect 252744 4082 252796 4088
rect 252652 3732 252704 3738
rect 252652 3674 252704 3680
rect 252560 3528 252612 3534
rect 252560 3470 252612 3476
rect 252756 2122 252784 4082
rect 255332 3806 255360 102054
rect 256436 95266 256464 102068
rect 256712 102054 257370 102082
rect 258092 102054 258198 102082
rect 255872 95260 255924 95266
rect 255872 95202 255924 95208
rect 256424 95260 256476 95266
rect 256424 95202 256476 95208
rect 255884 87145 255912 95202
rect 255870 87136 255926 87145
rect 255870 87071 255926 87080
rect 255410 87000 255466 87009
rect 255410 86935 255466 86944
rect 255424 67810 255452 86935
rect 255424 67782 255544 67810
rect 255516 67658 255544 67782
rect 255412 67652 255464 67658
rect 255412 67594 255464 67600
rect 255504 67652 255556 67658
rect 255504 67594 255556 67600
rect 255424 27606 255452 67594
rect 255412 27600 255464 27606
rect 255412 27542 255464 27548
rect 255412 18012 255464 18018
rect 255412 17954 255464 17960
rect 255424 3942 255452 17954
rect 256712 4826 256740 102054
rect 256700 4820 256752 4826
rect 256700 4762 256752 4768
rect 255412 3936 255464 3942
rect 255412 3878 255464 3884
rect 255320 3800 255372 3806
rect 255320 3742 255372 3748
rect 256240 3800 256292 3806
rect 256240 3742 256292 3748
rect 253848 3528 253900 3534
rect 253848 3470 253900 3476
rect 252664 2094 252784 2122
rect 252664 480 252692 2094
rect 253860 480 253888 3470
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 255056 480 255084 3402
rect 256252 480 256280 3742
rect 257436 3732 257488 3738
rect 257436 3674 257488 3680
rect 257448 480 257476 3674
rect 258092 3670 258120 102054
rect 259012 95266 259040 102068
rect 259564 102054 259854 102082
rect 260392 102054 260774 102082
rect 261220 102054 261602 102082
rect 262324 102054 262430 102082
rect 262968 102054 263350 102082
rect 263612 102054 264178 102082
rect 258356 95260 258408 95266
rect 258356 95202 258408 95208
rect 259000 95260 259052 95266
rect 259000 95202 259052 95208
rect 258368 93838 258396 95202
rect 258356 93832 258408 93838
rect 258356 93774 258408 93780
rect 259460 91316 259512 91322
rect 259460 91258 259512 91264
rect 258264 84244 258316 84250
rect 258264 84186 258316 84192
rect 258276 77382 258304 84186
rect 258264 77376 258316 77382
rect 258264 77318 258316 77324
rect 258264 77240 258316 77246
rect 258264 77182 258316 77188
rect 258276 66298 258304 77182
rect 258172 66292 258224 66298
rect 258172 66234 258224 66240
rect 258264 66292 258316 66298
rect 258264 66234 258316 66240
rect 258184 56506 258212 66234
rect 258172 56500 258224 56506
rect 258172 56442 258224 56448
rect 258172 46980 258224 46986
rect 258172 46922 258224 46928
rect 258184 38622 258212 46922
rect 258172 38616 258224 38622
rect 258172 38558 258224 38564
rect 258264 38616 258316 38622
rect 258264 38558 258316 38564
rect 258276 12458 258304 38558
rect 258276 12430 258396 12458
rect 258368 3874 258396 12430
rect 259472 4078 259500 91258
rect 259460 4072 259512 4078
rect 259460 4014 259512 4020
rect 259564 4010 259592 102054
rect 260392 91322 260420 102054
rect 260380 91316 260432 91322
rect 260380 91258 260432 91264
rect 261220 77353 261248 102054
rect 262220 92404 262272 92410
rect 262220 92346 262272 92352
rect 261206 77344 261262 77353
rect 261206 77279 261262 77288
rect 260838 77208 260894 77217
rect 260838 77143 260894 77152
rect 260852 57934 260880 77143
rect 260840 57928 260892 57934
rect 260840 57870 260892 57876
rect 260840 48340 260892 48346
rect 260840 48282 260892 48288
rect 260852 48210 260880 48282
rect 260840 48204 260892 48210
rect 260840 48146 260892 48152
rect 260840 38752 260892 38758
rect 260840 38694 260892 38700
rect 260852 19310 260880 38694
rect 260840 19304 260892 19310
rect 260840 19246 260892 19252
rect 261024 9716 261076 9722
rect 261024 9658 261076 9664
rect 259552 4004 259604 4010
rect 259552 3946 259604 3952
rect 259828 3936 259880 3942
rect 259828 3878 259880 3884
rect 258356 3868 258408 3874
rect 258356 3810 258408 3816
rect 258080 3664 258132 3670
rect 258080 3606 258132 3612
rect 258632 3324 258684 3330
rect 258632 3266 258684 3272
rect 258644 480 258672 3266
rect 259840 480 259868 3878
rect 261036 3398 261064 9658
rect 262232 4146 262260 92346
rect 262220 4140 262272 4146
rect 262220 4082 262272 4088
rect 262220 3868 262272 3874
rect 262220 3810 262272 3816
rect 261024 3392 261076 3398
rect 261024 3334 261076 3340
rect 261024 3052 261076 3058
rect 261024 2994 261076 3000
rect 261036 480 261064 2994
rect 262232 480 262260 3810
rect 262324 3602 262352 102054
rect 262968 92410 262996 102054
rect 262956 92404 263008 92410
rect 262956 92346 263008 92352
rect 262312 3596 262364 3602
rect 262312 3538 262364 3544
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 263428 480 263456 3538
rect 263612 3534 263640 102054
rect 264992 94738 265020 102068
rect 265544 102054 265834 102082
rect 266372 102054 266754 102082
rect 267016 102054 267582 102082
rect 267752 102054 268410 102082
rect 269132 102054 269238 102082
rect 269776 102054 270158 102082
rect 270604 102054 270986 102082
rect 271432 102054 271814 102082
rect 272260 102054 272734 102082
rect 273364 102054 273562 102082
rect 274008 102054 274390 102082
rect 274652 102054 275218 102082
rect 264992 94710 265112 94738
rect 264980 94580 265032 94586
rect 264980 94522 265032 94528
rect 264992 3806 265020 94522
rect 264980 3800 265032 3806
rect 264980 3742 265032 3748
rect 264612 3596 264664 3602
rect 264612 3538 264664 3544
rect 263600 3528 263652 3534
rect 263600 3470 263652 3476
rect 264624 480 264652 3538
rect 265084 3466 265112 94710
rect 265544 94586 265572 102054
rect 265532 94580 265584 94586
rect 265532 94522 265584 94528
rect 266372 3738 266400 102054
rect 267016 89842 267044 102054
rect 266832 89814 267044 89842
rect 266832 80016 266860 89814
rect 266648 79988 266860 80016
rect 266648 60858 266676 79988
rect 266636 60852 266688 60858
rect 266636 60794 266688 60800
rect 266544 60784 266596 60790
rect 266544 60726 266596 60732
rect 266556 57934 266584 60726
rect 266544 57928 266596 57934
rect 266544 57870 266596 57876
rect 266452 48340 266504 48346
rect 266452 48282 266504 48288
rect 266464 38690 266492 48282
rect 266452 38684 266504 38690
rect 266452 38626 266504 38632
rect 266544 38684 266596 38690
rect 266544 38626 266596 38632
rect 266556 22114 266584 38626
rect 266464 22086 266584 22114
rect 266464 21978 266492 22086
rect 266464 21950 266584 21978
rect 266360 3732 266412 3738
rect 266360 3674 266412 3680
rect 265072 3460 265124 3466
rect 265072 3402 265124 3408
rect 266556 3330 266584 21950
rect 267752 3942 267780 102054
rect 267740 3936 267792 3942
rect 267740 3878 267792 3884
rect 268108 3664 268160 3670
rect 268108 3606 268160 3612
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 266544 3324 266596 3330
rect 266544 3266 266596 3272
rect 265808 3188 265860 3194
rect 265808 3130 265860 3136
rect 265820 480 265848 3130
rect 267016 480 267044 3402
rect 268120 480 268148 3606
rect 269132 3058 269160 102054
rect 269776 89842 269804 102054
rect 270500 91588 270552 91594
rect 270500 91530 270552 91536
rect 269592 89814 269804 89842
rect 269592 80016 269620 89814
rect 269408 79988 269620 80016
rect 269408 60874 269436 79988
rect 269316 60846 269436 60874
rect 269316 60738 269344 60846
rect 269224 60710 269344 60738
rect 269224 60602 269252 60710
rect 269224 60574 269344 60602
rect 269316 41426 269344 60574
rect 269224 41398 269344 41426
rect 269224 41290 269252 41398
rect 269224 41262 269344 41290
rect 269316 22114 269344 41262
rect 269224 22086 269344 22114
rect 269224 21978 269252 22086
rect 269224 21950 269344 21978
rect 269316 3874 269344 21950
rect 269304 3868 269356 3874
rect 269304 3810 269356 3816
rect 269304 3732 269356 3738
rect 269304 3674 269356 3680
rect 269120 3052 269172 3058
rect 269120 2994 269172 3000
rect 269316 480 269344 3674
rect 270512 3602 270540 91530
rect 270500 3596 270552 3602
rect 270500 3538 270552 3544
rect 270604 3534 270632 102054
rect 271432 91594 271460 102054
rect 271420 91588 271472 91594
rect 271420 91530 271472 91536
rect 272260 89842 272288 102054
rect 273260 92404 273312 92410
rect 273260 92346 273312 92352
rect 272168 89814 272288 89842
rect 272168 80238 272196 89814
rect 272156 80232 272208 80238
rect 272156 80174 272208 80180
rect 272064 77308 272116 77314
rect 272064 77250 272116 77256
rect 272076 58002 272104 77250
rect 271972 57996 272024 58002
rect 271972 57938 272024 57944
rect 272064 57996 272116 58002
rect 272064 57938 272116 57944
rect 271984 57882 272012 57938
rect 271984 57854 272104 57882
rect 272076 48346 272104 57854
rect 271972 48340 272024 48346
rect 271972 48282 272024 48288
rect 272064 48340 272116 48346
rect 272064 48282 272116 48288
rect 271984 43518 272012 48282
rect 271972 43512 272024 43518
rect 271972 43454 272024 43460
rect 272248 43512 272300 43518
rect 272248 43454 272300 43460
rect 272260 38729 272288 43454
rect 272062 38720 272118 38729
rect 271984 38678 272062 38706
rect 271984 38622 272012 38678
rect 272062 38655 272118 38664
rect 272246 38720 272302 38729
rect 272246 38655 272302 38664
rect 271788 38616 271840 38622
rect 271788 38558 271840 38564
rect 271972 38616 272024 38622
rect 271972 38558 272024 38564
rect 271800 29073 271828 38558
rect 271786 29064 271842 29073
rect 271786 28999 271842 29008
rect 271970 29064 272026 29073
rect 271970 28999 272026 29008
rect 271984 28966 272012 28999
rect 271972 28960 272024 28966
rect 271972 28902 272024 28908
rect 271972 19372 272024 19378
rect 271972 19314 272024 19320
rect 271984 9654 272012 19314
rect 271972 9648 272024 9654
rect 271972 9590 272024 9596
rect 271696 4140 271748 4146
rect 271696 4082 271748 4088
rect 270592 3528 270644 3534
rect 270592 3470 270644 3476
rect 270500 3392 270552 3398
rect 270500 3334 270552 3340
rect 270512 480 270540 3334
rect 271708 480 271736 4082
rect 273272 3670 273300 92346
rect 273260 3664 273312 3670
rect 273260 3606 273312 3612
rect 272892 3528 272944 3534
rect 272892 3470 272944 3476
rect 272904 480 272932 3470
rect 273364 3466 273392 102054
rect 274008 92410 274036 102054
rect 273996 92404 274048 92410
rect 273996 92346 274048 92352
rect 274652 3738 274680 102054
rect 276020 94580 276072 94586
rect 276020 94522 276072 94528
rect 276032 4146 276060 94522
rect 276020 4140 276072 4146
rect 276020 4082 276072 4088
rect 275284 4072 275336 4078
rect 275284 4014 275336 4020
rect 274640 3732 274692 3738
rect 274640 3674 274692 3680
rect 273352 3460 273404 3466
rect 273352 3402 273404 3408
rect 274088 3052 274140 3058
rect 274088 2994 274140 3000
rect 274100 480 274128 2994
rect 275296 480 275324 4014
rect 276124 3398 276152 102068
rect 276584 102054 276966 102082
rect 277412 102054 277794 102082
rect 276584 94586 276612 102054
rect 276572 94580 276624 94586
rect 276572 94522 276624 94528
rect 276480 3800 276532 3806
rect 276480 3742 276532 3748
rect 276112 3392 276164 3398
rect 276112 3334 276164 3340
rect 276492 480 276520 3742
rect 277412 3534 277440 102054
rect 277964 89842 277992 102190
rect 279160 102054 279542 102082
rect 280172 102054 280370 102082
rect 279160 89842 279188 102054
rect 277688 89814 277992 89842
rect 278976 89814 279188 89842
rect 277688 77314 277716 89814
rect 278976 77314 279004 89814
rect 277584 77308 277636 77314
rect 277584 77250 277636 77256
rect 277676 77308 277728 77314
rect 277676 77250 277728 77256
rect 278872 77308 278924 77314
rect 278872 77250 278924 77256
rect 278964 77308 279016 77314
rect 278964 77250 279016 77256
rect 277596 70446 277624 77250
rect 277584 70440 277636 70446
rect 277584 70382 277636 70388
rect 277492 70372 277544 70378
rect 277492 70314 277544 70320
rect 277504 60926 277532 70314
rect 277492 60920 277544 60926
rect 277492 60862 277544 60868
rect 277584 60716 277636 60722
rect 277584 60658 277636 60664
rect 277596 41426 277624 60658
rect 278884 41426 278912 77250
rect 277504 41398 277624 41426
rect 278792 41398 278912 41426
rect 277504 41290 277532 41398
rect 278792 41290 278820 41398
rect 277504 41262 277624 41290
rect 278792 41262 278912 41290
rect 277596 22114 277624 41262
rect 278884 22114 278912 41262
rect 277504 22086 277624 22114
rect 278792 22086 278912 22114
rect 277504 21978 277532 22086
rect 278792 21978 278820 22086
rect 277504 21950 277624 21978
rect 278792 21950 278912 21978
rect 277400 3528 277452 3534
rect 277400 3470 277452 3476
rect 277596 3058 277624 21950
rect 278884 4162 278912 21950
rect 277676 4140 277728 4146
rect 277676 4082 277728 4088
rect 278700 4134 278912 4162
rect 277584 3052 277636 3058
rect 277584 2994 277636 3000
rect 277688 480 277716 4082
rect 278700 4078 278728 4134
rect 278688 4072 278740 4078
rect 278688 4014 278740 4020
rect 278872 4072 278924 4078
rect 278872 4014 278924 4020
rect 278884 480 278912 4014
rect 280172 3806 280200 102054
rect 280540 89842 280568 102190
rect 280448 89814 280568 89842
rect 281552 102054 282118 102082
rect 280448 67658 280476 89814
rect 280344 67652 280396 67658
rect 280344 67594 280396 67600
rect 280436 67652 280488 67658
rect 280436 67594 280488 67600
rect 280356 41426 280384 67594
rect 280264 41398 280384 41426
rect 280264 41290 280292 41398
rect 280264 41262 280384 41290
rect 280356 22114 280384 41262
rect 280264 22086 280384 22114
rect 280264 21978 280292 22086
rect 280264 21950 280384 21978
rect 280356 4146 280384 21950
rect 280344 4140 280396 4146
rect 280344 4082 280396 4088
rect 281552 4078 281580 102054
rect 281540 4072 281592 4078
rect 281540 4014 281592 4020
rect 282460 4072 282512 4078
rect 282460 4014 282512 4020
rect 280160 3800 280212 3806
rect 280160 3742 280212 3748
rect 280068 3460 280120 3466
rect 280068 3402 280120 3408
rect 280080 480 280108 3402
rect 281264 3052 281316 3058
rect 281264 2994 281316 3000
rect 281276 480 281304 2994
rect 282472 480 282500 4014
rect 282932 3466 282960 102068
rect 283392 102054 283774 102082
rect 284312 102054 284602 102082
rect 283392 89842 283420 102054
rect 283208 89814 283420 89842
rect 283208 70258 283236 89814
rect 283116 70230 283236 70258
rect 283116 67590 283144 70230
rect 283104 67584 283156 67590
rect 283104 67526 283156 67532
rect 283104 57996 283156 58002
rect 283104 57938 283156 57944
rect 283116 41426 283144 57938
rect 283024 41398 283144 41426
rect 283024 41290 283052 41398
rect 283024 41262 283144 41290
rect 283116 22114 283144 41262
rect 283024 22086 283144 22114
rect 283024 21978 283052 22086
rect 283024 21950 283144 21978
rect 282920 3460 282972 3466
rect 282920 3402 282972 3408
rect 283116 3058 283144 21950
rect 283656 9648 283708 9654
rect 283656 9590 283708 9596
rect 283104 3052 283156 3058
rect 283104 2994 283156 3000
rect 283668 480 283696 9590
rect 284312 4078 284340 102054
rect 284772 85610 284800 102190
rect 285692 102054 286350 102082
rect 287072 102054 287178 102082
rect 287808 102054 288098 102082
rect 288452 102054 288926 102082
rect 284576 85604 284628 85610
rect 284576 85546 284628 85552
rect 284760 85604 284812 85610
rect 284760 85546 284812 85552
rect 284588 77382 284616 85546
rect 284576 77376 284628 77382
rect 284576 77318 284628 77324
rect 284392 77240 284444 77246
rect 284392 77182 284444 77188
rect 284404 67658 284432 77182
rect 284392 67652 284444 67658
rect 284392 67594 284444 67600
rect 284484 67652 284536 67658
rect 284484 67594 284536 67600
rect 284496 41426 284524 67594
rect 284496 41398 284616 41426
rect 284588 38706 284616 41398
rect 284496 38678 284616 38706
rect 284496 38622 284524 38678
rect 284484 38616 284536 38622
rect 284484 38558 284536 38564
rect 284484 29096 284536 29102
rect 284484 29038 284536 29044
rect 284496 28966 284524 29038
rect 284484 28960 284536 28966
rect 284484 28902 284536 28908
rect 284484 19372 284536 19378
rect 284484 19314 284536 19320
rect 284496 9654 284524 19314
rect 284484 9648 284536 9654
rect 284484 9590 284536 9596
rect 285692 4146 285720 102054
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 285680 4140 285732 4146
rect 285680 4082 285732 4088
rect 284300 4072 284352 4078
rect 284300 4014 284352 4020
rect 284772 480 284800 4082
rect 287072 3602 287100 102054
rect 287808 89842 287836 102054
rect 287440 89814 287836 89842
rect 287440 80238 287468 89814
rect 287428 80232 287480 80238
rect 287428 80174 287480 80180
rect 287336 77308 287388 77314
rect 287336 77250 287388 77256
rect 287348 66230 287376 77250
rect 287336 66224 287388 66230
rect 287336 66166 287388 66172
rect 287244 56636 287296 56642
rect 287244 56578 287296 56584
rect 287256 48278 287284 56578
rect 287244 48272 287296 48278
rect 287244 48214 287296 48220
rect 287244 39840 287296 39846
rect 287244 39782 287296 39788
rect 287256 28966 287284 39782
rect 287244 28960 287296 28966
rect 287244 28902 287296 28908
rect 287336 19372 287388 19378
rect 287336 19314 287388 19320
rect 285956 3596 286008 3602
rect 285956 3538 286008 3544
rect 287060 3596 287112 3602
rect 287060 3538 287112 3544
rect 285968 480 285996 3538
rect 287348 610 287376 19314
rect 288452 4060 288480 102054
rect 289096 89842 289124 102190
rect 290200 102054 290582 102082
rect 291304 102054 291502 102082
rect 292330 102054 292528 102082
rect 290200 89842 290228 102054
rect 288636 89814 289124 89842
rect 290108 89814 290228 89842
rect 288636 80186 288664 89814
rect 290108 86970 290136 89814
rect 290096 86964 290148 86970
rect 290096 86906 290148 86912
rect 288544 80158 288664 80186
rect 288544 4146 288572 80158
rect 290004 77308 290056 77314
rect 290004 77250 290056 77256
rect 290016 60874 290044 77250
rect 289924 60846 290044 60874
rect 289924 60738 289952 60846
rect 289832 60710 289952 60738
rect 289832 60602 289860 60710
rect 289832 60574 289952 60602
rect 289924 41426 289952 60574
rect 289832 41398 289952 41426
rect 289832 41290 289860 41398
rect 289832 41262 289952 41290
rect 289924 22114 289952 41262
rect 289832 22086 289952 22114
rect 289832 21978 289860 22086
rect 289832 21950 289952 21978
rect 289924 4146 289952 21950
rect 291304 4146 291332 102054
rect 288532 4140 288584 4146
rect 288532 4082 288584 4088
rect 289544 4140 289596 4146
rect 289544 4082 289596 4088
rect 289912 4140 289964 4146
rect 289912 4082 289964 4088
rect 290740 4140 290792 4146
rect 290740 4082 290792 4088
rect 291292 4140 291344 4146
rect 291292 4082 291344 4088
rect 291936 4140 291988 4146
rect 291936 4082 291988 4088
rect 288360 4032 288480 4060
rect 287152 604 287204 610
rect 287152 546 287204 552
rect 287336 604 287388 610
rect 287336 546 287388 552
rect 287164 480 287192 546
rect 288360 480 288388 4032
rect 289556 480 289584 4082
rect 290752 480 290780 4082
rect 291948 480 291976 4082
rect 292500 3466 292528 102054
rect 293144 99414 293172 102068
rect 294064 99414 294092 102068
rect 294906 102054 295288 102082
rect 293132 99408 293184 99414
rect 293132 99350 293184 99356
rect 293868 99408 293920 99414
rect 293868 99350 293920 99356
rect 294052 99408 294104 99414
rect 294052 99350 294104 99356
rect 295156 99408 295208 99414
rect 295156 99350 295208 99356
rect 292488 3460 292540 3466
rect 292488 3402 292540 3408
rect 293132 3460 293184 3466
rect 293132 3402 293184 3408
rect 293144 480 293172 3402
rect 293880 3194 293908 99350
rect 295168 3482 295196 99350
rect 295260 4146 295288 102054
rect 295720 99414 295748 102068
rect 295708 99408 295760 99414
rect 295708 99350 295760 99356
rect 295248 4140 295300 4146
rect 295248 4082 295300 4088
rect 295168 3454 295564 3482
rect 293868 3188 293920 3194
rect 293868 3130 293920 3136
rect 294328 3188 294380 3194
rect 294328 3130 294380 3136
rect 294340 480 294368 3130
rect 295536 480 295564 3454
rect 296548 2922 296576 102068
rect 297482 102054 298048 102082
rect 296628 99408 296680 99414
rect 296628 99350 296680 99356
rect 296640 4078 296668 99350
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 296628 4072 296680 4078
rect 296628 4014 296680 4020
rect 296536 2916 296588 2922
rect 296536 2858 296588 2864
rect 296732 480 296760 4082
rect 297916 4072 297968 4078
rect 297916 4014 297968 4020
rect 297928 480 297956 4014
rect 298020 3126 298048 102054
rect 298296 99414 298324 102068
rect 299138 102054 299336 102082
rect 300058 102054 300808 102082
rect 298284 99408 298336 99414
rect 298284 99350 298336 99356
rect 299308 3398 299336 102054
rect 299388 99408 299440 99414
rect 299388 99350 299440 99356
rect 299296 3392 299348 3398
rect 299296 3334 299348 3340
rect 298008 3120 298060 3126
rect 298008 3062 298060 3068
rect 299400 3058 299428 99350
rect 300780 3534 300808 102054
rect 300872 99414 300900 102068
rect 301714 102054 302096 102082
rect 300860 99408 300912 99414
rect 300860 99350 300912 99356
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 302068 3330 302096 102054
rect 302528 100706 302556 102068
rect 302516 100700 302568 100706
rect 302516 100642 302568 100648
rect 302148 99408 302200 99414
rect 302148 99350 302200 99356
rect 302056 3324 302108 3330
rect 302056 3266 302108 3272
rect 302160 3194 302188 99350
rect 303448 3942 303476 102068
rect 304290 102054 304948 102082
rect 303528 100700 303580 100706
rect 303528 100642 303580 100648
rect 303540 4146 303568 100642
rect 303528 4140 303580 4146
rect 303528 4082 303580 4088
rect 304920 4010 304948 102054
rect 305104 100638 305132 102068
rect 305946 102054 306236 102082
rect 306866 102054 307616 102082
rect 305092 100632 305144 100638
rect 305092 100574 305144 100580
rect 304908 4004 304960 4010
rect 304908 3946 304960 3952
rect 303436 3936 303488 3942
rect 303436 3878 303488 3884
rect 306208 3534 306236 102054
rect 306288 100632 306340 100638
rect 306288 100574 306340 100580
rect 306300 4078 306328 100574
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 306288 4072 306340 4078
rect 306288 4014 306340 4020
rect 303804 3528 303856 3534
rect 303804 3470 303856 3476
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 302608 3392 302660 3398
rect 302608 3334 302660 3340
rect 302148 3188 302200 3194
rect 302148 3130 302200 3136
rect 300308 3120 300360 3126
rect 300308 3062 300360 3068
rect 299388 3052 299440 3058
rect 299388 2994 299440 3000
rect 299112 2916 299164 2922
rect 299112 2858 299164 2864
rect 299124 480 299152 2858
rect 300320 480 300348 3062
rect 301412 3052 301464 3058
rect 301412 2994 301464 3000
rect 301424 480 301452 2994
rect 302620 480 302648 3334
rect 303816 480 303844 3470
rect 306196 3324 306248 3330
rect 306196 3266 306248 3272
rect 305000 3188 305052 3194
rect 305000 3130 305052 3136
rect 305012 480 305040 3130
rect 306208 480 306236 3266
rect 307404 480 307432 4082
rect 307588 2990 307616 102054
rect 307680 3330 307708 102068
rect 308522 102054 309088 102082
rect 308588 3936 308640 3942
rect 308588 3878 308640 3884
rect 307668 3324 307720 3330
rect 307668 3266 307720 3272
rect 307576 2984 307628 2990
rect 307576 2926 307628 2932
rect 308600 480 308628 3878
rect 309060 3058 309088 102054
rect 309428 100706 309456 102068
rect 310164 102054 310270 102082
rect 311098 102054 311848 102082
rect 309416 100700 309468 100706
rect 309416 100642 309468 100648
rect 310164 96665 310192 102054
rect 310428 100700 310480 100706
rect 310428 100642 310480 100648
rect 310150 96656 310206 96665
rect 310150 96591 310206 96600
rect 310334 96656 310390 96665
rect 310334 96591 310390 96600
rect 310348 89706 310376 96591
rect 310164 89678 310376 89706
rect 310164 86970 310192 89678
rect 310152 86964 310204 86970
rect 310152 86906 310204 86912
rect 310244 80028 310296 80034
rect 310244 79970 310296 79976
rect 310256 66434 310284 79970
rect 310060 66428 310112 66434
rect 310060 66370 310112 66376
rect 310244 66428 310296 66434
rect 310244 66370 310296 66376
rect 310072 63510 310100 66370
rect 310060 63504 310112 63510
rect 310060 63446 310112 63452
rect 310244 59220 310296 59226
rect 310244 59162 310296 59168
rect 310256 45642 310284 59162
rect 310072 45614 310284 45642
rect 310072 45558 310100 45614
rect 310060 45552 310112 45558
rect 310060 45494 310112 45500
rect 310244 40724 310296 40730
rect 310244 40666 310296 40672
rect 310256 31822 310284 40666
rect 310244 31816 310296 31822
rect 310244 31758 310296 31764
rect 310152 31748 310204 31754
rect 310152 31690 310204 31696
rect 310164 27554 310192 31690
rect 310072 27538 310192 27554
rect 310060 27532 310192 27538
rect 310112 27526 310192 27532
rect 310060 27474 310112 27480
rect 310336 12368 310388 12374
rect 310336 12310 310388 12316
rect 310348 9602 310376 12310
rect 310256 9574 310376 9602
rect 310256 4894 310284 9574
rect 310244 4888 310296 4894
rect 310244 4830 310296 4836
rect 309784 4004 309836 4010
rect 309784 3946 309836 3952
rect 309048 3052 309100 3058
rect 309048 2994 309100 3000
rect 309796 480 309824 3946
rect 310440 2718 310468 100642
rect 310980 4072 311032 4078
rect 310980 4014 311032 4020
rect 310428 2712 310480 2718
rect 310428 2654 310480 2660
rect 310992 480 311020 4014
rect 311820 3942 311848 102054
rect 311912 100706 311940 102068
rect 312846 102054 313228 102082
rect 311900 100700 311952 100706
rect 311900 100642 311952 100648
rect 313096 100700 313148 100706
rect 313096 100642 313148 100648
rect 313108 4010 313136 100642
rect 313096 4004 313148 4010
rect 313096 3946 313148 3952
rect 311808 3936 311860 3942
rect 311808 3878 311860 3884
rect 313200 3602 313228 102054
rect 313660 100706 313688 102068
rect 313648 100700 313700 100706
rect 313648 100642 313700 100648
rect 313188 3596 313240 3602
rect 313188 3538 313240 3544
rect 312176 3528 312228 3534
rect 312176 3470 312228 3476
rect 312188 480 312216 3470
rect 314488 3466 314516 102068
rect 315422 102054 315988 102082
rect 314568 100700 314620 100706
rect 314568 100642 314620 100648
rect 314580 4078 314608 100642
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 315960 3534 315988 102054
rect 316236 100706 316264 102068
rect 317078 102054 317368 102082
rect 316224 100700 316276 100706
rect 316224 100642 316276 100648
rect 317236 100700 317288 100706
rect 317236 100642 317288 100648
rect 317248 4758 317276 100642
rect 317236 4752 317288 4758
rect 317236 4694 317288 4700
rect 317340 3806 317368 102054
rect 317892 100706 317920 102068
rect 317880 100700 317932 100706
rect 317880 100642 317932 100648
rect 318708 100700 318760 100706
rect 318708 100642 318760 100648
rect 318064 4888 318116 4894
rect 318064 4830 318116 4836
rect 317328 3800 317380 3806
rect 317328 3742 317380 3748
rect 315948 3528 316000 3534
rect 315948 3470 316000 3476
rect 314476 3460 314528 3466
rect 314476 3402 314528 3408
rect 314568 3324 314620 3330
rect 314568 3266 314620 3272
rect 313372 2984 313424 2990
rect 313372 2926 313424 2932
rect 313384 480 313412 2926
rect 314580 480 314608 3266
rect 315764 3052 315816 3058
rect 315764 2994 315816 3000
rect 315776 480 315804 2994
rect 316960 2712 317012 2718
rect 316960 2654 317012 2660
rect 316972 480 317000 2654
rect 318076 480 318104 4830
rect 318720 3738 318748 100642
rect 318812 99482 318840 102068
rect 319654 102054 320128 102082
rect 318800 99476 318852 99482
rect 318800 99418 318852 99424
rect 319260 3936 319312 3942
rect 319260 3878 319312 3884
rect 318708 3732 318760 3738
rect 318708 3674 318760 3680
rect 319272 480 319300 3878
rect 320100 3670 320128 102054
rect 320468 95334 320496 102068
rect 321204 102054 321310 102082
rect 322230 102054 322888 102082
rect 320456 95328 320508 95334
rect 320456 95270 320508 95276
rect 321204 95266 321232 102054
rect 321468 95328 321520 95334
rect 321468 95270 321520 95276
rect 321192 95260 321244 95266
rect 321192 95202 321244 95208
rect 321376 95260 321428 95266
rect 321376 95202 321428 95208
rect 321388 95146 321416 95202
rect 321204 95118 321416 95146
rect 321204 85610 321232 95118
rect 321192 85604 321244 85610
rect 321192 85546 321244 85552
rect 321284 85604 321336 85610
rect 321284 85546 321336 85552
rect 321296 80730 321324 85546
rect 321204 80702 321324 80730
rect 321204 71126 321232 80702
rect 321192 71120 321244 71126
rect 321192 71062 321244 71068
rect 321376 71120 321428 71126
rect 321376 71062 321428 71068
rect 321388 66337 321416 71062
rect 321190 66328 321246 66337
rect 321112 66286 321190 66314
rect 321112 64870 321140 66286
rect 321190 66263 321246 66272
rect 321374 66328 321430 66337
rect 321374 66263 321430 66272
rect 321100 64864 321152 64870
rect 321100 64806 321152 64812
rect 321192 55276 321244 55282
rect 321192 55218 321244 55224
rect 321204 51134 321232 55218
rect 321192 51128 321244 51134
rect 321192 51070 321244 51076
rect 321100 51060 321152 51066
rect 321100 51002 321152 51008
rect 321112 46866 321140 51002
rect 321190 46880 321246 46889
rect 321112 46838 321190 46866
rect 321190 46815 321246 46824
rect 321190 37360 321246 37369
rect 321190 37295 321246 37304
rect 321204 37262 321232 37295
rect 321192 37256 321244 37262
rect 321192 37198 321244 37204
rect 321100 27668 321152 27674
rect 321100 27610 321152 27616
rect 321112 22166 321140 27610
rect 321100 22160 321152 22166
rect 321100 22102 321152 22108
rect 321100 18012 321152 18018
rect 321100 17954 321152 17960
rect 321112 9586 321140 17954
rect 321100 9580 321152 9586
rect 321100 9522 321152 9528
rect 321480 4010 321508 95270
rect 322860 4162 322888 102054
rect 323044 100706 323072 102068
rect 323886 102054 324176 102082
rect 323032 100700 323084 100706
rect 323032 100642 323084 100648
rect 324148 7614 324176 102054
rect 324792 100706 324820 102068
rect 324228 100700 324280 100706
rect 324228 100642 324280 100648
rect 324780 100700 324832 100706
rect 324780 100642 324832 100648
rect 325516 100700 325568 100706
rect 325516 100642 325568 100648
rect 324136 7608 324188 7614
rect 324136 7550 324188 7556
rect 322860 4134 322980 4162
rect 322848 4072 322900 4078
rect 322848 4014 322900 4020
rect 320456 4004 320508 4010
rect 320456 3946 320508 3952
rect 321468 4004 321520 4010
rect 321468 3946 321520 3952
rect 320088 3664 320140 3670
rect 320088 3606 320140 3612
rect 320468 480 320496 3946
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 321664 480 321692 3538
rect 322860 480 322888 4014
rect 322952 3602 322980 4134
rect 324240 3942 324268 100642
rect 324228 3936 324280 3942
rect 324228 3878 324280 3884
rect 322940 3596 322992 3602
rect 322940 3538 322992 3544
rect 325528 3534 325556 100642
rect 325240 3528 325292 3534
rect 325240 3470 325292 3476
rect 325516 3528 325568 3534
rect 325516 3470 325568 3476
rect 324044 3460 324096 3466
rect 324044 3402 324096 3408
rect 324056 480 324084 3402
rect 325252 480 325280 3470
rect 325620 3466 325648 102068
rect 326448 100026 326476 102068
rect 327276 100706 327304 102068
rect 328104 102054 328210 102082
rect 327264 100700 327316 100706
rect 327264 100642 327316 100648
rect 326436 100020 326488 100026
rect 326436 99962 326488 99968
rect 326344 99476 326396 99482
rect 326344 99418 326396 99424
rect 326356 5506 326384 99418
rect 328104 96665 328132 102054
rect 329024 100706 329052 102068
rect 329852 100706 329880 102068
rect 330786 102054 331168 102082
rect 328368 100700 328420 100706
rect 328368 100642 328420 100648
rect 329012 100700 329064 100706
rect 329012 100642 329064 100648
rect 329748 100700 329800 100706
rect 329748 100642 329800 100648
rect 329840 100700 329892 100706
rect 329840 100642 329892 100648
rect 331036 100700 331088 100706
rect 331036 100642 331088 100648
rect 328090 96656 328146 96665
rect 328274 96656 328330 96665
rect 328090 96591 328146 96600
rect 328184 96620 328236 96626
rect 328274 96591 328276 96600
rect 328184 96562 328236 96568
rect 328328 96591 328330 96600
rect 328276 96562 328328 96568
rect 328196 87009 328224 96562
rect 327998 87000 328054 87009
rect 327998 86935 328054 86944
rect 328182 87000 328238 87009
rect 328182 86935 328238 86944
rect 328012 80102 328040 86935
rect 328000 80096 328052 80102
rect 328000 80038 328052 80044
rect 328092 79960 328144 79966
rect 328092 79902 328144 79908
rect 328104 75886 328132 79902
rect 328092 75880 328144 75886
rect 328092 75822 328144 75828
rect 328000 66292 328052 66298
rect 328000 66234 328052 66240
rect 328012 66162 328040 66234
rect 328000 66156 328052 66162
rect 328000 66098 328052 66104
rect 328000 56636 328052 56642
rect 328000 56578 328052 56584
rect 328012 51082 328040 56578
rect 327920 51054 328040 51082
rect 327920 47054 327948 51054
rect 327908 47048 327960 47054
rect 327908 46990 327960 46996
rect 328000 47048 328052 47054
rect 328000 46990 328052 46996
rect 328012 45558 328040 46990
rect 328000 45552 328052 45558
rect 328000 45494 328052 45500
rect 328092 45552 328144 45558
rect 328092 45494 328144 45500
rect 328104 31754 328132 45494
rect 328092 31748 328144 31754
rect 328092 31690 328144 31696
rect 327908 26376 327960 26382
rect 327908 26318 327960 26324
rect 327920 26246 327948 26318
rect 327908 26240 327960 26246
rect 327908 26182 327960 26188
rect 328092 21956 328144 21962
rect 328092 21898 328144 21904
rect 328104 9790 328132 21898
rect 328092 9784 328144 9790
rect 328092 9726 328144 9732
rect 328092 9648 328144 9654
rect 328092 9590 328144 9596
rect 326344 5500 326396 5506
rect 326344 5442 326396 5448
rect 326436 4752 326488 4758
rect 326436 4694 326488 4700
rect 325608 3460 325660 3466
rect 325608 3402 325660 3408
rect 326448 480 326476 4694
rect 328104 3806 328132 9590
rect 328380 3874 328408 100642
rect 329760 10334 329788 100642
rect 331048 11762 331076 100642
rect 331036 11756 331088 11762
rect 331036 11698 331088 11704
rect 329748 10328 329800 10334
rect 329748 10270 329800 10276
rect 330024 5500 330076 5506
rect 330024 5442 330076 5448
rect 328368 3868 328420 3874
rect 328368 3810 328420 3816
rect 327632 3800 327684 3806
rect 327632 3742 327684 3748
rect 328092 3800 328144 3806
rect 328092 3742 328144 3748
rect 327644 480 327672 3742
rect 328828 3732 328880 3738
rect 328828 3674 328880 3680
rect 328840 480 328868 3674
rect 330036 480 330064 5442
rect 331140 3738 331168 102054
rect 331600 100706 331628 102068
rect 332336 102054 332442 102082
rect 333270 102054 333928 102082
rect 331588 100700 331640 100706
rect 331588 100642 331640 100648
rect 332336 96665 332364 102054
rect 333244 100700 333296 100706
rect 333244 100642 333296 100648
rect 332322 96656 332378 96665
rect 332322 96591 332378 96600
rect 332506 96656 332562 96665
rect 332506 96591 332562 96600
rect 332520 89758 332548 96591
rect 332324 89752 332376 89758
rect 332508 89752 332560 89758
rect 332376 89700 332508 89706
rect 332324 89694 332560 89700
rect 332336 89678 332548 89694
rect 332520 80102 332548 89678
rect 332508 80096 332560 80102
rect 332508 80038 332560 80044
rect 332416 80028 332468 80034
rect 332416 79970 332468 79976
rect 332428 72486 332456 79970
rect 332416 72480 332468 72486
rect 332416 72422 332468 72428
rect 332600 72480 332652 72486
rect 332600 72422 332652 72428
rect 332612 67697 332640 72422
rect 332414 67688 332470 67697
rect 332336 67646 332414 67674
rect 332336 66230 332364 67646
rect 332414 67623 332470 67632
rect 332598 67688 332654 67697
rect 332598 67623 332654 67632
rect 332324 66224 332376 66230
rect 332324 66166 332376 66172
rect 332416 56636 332468 56642
rect 332416 56578 332468 56584
rect 332428 48414 332456 56578
rect 332416 48408 332468 48414
rect 332416 48350 332468 48356
rect 332324 46980 332376 46986
rect 332324 46922 332376 46928
rect 332336 46850 332364 46922
rect 332324 46844 332376 46850
rect 332324 46786 332376 46792
rect 332416 46844 332468 46850
rect 332416 46786 332468 46792
rect 332428 31822 332456 46786
rect 332416 31816 332468 31822
rect 332416 31758 332468 31764
rect 332324 31748 332376 31754
rect 332324 31690 332376 31696
rect 332336 22166 332364 31690
rect 332324 22160 332376 22166
rect 332324 22102 332376 22108
rect 332324 22024 332376 22030
rect 332324 21966 332376 21972
rect 332336 13122 332364 21966
rect 332324 13116 332376 13122
rect 332324 13058 332376 13064
rect 333256 6186 333284 100642
rect 333244 6180 333296 6186
rect 333244 6122 333296 6128
rect 333612 6044 333664 6050
rect 333612 5986 333664 5992
rect 332416 4004 332468 4010
rect 332416 3946 332468 3952
rect 331128 3732 331180 3738
rect 331128 3674 331180 3680
rect 331220 3664 331272 3670
rect 331220 3606 331272 3612
rect 331232 480 331260 3606
rect 332428 480 332456 3946
rect 333624 480 333652 5986
rect 333900 3670 333928 102054
rect 334176 100706 334204 102068
rect 335018 102054 335216 102082
rect 334164 100700 334216 100706
rect 334164 100642 334216 100648
rect 335188 15910 335216 102054
rect 335832 100706 335860 102068
rect 335268 100700 335320 100706
rect 335268 100642 335320 100648
rect 335820 100700 335872 100706
rect 335820 100642 335872 100648
rect 336556 100700 336608 100706
rect 336556 100642 336608 100648
rect 335176 15904 335228 15910
rect 335176 15846 335228 15852
rect 335280 4826 335308 100642
rect 335268 4820 335320 4826
rect 335268 4762 335320 4768
rect 335912 3936 335964 3942
rect 335912 3878 335964 3884
rect 333888 3664 333940 3670
rect 333888 3606 333940 3612
rect 334716 3596 334768 3602
rect 334716 3538 334768 3544
rect 334728 480 334756 3538
rect 335924 480 335952 3878
rect 336568 3602 336596 100642
rect 336660 98666 336688 102068
rect 337580 100162 337608 102068
rect 338408 100706 338436 102068
rect 338396 100700 338448 100706
rect 338396 100642 338448 100648
rect 337568 100156 337620 100162
rect 337568 100098 337620 100104
rect 338764 100156 338816 100162
rect 338764 100098 338816 100104
rect 337384 100020 337436 100026
rect 337384 99962 337436 99968
rect 336648 98660 336700 98666
rect 336648 98602 336700 98608
rect 337396 8566 337424 99962
rect 338776 8974 338804 100098
rect 339236 99550 339264 102068
rect 340170 102054 340828 102082
rect 339408 100700 339460 100706
rect 339408 100642 339460 100648
rect 339224 99544 339276 99550
rect 339224 99486 339276 99492
rect 338764 8968 338816 8974
rect 338764 8910 338816 8916
rect 337384 8560 337436 8566
rect 337384 8502 337436 8508
rect 337108 7608 337160 7614
rect 337108 7550 337160 7556
rect 336556 3596 336608 3602
rect 336556 3538 336608 3544
rect 337120 480 337148 7550
rect 339420 3534 339448 100642
rect 340800 17270 340828 102054
rect 340984 100638 341012 102068
rect 341826 102054 342116 102082
rect 340972 100632 341024 100638
rect 340972 100574 341024 100580
rect 342088 73846 342116 102054
rect 342640 100638 342668 102068
rect 342168 100632 342220 100638
rect 342168 100574 342220 100580
rect 342628 100632 342680 100638
rect 342628 100574 342680 100580
rect 342076 73840 342128 73846
rect 342076 73782 342128 73788
rect 340788 17264 340840 17270
rect 340788 17206 340840 17212
rect 340696 8560 340748 8566
rect 340696 8502 340748 8508
rect 338304 3528 338356 3534
rect 338304 3470 338356 3476
rect 339408 3528 339460 3534
rect 339408 3470 339460 3476
rect 338316 480 338344 3470
rect 339500 3460 339552 3466
rect 339500 3402 339552 3408
rect 339512 480 339540 3402
rect 340708 480 340736 8502
rect 341892 3868 341944 3874
rect 341892 3810 341944 3816
rect 341904 480 341932 3810
rect 342180 3466 342208 100574
rect 343560 3942 343588 102068
rect 344402 102054 344968 102082
rect 344284 99544 344336 99550
rect 344284 99486 344336 99492
rect 344296 14482 344324 99486
rect 344284 14476 344336 14482
rect 344284 14418 344336 14424
rect 343640 10328 343692 10334
rect 343640 10270 343692 10276
rect 343548 3936 343600 3942
rect 343548 3878 343600 3884
rect 343088 3800 343140 3806
rect 343088 3742 343140 3748
rect 342168 3460 342220 3466
rect 342168 3402 342220 3408
rect 343100 480 343128 3742
rect 343652 3346 343680 10270
rect 344940 7614 344968 102054
rect 345216 100706 345244 102068
rect 346150 102054 346348 102082
rect 345204 100700 345256 100706
rect 345204 100642 345256 100648
rect 346216 100700 346268 100706
rect 346216 100642 346268 100648
rect 346228 18630 346256 100642
rect 346216 18624 346268 18630
rect 346216 18566 346268 18572
rect 345020 11756 345072 11762
rect 345020 11698 345072 11704
rect 344928 7608 344980 7614
rect 344928 7550 344980 7556
rect 343652 3318 344324 3346
rect 344296 480 344324 3318
rect 345032 626 345060 11698
rect 346320 4010 346348 102054
rect 346964 100026 346992 102068
rect 347792 100638 347820 102068
rect 348634 102054 349108 102082
rect 347044 100632 347096 100638
rect 347044 100574 347096 100580
rect 347780 100632 347832 100638
rect 347780 100574 347832 100580
rect 348976 100632 349028 100638
rect 348976 100574 349028 100580
rect 346952 100020 347004 100026
rect 346952 99962 347004 99968
rect 347056 11762 347084 100574
rect 348988 21418 349016 100574
rect 348976 21412 349028 21418
rect 348976 21354 349028 21360
rect 347780 13116 347832 13122
rect 347780 13058 347832 13064
rect 347044 11756 347096 11762
rect 347044 11698 347096 11704
rect 346308 4004 346360 4010
rect 346308 3946 346360 3952
rect 346676 3732 346728 3738
rect 346676 3674 346728 3680
rect 345032 598 345520 626
rect 345492 480 345520 598
rect 346688 480 346716 3674
rect 347792 3602 347820 13058
rect 347872 6180 347924 6186
rect 347872 6122 347924 6128
rect 347780 3596 347832 3602
rect 347780 3538 347832 3544
rect 347884 480 347912 6122
rect 349080 3874 349108 102054
rect 349540 97306 349568 102068
rect 349528 97300 349580 97306
rect 349528 97242 349580 97248
rect 350552 96642 350580 102190
rect 356900 102190 357190 102218
rect 468772 102190 469062 102218
rect 351210 102054 351868 102082
rect 350460 96614 350580 96642
rect 350460 87009 350488 96614
rect 350262 87000 350318 87009
rect 350262 86935 350318 86944
rect 350446 87000 350502 87009
rect 350446 86935 350502 86944
rect 350276 80170 350304 86935
rect 350264 80164 350316 80170
rect 350264 80106 350316 80112
rect 350172 75948 350224 75954
rect 350172 75890 350224 75896
rect 350184 67658 350212 75890
rect 350172 67652 350224 67658
rect 350172 67594 350224 67600
rect 350356 67652 350408 67658
rect 350356 67594 350408 67600
rect 350368 66230 350396 67594
rect 350356 66224 350408 66230
rect 350356 66166 350408 66172
rect 350356 63912 350408 63918
rect 350356 63854 350408 63860
rect 350368 54097 350396 63854
rect 350354 54088 350410 54097
rect 350354 54023 350410 54032
rect 350354 53952 350410 53961
rect 350354 53887 350410 53896
rect 350368 53825 350396 53887
rect 350354 53816 350410 53825
rect 350354 53751 350410 53760
rect 350538 53816 350594 53825
rect 350538 53751 350594 53760
rect 350552 44266 350580 53751
rect 350356 44260 350408 44266
rect 350356 44202 350408 44208
rect 350540 44260 350592 44266
rect 350540 44202 350592 44208
rect 350368 44130 350396 44202
rect 350356 44124 350408 44130
rect 350356 44066 350408 44072
rect 350356 31680 350408 31686
rect 350356 31622 350408 31628
rect 350368 16658 350396 31622
rect 350264 16652 350316 16658
rect 350264 16594 350316 16600
rect 350356 16652 350408 16658
rect 350356 16594 350408 16600
rect 350276 13122 350304 16594
rect 350264 13116 350316 13122
rect 350264 13058 350316 13064
rect 351368 4820 351420 4826
rect 351368 4762 351420 4768
rect 349068 3868 349120 3874
rect 349068 3810 349120 3816
rect 350264 3664 350316 3670
rect 350264 3606 350316 3612
rect 349068 3596 349120 3602
rect 349068 3538 349120 3544
rect 349080 480 349108 3538
rect 350276 480 350304 3606
rect 351380 480 351408 4762
rect 351840 3806 351868 102054
rect 352024 100638 352052 102068
rect 352958 102054 353156 102082
rect 352012 100632 352064 100638
rect 352012 100574 352064 100580
rect 353128 22778 353156 102054
rect 353772 100706 353800 102068
rect 354508 102054 354614 102082
rect 355534 102054 356008 102082
rect 353760 100700 353812 100706
rect 353760 100642 353812 100648
rect 353208 100632 353260 100638
rect 353208 100574 353260 100580
rect 353116 22772 353168 22778
rect 353116 22714 353168 22720
rect 351920 15904 351972 15910
rect 351920 15846 351972 15852
rect 351828 3800 351880 3806
rect 351828 3742 351880 3748
rect 351932 610 351960 15846
rect 353220 4826 353248 100574
rect 354508 95946 354536 102054
rect 354588 100700 354640 100706
rect 354588 100642 354640 100648
rect 354496 95940 354548 95946
rect 354496 95882 354548 95888
rect 353208 4820 353260 4826
rect 353208 4762 353260 4768
rect 354600 3738 354628 100642
rect 354680 98660 354732 98666
rect 354680 98602 354732 98608
rect 354588 3732 354640 3738
rect 354588 3674 354640 3680
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 351920 604 351972 610
rect 351920 546 351972 552
rect 352564 604 352616 610
rect 352564 546 352616 552
rect 352576 480 352604 546
rect 353772 480 353800 3334
rect 354692 1034 354720 98602
rect 355980 15910 356008 102054
rect 356348 100706 356376 102068
rect 356336 100700 356388 100706
rect 356336 100642 356388 100648
rect 356900 96694 356928 102190
rect 358018 102054 358768 102082
rect 357348 100700 357400 100706
rect 357348 100642 357400 100648
rect 356888 96688 356940 96694
rect 356888 96630 356940 96636
rect 356980 96688 357032 96694
rect 356980 96630 357032 96636
rect 356992 89706 357020 96630
rect 356992 89678 357112 89706
rect 357084 80238 357112 89678
rect 357072 80232 357124 80238
rect 357072 80174 357124 80180
rect 357072 80028 357124 80034
rect 357072 79970 357124 79976
rect 357084 67674 357112 79970
rect 356992 67646 357112 67674
rect 356992 66230 357020 67646
rect 356980 66224 357032 66230
rect 356980 66166 357032 66172
rect 357072 56636 357124 56642
rect 357072 56578 357124 56584
rect 357084 50946 357112 56578
rect 356992 50918 357112 50946
rect 356992 41478 357020 50918
rect 356980 41472 357032 41478
rect 356980 41414 357032 41420
rect 357072 41336 357124 41342
rect 357072 41278 357124 41284
rect 357084 37262 357112 41278
rect 357072 37256 357124 37262
rect 357072 37198 357124 37204
rect 357072 31748 357124 31754
rect 357072 31690 357124 31696
rect 357084 27690 357112 31690
rect 357084 27662 357204 27690
rect 357176 27606 357204 27662
rect 357164 27600 357216 27606
rect 357164 27542 357216 27548
rect 357256 18012 357308 18018
rect 357256 17954 357308 17960
rect 355968 15904 356020 15910
rect 355968 15846 356020 15852
rect 357268 12458 357296 17954
rect 357176 12430 357296 12458
rect 356152 8968 356204 8974
rect 356152 8910 356204 8916
rect 354692 1006 354996 1034
rect 354968 480 354996 1006
rect 356164 480 356192 8910
rect 357176 6186 357204 12430
rect 357164 6180 357216 6186
rect 357164 6122 357216 6128
rect 357360 3670 357388 100642
rect 358740 14482 358768 102054
rect 358924 99890 358952 102068
rect 359766 102054 360056 102082
rect 358912 99884 358964 99890
rect 358912 99826 358964 99832
rect 358820 17264 358872 17270
rect 358820 17206 358872 17212
rect 357440 14476 357492 14482
rect 357440 14418 357492 14424
rect 358728 14476 358780 14482
rect 358728 14418 358780 14424
rect 357452 9654 357480 14418
rect 358832 9654 358860 17206
rect 357440 9648 357492 9654
rect 357440 9590 357492 9596
rect 358820 9648 358872 9654
rect 358820 9590 358872 9596
rect 360028 8974 360056 102054
rect 360580 100094 360608 102068
rect 360568 100088 360620 100094
rect 360568 100030 360620 100036
rect 360108 99884 360160 99890
rect 360108 99826 360160 99832
rect 360016 8968 360068 8974
rect 360016 8910 360068 8916
rect 360120 3670 360148 99826
rect 357348 3664 357400 3670
rect 357348 3606 357400 3612
rect 360108 3664 360160 3670
rect 360108 3606 360160 3612
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 357360 480 357388 3470
rect 361500 3466 361528 102068
rect 362342 102054 362908 102082
rect 361580 73840 361632 73846
rect 361580 73782 361632 73788
rect 360936 3460 360988 3466
rect 360936 3402 360988 3408
rect 361488 3460 361540 3466
rect 361488 3402 361540 3408
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 358556 480 358584 546
rect 359752 480 359780 546
rect 360948 480 360976 3402
rect 361592 3210 361620 73782
rect 362880 10334 362908 102054
rect 363156 99414 363184 102068
rect 363998 102054 364288 102082
rect 363144 99408 363196 99414
rect 363144 99350 363196 99356
rect 364156 99408 364208 99414
rect 364156 99350 364208 99356
rect 364168 17270 364196 99350
rect 364156 17264 364208 17270
rect 364156 17206 364208 17212
rect 362960 11756 363012 11762
rect 362960 11698 363012 11704
rect 362868 10328 362920 10334
rect 362868 10270 362920 10276
rect 362972 3210 363000 11698
rect 364260 3534 364288 102054
rect 364904 99414 364932 102068
rect 365732 99414 365760 102068
rect 366574 102054 366956 102082
rect 364892 99408 364944 99414
rect 364892 99350 364944 99356
rect 365628 99408 365680 99414
rect 365628 99350 365680 99356
rect 365720 99408 365772 99414
rect 365720 99350 365772 99356
rect 365640 11762 365668 99350
rect 366928 32502 366956 102054
rect 367008 99408 367060 99414
rect 367008 99350 367060 99356
rect 366916 32496 366968 32502
rect 366916 32438 366968 32444
rect 367020 18630 367048 99350
rect 367480 98666 367508 102068
rect 367468 98660 367520 98666
rect 367468 98602 367520 98608
rect 368308 24138 368336 102068
rect 369150 102054 369808 102082
rect 368572 100020 368624 100026
rect 368572 99962 368624 99968
rect 368296 24132 368348 24138
rect 368296 24074 368348 24080
rect 365720 18624 365772 18630
rect 365720 18566 365772 18572
rect 367008 18624 367060 18630
rect 367008 18566 367060 18572
rect 365628 11756 365680 11762
rect 365628 11698 365680 11704
rect 364524 3936 364576 3942
rect 364524 3878 364576 3884
rect 364248 3528 364300 3534
rect 364248 3470 364300 3476
rect 361592 3182 362172 3210
rect 362972 3182 363368 3210
rect 362144 480 362172 3182
rect 363340 480 363368 3182
rect 364536 480 364564 3878
rect 365732 3874 365760 18566
rect 365812 7608 365864 7614
rect 365812 7550 365864 7556
rect 365720 3868 365772 3874
rect 365720 3810 365772 3816
rect 365824 3482 365852 7550
rect 368020 4004 368072 4010
rect 368020 3946 368072 3952
rect 366916 3868 366968 3874
rect 366916 3810 366968 3816
rect 365732 3454 365852 3482
rect 365732 480 365760 3454
rect 366928 480 366956 3810
rect 368032 480 368060 3946
rect 368584 3482 368612 99962
rect 369780 36650 369808 102054
rect 369964 100570 369992 102068
rect 370898 102054 371188 102082
rect 369952 100564 370004 100570
rect 369952 100506 370004 100512
rect 370504 100088 370556 100094
rect 370504 100030 370556 100036
rect 369768 36644 369820 36650
rect 369768 36586 369820 36592
rect 369860 21412 369912 21418
rect 369860 21354 369912 21360
rect 369872 3482 369900 21354
rect 370516 19990 370544 100030
rect 371160 21418 371188 102054
rect 371712 100638 371740 102068
rect 372540 100722 372568 102068
rect 373382 102054 373948 102082
rect 372540 100694 372660 100722
rect 371700 100632 371752 100638
rect 371700 100574 371752 100580
rect 372528 100632 372580 100638
rect 372528 100574 372580 100580
rect 372540 37942 372568 100574
rect 372632 97374 372660 100694
rect 372620 97368 372672 97374
rect 372620 97310 372672 97316
rect 372620 97232 372672 97238
rect 372620 97174 372672 97180
rect 372528 37936 372580 37942
rect 372528 37878 372580 37884
rect 371148 21412 371200 21418
rect 371148 21354 371200 21360
rect 370504 19984 370556 19990
rect 370504 19926 370556 19932
rect 371608 3936 371660 3942
rect 371608 3878 371660 3884
rect 368584 3454 369256 3482
rect 369872 3454 370452 3482
rect 369228 480 369256 3454
rect 370424 480 370452 3454
rect 371620 480 371648 3878
rect 372632 3482 372660 97174
rect 373920 25566 373948 102054
rect 374288 100706 374316 102068
rect 375130 102054 375328 102082
rect 374276 100700 374328 100706
rect 374276 100642 374328 100648
rect 375196 100700 375248 100706
rect 375196 100642 375248 100648
rect 375208 42090 375236 100642
rect 375196 42084 375248 42090
rect 375196 42026 375248 42032
rect 373908 25560 373960 25566
rect 373908 25502 373960 25508
rect 375300 13190 375328 102054
rect 375944 100026 375972 102068
rect 376024 100564 376076 100570
rect 376024 100506 376076 100512
rect 375932 100020 375984 100026
rect 375932 99962 375984 99968
rect 375288 13184 375340 13190
rect 375288 13126 375340 13132
rect 374092 13116 374144 13122
rect 374092 13058 374144 13064
rect 372632 3454 372844 3482
rect 372816 480 372844 3454
rect 374104 1442 374132 13058
rect 376036 4894 376064 100506
rect 376864 99686 376892 102068
rect 377692 100026 377720 102068
rect 377404 100020 377456 100026
rect 377404 99962 377456 99968
rect 377680 100020 377732 100026
rect 377680 99962 377732 99968
rect 376852 99680 376904 99686
rect 376852 99622 376904 99628
rect 377416 22778 377444 99962
rect 378048 99680 378100 99686
rect 378048 99622 378100 99628
rect 378060 44878 378088 99622
rect 378520 94518 378548 102068
rect 379256 102054 379362 102082
rect 380282 102054 380848 102082
rect 379256 96665 379284 102054
rect 379242 96656 379298 96665
rect 379242 96591 379298 96600
rect 379426 96656 379482 96665
rect 379426 96591 379482 96600
rect 378508 94512 378560 94518
rect 378508 94454 378560 94460
rect 379440 89758 379468 96591
rect 379520 95940 379572 95946
rect 379520 95882 379572 95888
rect 379244 89752 379296 89758
rect 379428 89752 379480 89758
rect 379296 89700 379376 89706
rect 379244 89694 379376 89700
rect 379428 89694 379480 89700
rect 379256 89678 379376 89694
rect 379348 80170 379376 89678
rect 379336 80164 379388 80170
rect 379336 80106 379388 80112
rect 379336 80028 379388 80034
rect 379336 79970 379388 79976
rect 379348 70394 379376 79970
rect 379256 70366 379376 70394
rect 379256 70258 379284 70366
rect 379256 70230 379376 70258
rect 379348 51082 379376 70230
rect 379256 51054 379376 51082
rect 379256 47598 379284 51054
rect 379244 47592 379296 47598
rect 379244 47534 379296 47540
rect 378048 44872 378100 44878
rect 378048 44814 378100 44820
rect 376760 22772 376812 22778
rect 376760 22714 376812 22720
rect 377404 22772 377456 22778
rect 377404 22714 377456 22720
rect 376024 4888 376076 4894
rect 376024 4830 376076 4836
rect 376392 4820 376444 4826
rect 376392 4762 376444 4768
rect 375196 3800 375248 3806
rect 375196 3742 375248 3748
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3742
rect 376404 480 376432 4762
rect 376772 3346 376800 22714
rect 378784 3732 378836 3738
rect 378784 3674 378836 3680
rect 376772 3318 377628 3346
rect 377600 480 377628 3318
rect 378796 480 378824 3674
rect 379532 3346 379560 95882
rect 380820 7614 380848 102054
rect 381096 99890 381124 102068
rect 381938 102054 382136 102082
rect 382858 102054 383608 102082
rect 381084 99884 381136 99890
rect 381084 99826 381136 99832
rect 382108 49026 382136 102054
rect 382188 99884 382240 99890
rect 382188 99826 382240 99832
rect 382096 49020 382148 49026
rect 382096 48962 382148 48968
rect 382200 26926 382228 99826
rect 382188 26920 382240 26926
rect 382188 26862 382240 26868
rect 380900 15904 380952 15910
rect 380900 15846 380952 15852
rect 380808 7608 380860 7614
rect 380808 7550 380860 7556
rect 380912 3346 380940 15846
rect 383580 6186 383608 102054
rect 383672 100706 383700 102068
rect 384514 102054 384896 102082
rect 383660 100700 383712 100706
rect 383660 100642 383712 100648
rect 384868 51746 384896 102054
rect 384948 100700 385000 100706
rect 384948 100642 385000 100648
rect 384856 51740 384908 51746
rect 384856 51682 384908 51688
rect 384960 28286 384988 100642
rect 385328 95946 385356 102068
rect 386156 102054 386262 102082
rect 387090 102054 387748 102082
rect 386156 99346 386184 102054
rect 386144 99340 386196 99346
rect 386144 99282 386196 99288
rect 386328 99340 386380 99346
rect 386328 99282 386380 99288
rect 385316 95940 385368 95946
rect 385316 95882 385368 95888
rect 386340 75954 386368 99282
rect 386144 75948 386196 75954
rect 386144 75890 386196 75896
rect 386328 75948 386380 75954
rect 386328 75890 386380 75896
rect 386156 56030 386184 75890
rect 386144 56024 386196 56030
rect 386144 55966 386196 55972
rect 386328 48340 386380 48346
rect 386328 48282 386380 48288
rect 386340 41478 386368 48282
rect 386328 41472 386380 41478
rect 386328 41414 386380 41420
rect 386236 41404 386288 41410
rect 386236 41346 386288 41352
rect 386248 38622 386276 41346
rect 386236 38616 386288 38622
rect 386236 38558 386288 38564
rect 384948 28280 385000 28286
rect 384948 28222 385000 28228
rect 383660 14476 383712 14482
rect 383660 14418 383712 14424
rect 383476 6180 383528 6186
rect 383476 6122 383528 6128
rect 383568 6180 383620 6186
rect 383568 6122 383620 6128
rect 383488 6066 383516 6122
rect 383488 6038 383608 6066
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 379532 3318 380020 3346
rect 380912 3318 381216 3346
rect 379992 480 380020 3318
rect 381188 480 381216 3318
rect 382384 480 382412 3538
rect 383580 480 383608 6038
rect 383672 3482 383700 14418
rect 387064 8968 387116 8974
rect 387064 8910 387116 8916
rect 385868 3664 385920 3670
rect 385868 3606 385920 3612
rect 383672 3454 384712 3482
rect 384684 480 384712 3454
rect 385880 480 385908 3606
rect 387076 480 387104 8910
rect 387720 4826 387748 102054
rect 387904 100638 387932 102068
rect 388746 102054 389036 102082
rect 387892 100632 387944 100638
rect 387892 100574 387944 100580
rect 389008 31074 389036 102054
rect 389088 100632 389140 100638
rect 389088 100574 389140 100580
rect 388996 31068 389048 31074
rect 388996 31010 389048 31016
rect 387800 19984 387852 19990
rect 387800 19926 387852 19932
rect 387708 4820 387760 4826
rect 387708 4762 387760 4768
rect 387812 3482 387840 19926
rect 389100 8974 389128 100574
rect 389652 99414 389680 102068
rect 390480 99414 390508 102068
rect 391322 102054 391888 102082
rect 389640 99408 389692 99414
rect 389640 99350 389692 99356
rect 390468 99408 390520 99414
rect 390468 99350 390520 99356
rect 391204 99408 391256 99414
rect 391204 99350 391256 99356
rect 390468 99272 390520 99278
rect 390468 99214 390520 99220
rect 390480 93786 390508 99214
rect 390388 93758 390508 93786
rect 390388 89706 390416 93758
rect 390204 89678 390416 89706
rect 390204 82142 390232 89678
rect 390192 82136 390244 82142
rect 390192 82078 390244 82084
rect 390376 82136 390428 82142
rect 390376 82078 390428 82084
rect 390388 77353 390416 82078
rect 390190 77344 390246 77353
rect 390112 77302 390190 77330
rect 390112 62150 390140 77302
rect 390190 77279 390246 77288
rect 390374 77344 390430 77353
rect 390374 77279 390430 77288
rect 390008 62144 390060 62150
rect 390008 62086 390060 62092
rect 390100 62144 390152 62150
rect 390100 62086 390152 62092
rect 390020 60874 390048 62086
rect 390020 60846 390232 60874
rect 390204 52494 390232 60846
rect 391216 54534 391244 99350
rect 391204 54528 391256 54534
rect 391204 54470 391256 54476
rect 390192 52488 390244 52494
rect 390192 52430 390244 52436
rect 390284 52488 390336 52494
rect 390284 52430 390336 52436
rect 390296 48278 390324 52430
rect 390284 48272 390336 48278
rect 390284 48214 390336 48220
rect 390192 38684 390244 38690
rect 390192 38626 390244 38632
rect 390204 32434 390232 38626
rect 391860 33794 391888 102054
rect 392228 99414 392256 102068
rect 393070 102054 393268 102082
rect 393898 102054 394648 102082
rect 392216 99408 392268 99414
rect 392216 99350 392268 99356
rect 393136 99408 393188 99414
rect 393136 99350 393188 99356
rect 393148 57254 393176 99350
rect 393136 57248 393188 57254
rect 393136 57190 393188 57196
rect 391848 33788 391900 33794
rect 391848 33730 391900 33736
rect 390192 32428 390244 32434
rect 390192 32370 390244 32376
rect 390560 17264 390612 17270
rect 390560 17206 390612 17212
rect 389088 8968 389140 8974
rect 389088 8910 389140 8916
rect 390572 7682 390600 17206
rect 393240 10334 393268 102054
rect 394620 35222 394648 102054
rect 394712 99414 394740 102068
rect 395646 102054 396028 102082
rect 394700 99408 394752 99414
rect 394700 99350 394752 99356
rect 395896 99408 395948 99414
rect 395896 99350 395948 99356
rect 395908 58682 395936 99350
rect 395896 58676 395948 58682
rect 395896 58618 395948 58624
rect 394608 35216 394660 35222
rect 394608 35158 394660 35164
rect 396000 11762 396028 102054
rect 396460 99414 396488 102068
rect 397288 99482 397316 102068
rect 398222 102054 398788 102082
rect 397276 99476 397328 99482
rect 397276 99418 397328 99424
rect 396448 99408 396500 99414
rect 396448 99350 396500 99356
rect 397368 99408 397420 99414
rect 397368 99350 397420 99356
rect 397380 89010 397408 99350
rect 397460 98660 397512 98666
rect 397460 98602 397512 98608
rect 397368 89004 397420 89010
rect 397368 88946 397420 88952
rect 396080 32496 396132 32502
rect 396080 32438 396132 32444
rect 396092 12442 396120 32438
rect 397472 14498 397500 98602
rect 397472 14470 397592 14498
rect 398760 14482 398788 102054
rect 399036 99414 399064 102068
rect 399484 99476 399536 99482
rect 399484 99418 399536 99424
rect 399024 99408 399076 99414
rect 399024 99350 399076 99356
rect 399496 36582 399524 99418
rect 399864 98734 399892 102068
rect 400692 99414 400720 102068
rect 401612 99414 401640 102068
rect 402454 102054 402928 102082
rect 400036 99408 400088 99414
rect 400036 99350 400088 99356
rect 400680 99408 400732 99414
rect 400680 99350 400732 99356
rect 401508 99408 401560 99414
rect 401508 99350 401560 99356
rect 401600 99408 401652 99414
rect 401600 99350 401652 99356
rect 402796 99408 402848 99414
rect 402796 99350 402848 99356
rect 399852 98728 399904 98734
rect 399852 98670 399904 98676
rect 400048 90370 400076 99350
rect 400036 90364 400088 90370
rect 400036 90306 400088 90312
rect 400220 36644 400272 36650
rect 400220 36586 400272 36592
rect 399484 36576 399536 36582
rect 399484 36518 399536 36524
rect 398840 24132 398892 24138
rect 398840 24074 398892 24080
rect 396080 12436 396132 12442
rect 396080 12378 396132 12384
rect 396632 12436 396684 12442
rect 396632 12378 396684 12384
rect 394240 11756 394292 11762
rect 394240 11698 394292 11704
rect 395988 11756 396040 11762
rect 395988 11698 396040 11704
rect 390652 10328 390704 10334
rect 390652 10270 390704 10276
rect 393228 10328 393280 10334
rect 393228 10270 393280 10276
rect 390560 7676 390612 7682
rect 390560 7618 390612 7624
rect 387812 3454 388300 3482
rect 388272 480 388300 3454
rect 389456 3460 389508 3466
rect 389456 3402 389508 3408
rect 389468 480 389496 3402
rect 390664 480 390692 10270
rect 391848 7676 391900 7682
rect 391848 7618 391900 7624
rect 391860 480 391888 7618
rect 393044 3528 393096 3534
rect 393044 3470 393096 3476
rect 393056 480 393084 3470
rect 394252 480 394280 11698
rect 395436 9716 395488 9722
rect 395436 9658 395488 9664
rect 395448 480 395476 9658
rect 396644 480 396672 12378
rect 397564 12374 397592 14470
rect 398748 14476 398800 14482
rect 398748 14418 398800 14424
rect 398852 12510 398880 24074
rect 398840 12504 398892 12510
rect 398840 12446 398892 12452
rect 397552 12368 397604 12374
rect 397552 12310 397604 12316
rect 397828 12368 397880 12374
rect 397828 12310 397880 12316
rect 399024 12368 399076 12374
rect 399024 12310 399076 12316
rect 397840 9654 397868 12310
rect 399036 9654 399064 12310
rect 397828 9648 397880 9654
rect 397828 9590 397880 9596
rect 399024 9648 399076 9654
rect 399024 9590 399076 9596
rect 397828 9512 397880 9518
rect 397828 9454 397880 9460
rect 399024 9512 399076 9518
rect 399024 9454 399076 9460
rect 397840 480 397868 9454
rect 399036 480 399064 9454
rect 400232 480 400260 36586
rect 401520 15910 401548 99350
rect 402808 39370 402836 99350
rect 402796 39364 402848 39370
rect 402796 39306 402848 39312
rect 401600 21412 401652 21418
rect 401600 21354 401652 21360
rect 401508 15904 401560 15910
rect 401508 15846 401560 15852
rect 401612 12442 401640 21354
rect 401600 12436 401652 12442
rect 401600 12378 401652 12384
rect 402520 12436 402572 12442
rect 402520 12378 402572 12384
rect 401324 4888 401376 4894
rect 401324 4830 401376 4836
rect 401336 480 401364 4830
rect 402532 480 402560 12378
rect 402900 4146 402928 102054
rect 403268 99414 403296 102068
rect 404110 102054 404308 102082
rect 405030 102054 405688 102082
rect 403256 99408 403308 99414
rect 403256 99350 403308 99356
rect 404176 99408 404228 99414
rect 404176 99350 404228 99356
rect 402980 37936 403032 37942
rect 402980 37878 403032 37884
rect 402992 12510 403020 37878
rect 404188 17270 404216 99350
rect 404176 17264 404228 17270
rect 404176 17206 404228 17212
rect 404280 13122 404308 102054
rect 404360 97300 404412 97306
rect 404360 97242 404412 97248
rect 404268 13116 404320 13122
rect 404268 13058 404320 13064
rect 402980 12504 403032 12510
rect 402980 12446 403032 12452
rect 404372 12442 404400 97242
rect 404360 12436 404412 12442
rect 404360 12378 404412 12384
rect 404912 12436 404964 12442
rect 404912 12378 404964 12384
rect 403716 12368 403768 12374
rect 403716 12310 403768 12316
rect 403728 9654 403756 12310
rect 403716 9648 403768 9654
rect 403716 9590 403768 9596
rect 403716 9512 403768 9518
rect 403716 9454 403768 9460
rect 402888 4140 402940 4146
rect 402888 4082 402940 4088
rect 403728 480 403756 9454
rect 404924 480 404952 12378
rect 405660 4010 405688 102054
rect 405844 99414 405872 102068
rect 406686 102054 406976 102082
rect 405832 99408 405884 99414
rect 405832 99350 405884 99356
rect 406948 40730 406976 102054
rect 407028 99408 407080 99414
rect 407028 99350 407080 99356
rect 406936 40724 406988 40730
rect 406936 40666 406988 40672
rect 405740 25560 405792 25566
rect 405740 25502 405792 25508
rect 405752 14498 405780 25502
rect 407040 18630 407068 99350
rect 407592 95266 407620 102068
rect 408420 99414 408448 102068
rect 409262 102054 409828 102082
rect 408408 99408 408460 99414
rect 408408 99350 408460 99356
rect 409144 99408 409196 99414
rect 409144 99350 409196 99356
rect 407580 95260 407632 95266
rect 407580 95202 407632 95208
rect 408224 95260 408276 95266
rect 408224 95202 408276 95208
rect 408236 95130 408264 95202
rect 408224 95124 408276 95130
rect 408224 95066 408276 95072
rect 408224 85604 408276 85610
rect 408224 85546 408276 85552
rect 408236 76022 408264 85546
rect 408132 76016 408184 76022
rect 408132 75958 408184 75964
rect 408224 76016 408276 76022
rect 408224 75958 408276 75964
rect 408144 75886 408172 75958
rect 408132 75880 408184 75886
rect 408132 75822 408184 75828
rect 408224 66292 408276 66298
rect 408224 66234 408276 66240
rect 408236 60738 408264 66234
rect 408236 60710 408356 60738
rect 408328 45626 408356 60710
rect 408132 45620 408184 45626
rect 408132 45562 408184 45568
rect 408316 45620 408368 45626
rect 408316 45562 408368 45568
rect 407120 42084 407172 42090
rect 407120 42026 407172 42032
rect 407028 18624 407080 18630
rect 407028 18566 407080 18572
rect 405752 14470 405872 14498
rect 405844 12322 405872 14470
rect 407132 12424 407160 42026
rect 408144 32314 408172 45562
rect 408144 32286 408264 32314
rect 408236 27606 408264 32286
rect 408224 27600 408276 27606
rect 408224 27542 408276 27548
rect 408500 22772 408552 22778
rect 408500 22714 408552 22720
rect 408408 18012 408460 18018
rect 408408 17954 408460 17960
rect 408420 16862 408448 17954
rect 408408 16856 408460 16862
rect 408408 16798 408460 16804
rect 407132 12396 407344 12424
rect 405844 12294 406148 12322
rect 406120 9654 406148 12294
rect 407316 9654 407344 12396
rect 408408 9716 408460 9722
rect 408408 9658 408460 9664
rect 406108 9648 406160 9654
rect 406108 9590 406160 9596
rect 407304 9648 407356 9654
rect 407304 9590 407356 9596
rect 408420 4078 408448 9658
rect 408512 7682 408540 22714
rect 409156 19990 409184 99350
rect 409800 43450 409828 102054
rect 410076 99414 410104 102068
rect 410904 102054 411010 102082
rect 410064 99408 410116 99414
rect 410064 99350 410116 99356
rect 410904 95266 410932 102054
rect 411352 100020 411404 100026
rect 411352 99962 411404 99968
rect 411168 99408 411220 99414
rect 411168 99350 411220 99356
rect 410892 95260 410944 95266
rect 410892 95202 410944 95208
rect 411076 95260 411128 95266
rect 411076 95202 411128 95208
rect 411088 87145 411116 95202
rect 411074 87136 411130 87145
rect 411074 87071 411130 87080
rect 410982 87000 411038 87009
rect 410982 86935 411038 86944
rect 410996 79914 411024 86935
rect 410904 79886 411024 79914
rect 410904 74526 410932 79886
rect 410892 74520 410944 74526
rect 410892 74462 410944 74468
rect 410984 70032 411036 70038
rect 410984 69974 411036 69980
rect 410996 63510 411024 69974
rect 410984 63504 411036 63510
rect 410984 63446 411036 63452
rect 411076 63504 411128 63510
rect 411076 63446 411128 63452
rect 411088 46866 411116 63446
rect 410996 46838 411116 46866
rect 410996 45558 411024 46838
rect 410984 45552 411036 45558
rect 410984 45494 411036 45500
rect 410984 45416 411036 45422
rect 410984 45358 411036 45364
rect 409880 44872 409932 44878
rect 409880 44814 409932 44820
rect 409788 43444 409840 43450
rect 409788 43386 409840 43392
rect 409144 19984 409196 19990
rect 409144 19926 409196 19932
rect 408592 13184 408644 13190
rect 408592 13126 408644 13132
rect 408500 7676 408552 7682
rect 408500 7618 408552 7624
rect 408604 7562 408632 13126
rect 409892 12442 409920 44814
rect 410996 21418 411024 45358
rect 410984 21412 411036 21418
rect 410984 21354 411036 21360
rect 409880 12436 409932 12442
rect 409880 12378 409932 12384
rect 410892 12436 410944 12442
rect 410892 12378 410944 12384
rect 409696 7676 409748 7682
rect 409696 7618 409748 7624
rect 408512 7534 408632 7562
rect 408408 4072 408460 4078
rect 408408 4014 408460 4020
rect 405648 4004 405700 4010
rect 405648 3946 405700 3952
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 407304 604 407356 610
rect 407304 546 407356 552
rect 406120 480 406148 546
rect 407316 480 407344 546
rect 408512 480 408540 7534
rect 409708 480 409736 7618
rect 410904 480 410932 12378
rect 411180 3942 411208 99350
rect 411364 12442 411392 99962
rect 411824 99414 411852 102068
rect 412652 99414 412680 102068
rect 413572 99482 413600 102068
rect 413560 99476 413612 99482
rect 413560 99418 413612 99424
rect 411812 99408 411864 99414
rect 411812 99350 411864 99356
rect 412548 99408 412600 99414
rect 412548 99350 412600 99356
rect 412640 99408 412692 99414
rect 412640 99350 412692 99356
rect 413928 99408 413980 99414
rect 413928 99350 413980 99356
rect 412560 46238 412588 99350
rect 412640 94512 412692 94518
rect 412640 94454 412692 94460
rect 412548 46232 412600 46238
rect 412548 46174 412600 46180
rect 412652 12442 412680 94454
rect 411352 12436 411404 12442
rect 411352 12378 411404 12384
rect 412088 12436 412140 12442
rect 412088 12378 412140 12384
rect 412640 12436 412692 12442
rect 412640 12378 412692 12384
rect 413284 12436 413336 12442
rect 413284 12378 413336 12384
rect 411168 3936 411220 3942
rect 411168 3878 411220 3884
rect 412100 480 412128 12378
rect 413296 480 413324 12378
rect 413940 3874 413968 99350
rect 414400 94518 414428 102068
rect 415044 102054 415242 102082
rect 416070 102054 416728 102082
rect 414388 94512 414440 94518
rect 414388 94454 414440 94460
rect 415044 92478 415072 102054
rect 416044 99476 416096 99482
rect 416044 99418 416096 99424
rect 415032 92472 415084 92478
rect 415032 92414 415084 92420
rect 415032 82884 415084 82890
rect 415032 82826 415084 82832
rect 415044 80102 415072 82826
rect 415032 80096 415084 80102
rect 415032 80038 415084 80044
rect 415124 79960 415176 79966
rect 415124 79902 415176 79908
rect 415136 73166 415164 79902
rect 415124 73160 415176 73166
rect 415124 73102 415176 73108
rect 415400 73160 415452 73166
rect 415400 73102 415452 73108
rect 415412 48958 415440 73102
rect 415400 48952 415452 48958
rect 415400 48894 415452 48900
rect 414020 47592 414072 47598
rect 414020 47534 414072 47540
rect 414032 12442 414060 47534
rect 415308 35964 415360 35970
rect 415308 35906 415360 35912
rect 415320 12594 415348 35906
rect 416056 22778 416084 99418
rect 416700 24138 416728 102054
rect 416976 99414 417004 102068
rect 417818 102054 418108 102082
rect 416964 99408 417016 99414
rect 416964 99350 417016 99356
rect 417976 99408 418028 99414
rect 417976 99350 418028 99356
rect 417988 49026 418016 99350
rect 416780 49020 416832 49026
rect 416780 48962 416832 48968
rect 417976 49020 418028 49026
rect 417976 48962 418028 48968
rect 416688 24132 416740 24138
rect 416688 24074 416740 24080
rect 416044 22772 416096 22778
rect 416044 22714 416096 22720
rect 415228 12566 415348 12594
rect 415228 12458 415256 12566
rect 414020 12436 414072 12442
rect 414020 12378 414072 12384
rect 414480 12436 414532 12442
rect 414480 12378 414532 12384
rect 415136 12430 415256 12458
rect 414492 9654 414520 12378
rect 414480 9648 414532 9654
rect 414480 9590 414532 9596
rect 413928 3868 413980 3874
rect 413928 3810 413980 3816
rect 415136 3806 415164 12430
rect 416792 7614 416820 48962
rect 416872 26920 416924 26926
rect 416872 26862 416924 26868
rect 415676 7608 415728 7614
rect 415676 7550 415728 7556
rect 416780 7608 416832 7614
rect 416780 7550 416832 7556
rect 415124 3800 415176 3806
rect 415124 3742 415176 3748
rect 414480 604 414532 610
rect 414480 546 414532 552
rect 414492 480 414520 546
rect 415688 480 415716 7550
rect 416884 480 416912 26862
rect 417976 7608 418028 7614
rect 417976 7550 418028 7556
rect 417988 480 418016 7550
rect 418080 3670 418108 102054
rect 418632 99822 418660 102068
rect 418620 99816 418672 99822
rect 418620 99758 418672 99764
rect 419460 50454 419488 102068
rect 420394 102054 420868 102082
rect 420184 99816 420236 99822
rect 420184 99758 420236 99764
rect 419448 50448 419500 50454
rect 419448 50390 419500 50396
rect 419540 28280 419592 28286
rect 419540 28222 419592 28228
rect 419552 12442 419580 28222
rect 420196 25566 420224 99758
rect 420184 25560 420236 25566
rect 420184 25502 420236 25508
rect 419540 12436 419592 12442
rect 419540 12378 419592 12384
rect 420368 12436 420420 12442
rect 420368 12378 420420 12384
rect 419172 6180 419224 6186
rect 419172 6122 419224 6128
rect 418068 3664 418120 3670
rect 418068 3606 418120 3612
rect 419184 480 419212 6122
rect 420380 480 420408 12378
rect 420840 3738 420868 102054
rect 421208 100706 421236 102068
rect 421944 102054 422050 102082
rect 422970 102054 423628 102082
rect 421196 100700 421248 100706
rect 421196 100642 421248 100648
rect 421944 96665 421972 102054
rect 422208 100700 422260 100706
rect 422208 100642 422260 100648
rect 421930 96656 421986 96665
rect 421930 96591 421986 96600
rect 422114 96656 422170 96665
rect 422114 96591 422170 96600
rect 422128 92478 422156 96591
rect 422116 92472 422168 92478
rect 422116 92414 422168 92420
rect 421932 82952 421984 82958
rect 421984 82900 422064 82906
rect 421932 82894 422064 82900
rect 421944 82878 422064 82894
rect 422036 81394 422064 82878
rect 422024 81388 422076 81394
rect 422024 81330 422076 81336
rect 422024 63572 422076 63578
rect 422024 63514 422076 63520
rect 422036 53854 422064 63514
rect 421932 53848 421984 53854
rect 421932 53790 421984 53796
rect 422024 53848 422076 53854
rect 422024 53790 422076 53796
rect 421944 51814 421972 53790
rect 421932 51808 421984 51814
rect 421932 51750 421984 51756
rect 420920 51740 420972 51746
rect 420920 51682 420972 51688
rect 420932 12442 420960 51682
rect 422220 26926 422248 100642
rect 422300 95940 422352 95946
rect 422300 95882 422352 95888
rect 422312 57934 422340 95882
rect 422300 57928 422352 57934
rect 422300 57870 422352 57876
rect 422392 57928 422444 57934
rect 422392 57870 422444 57876
rect 422404 48362 422432 57870
rect 422312 48334 422432 48362
rect 422312 38622 422340 48334
rect 422300 38616 422352 38622
rect 422300 38558 422352 38564
rect 422392 38616 422444 38622
rect 422392 38558 422444 38564
rect 422404 29050 422432 38558
rect 422312 29022 422432 29050
rect 422312 27606 422340 29022
rect 422300 27600 422352 27606
rect 422300 27542 422352 27548
rect 422208 26920 422260 26926
rect 422208 26862 422260 26868
rect 420920 12436 420972 12442
rect 420920 12378 420972 12384
rect 421564 12436 421616 12442
rect 421564 12378 421616 12384
rect 420828 3732 420880 3738
rect 420828 3674 420880 3680
rect 421576 480 421604 12378
rect 422760 9716 422812 9722
rect 422760 9658 422812 9664
rect 422772 480 422800 9658
rect 423600 3534 423628 102054
rect 423784 100638 423812 102068
rect 424626 102054 424916 102082
rect 423772 100632 423824 100638
rect 423772 100574 423824 100580
rect 424888 53174 424916 102054
rect 425440 100706 425468 102068
rect 426360 100706 426388 102068
rect 425428 100700 425480 100706
rect 425428 100642 425480 100648
rect 426256 100700 426308 100706
rect 426256 100642 426308 100648
rect 426348 100700 426400 100706
rect 426348 100642 426400 100648
rect 427084 100700 427136 100706
rect 427084 100642 427136 100648
rect 424968 100632 425020 100638
rect 424968 100574 425020 100580
rect 424876 53168 424928 53174
rect 424876 53110 424928 53116
rect 423680 29640 423732 29646
rect 423680 29582 423732 29588
rect 423588 3528 423640 3534
rect 423588 3470 423640 3476
rect 423692 626 423720 29582
rect 424980 28354 425008 100574
rect 426268 89706 426296 100642
rect 426084 89678 426296 89706
rect 426084 85542 426112 89678
rect 426072 85536 426124 85542
rect 426072 85478 426124 85484
rect 426164 85536 426216 85542
rect 426164 85478 426216 85484
rect 426176 70258 426204 85478
rect 426084 70230 426204 70258
rect 426084 60738 426112 70230
rect 426084 60710 426204 60738
rect 426176 60602 426204 60710
rect 426176 60574 426296 60602
rect 426268 57934 426296 60574
rect 426256 57928 426308 57934
rect 426256 57870 426308 57876
rect 426348 48340 426400 48346
rect 426348 48282 426400 48288
rect 426360 41426 426388 48282
rect 426176 41410 426388 41426
rect 426164 41404 426400 41410
rect 426216 41398 426348 41404
rect 426164 41346 426216 41352
rect 426348 41346 426400 41352
rect 424968 28348 425020 28354
rect 424968 28290 425020 28296
rect 426360 22250 426388 41346
rect 427096 31074 427124 100642
rect 427188 99482 427216 102068
rect 427176 99476 427228 99482
rect 427176 99418 427228 99424
rect 428016 98666 428044 102068
rect 428844 102054 428950 102082
rect 429778 102054 430528 102082
rect 428004 98660 428056 98666
rect 428004 98602 428056 98608
rect 428844 95266 428872 102054
rect 429108 98660 429160 98666
rect 429108 98602 429160 98608
rect 428832 95260 428884 95266
rect 428832 95202 428884 95208
rect 429016 95260 429068 95266
rect 429016 95202 429068 95208
rect 429028 95146 429056 95202
rect 428844 95118 429056 95146
rect 428844 85610 428872 95118
rect 428832 85604 428884 85610
rect 428832 85546 428884 85552
rect 428924 85604 428976 85610
rect 428924 85546 428976 85552
rect 428936 85513 428964 85546
rect 428646 85504 428702 85513
rect 428646 85439 428702 85448
rect 428922 85504 428978 85513
rect 428922 85439 428978 85448
rect 428660 80782 428688 85439
rect 428648 80776 428700 80782
rect 428648 80718 428700 80724
rect 428924 67652 428976 67658
rect 428924 67594 428976 67600
rect 428936 60738 428964 67594
rect 428936 60710 429056 60738
rect 429028 51882 429056 60710
rect 429016 51876 429068 51882
rect 429016 51818 429068 51824
rect 428832 48340 428884 48346
rect 428832 48282 428884 48288
rect 428844 41426 428872 48282
rect 428844 41398 429056 41426
rect 427820 32428 427872 32434
rect 427820 32370 427872 32376
rect 426440 31068 426492 31074
rect 426440 31010 426492 31016
rect 427084 31068 427136 31074
rect 427084 31010 427136 31016
rect 426084 22222 426388 22250
rect 426084 22114 426112 22222
rect 425992 22086 426112 22114
rect 425992 18170 426020 22086
rect 425992 18142 426112 18170
rect 425152 4820 425204 4826
rect 425152 4762 425204 4768
rect 423692 598 423996 626
rect 423968 480 423996 598
rect 425164 480 425192 4762
rect 426084 3602 426112 18142
rect 426452 12442 426480 31010
rect 427832 12442 427860 32370
rect 429028 31890 429056 41398
rect 429016 31884 429068 31890
rect 429016 31826 429068 31832
rect 429016 27736 429068 27742
rect 429016 27678 429068 27684
rect 429028 27606 429056 27678
rect 428740 27600 428792 27606
rect 428740 27542 428792 27548
rect 429016 27600 429068 27606
rect 429016 27542 429068 27548
rect 428752 14362 428780 27542
rect 428752 14334 428964 14362
rect 426440 12436 426492 12442
rect 426440 12378 426492 12384
rect 427544 12436 427596 12442
rect 427544 12378 427596 12384
rect 427820 12436 427872 12442
rect 427820 12378 427872 12384
rect 428740 12436 428792 12442
rect 428740 12378 428792 12384
rect 426348 8968 426400 8974
rect 426348 8910 426400 8916
rect 426072 3596 426124 3602
rect 426072 3538 426124 3544
rect 426360 480 426388 8910
rect 427556 480 427584 12378
rect 428752 480 428780 12378
rect 428936 9654 428964 14334
rect 428924 9648 428976 9654
rect 428924 9590 428976 9596
rect 429120 3466 429148 98602
rect 429200 54528 429252 54534
rect 429200 54470 429252 54476
rect 429212 12442 429240 54470
rect 430500 32434 430528 102054
rect 430592 100706 430620 102068
rect 430580 100700 430632 100706
rect 430580 100642 430632 100648
rect 431420 100026 431448 102068
rect 432340 100706 432368 102068
rect 433076 102054 433182 102082
rect 434010 102054 434668 102082
rect 431868 100700 431920 100706
rect 431868 100642 431920 100648
rect 432328 100700 432380 100706
rect 432328 100642 432380 100648
rect 431408 100020 431460 100026
rect 431408 99962 431460 99968
rect 431224 99476 431276 99482
rect 431224 99418 431276 99424
rect 431236 54534 431264 99418
rect 431880 55894 431908 100642
rect 433076 96665 433104 102054
rect 433984 100700 434036 100706
rect 433984 100642 434036 100648
rect 433062 96656 433118 96665
rect 433062 96591 433118 96600
rect 433246 96656 433302 96665
rect 433246 96591 433302 96600
rect 433260 89706 433288 96591
rect 433076 89678 433288 89706
rect 433076 80102 433104 89678
rect 433260 80102 433288 80133
rect 433064 80096 433116 80102
rect 433248 80096 433300 80102
rect 433116 80044 433248 80050
rect 433064 80038 433300 80044
rect 433076 80022 433288 80038
rect 433076 70394 433104 80022
rect 433076 70366 433288 70394
rect 433260 57254 433288 70366
rect 433248 57248 433300 57254
rect 433248 57190 433300 57196
rect 431960 56636 432012 56642
rect 431960 56578 432012 56584
rect 431868 55888 431920 55894
rect 431868 55830 431920 55836
rect 431224 54528 431276 54534
rect 431224 54470 431276 54476
rect 431972 46918 432000 56578
rect 433996 47598 434024 100642
rect 433984 47592 434036 47598
rect 433984 47534 434036 47540
rect 431960 46912 432012 46918
rect 431960 46854 432012 46860
rect 431960 37324 432012 37330
rect 431960 37266 432012 37272
rect 430580 33788 430632 33794
rect 430580 33730 430632 33736
rect 430488 32428 430540 32434
rect 430488 32370 430540 32376
rect 430592 12442 430620 33730
rect 431972 27606 432000 37266
rect 433340 35216 433392 35222
rect 433340 35158 433392 35164
rect 431960 27600 432012 27606
rect 431960 27542 432012 27548
rect 431960 18012 432012 18018
rect 431960 17954 432012 17960
rect 431972 14906 432000 17954
rect 431972 14878 432092 14906
rect 429200 12436 429252 12442
rect 429200 12378 429252 12384
rect 429936 12436 429988 12442
rect 429936 12378 429988 12384
rect 430580 12436 430632 12442
rect 430580 12378 430632 12384
rect 431132 12436 431184 12442
rect 431132 12378 431184 12384
rect 429108 3460 429160 3466
rect 429108 3402 429160 3408
rect 429948 480 429976 12378
rect 431144 9654 431172 12378
rect 432064 12322 432092 14878
rect 432064 12294 432368 12322
rect 432340 9654 432368 12294
rect 431132 9648 431184 9654
rect 431132 9590 431184 9596
rect 432328 9648 432380 9654
rect 432328 9590 432380 9596
rect 433352 6050 433380 35158
rect 433524 10328 433576 10334
rect 433524 10270 433576 10276
rect 433340 6044 433392 6050
rect 433340 5986 433392 5992
rect 431132 604 431184 610
rect 431132 546 431184 552
rect 432328 604 432380 610
rect 432328 546 432380 552
rect 431144 480 431172 546
rect 432340 480 432368 546
rect 433536 480 433564 10270
rect 434640 6186 434668 102054
rect 434916 100706 434944 102068
rect 435758 102054 435956 102082
rect 434904 100700 434956 100706
rect 434904 100642 434956 100648
rect 435928 58682 435956 102054
rect 436008 100700 436060 100706
rect 436008 100642 436060 100648
rect 434720 58676 434772 58682
rect 434720 58618 434772 58624
rect 435916 58676 435968 58682
rect 435916 58618 435968 58624
rect 434732 12442 434760 58618
rect 436020 33794 436048 100642
rect 436572 99414 436600 102068
rect 436560 99408 436612 99414
rect 436560 99350 436612 99356
rect 437400 35222 437428 102068
rect 438334 102054 438808 102082
rect 438124 99408 438176 99414
rect 438124 99350 438176 99356
rect 437480 89004 437532 89010
rect 437480 88946 437532 88952
rect 437388 35216 437440 35222
rect 437388 35158 437440 35164
rect 436008 33788 436060 33794
rect 436008 33730 436060 33736
rect 434720 12436 434772 12442
rect 434720 12378 434772 12384
rect 435824 12436 435876 12442
rect 435824 12378 435876 12384
rect 434628 6180 434680 6186
rect 434628 6122 434680 6128
rect 434628 6044 434680 6050
rect 434628 5986 434680 5992
rect 434640 480 434668 5986
rect 435836 480 435864 12378
rect 437020 11756 437072 11762
rect 437020 11698 437072 11704
rect 437032 480 437060 11698
rect 437492 3482 437520 88946
rect 438136 7614 438164 99350
rect 438780 83502 438808 102054
rect 439148 100706 439176 102068
rect 439884 102054 439990 102082
rect 440818 102054 441568 102082
rect 439136 100700 439188 100706
rect 439136 100642 439188 100648
rect 439884 96665 439912 102054
rect 440148 100700 440200 100706
rect 440148 100642 440200 100648
rect 439870 96656 439926 96665
rect 439870 96591 439926 96600
rect 440054 96656 440110 96665
rect 440054 96591 440110 96600
rect 440068 89706 440096 96591
rect 439884 89678 440096 89706
rect 438768 83496 438820 83502
rect 438768 83438 438820 83444
rect 439884 80102 439912 89678
rect 439872 80096 439924 80102
rect 439872 80038 439924 80044
rect 439964 79960 440016 79966
rect 439964 79902 440016 79908
rect 439976 77246 440004 79902
rect 439964 77240 440016 77246
rect 439964 77182 440016 77188
rect 440056 67652 440108 67658
rect 440056 67594 440108 67600
rect 440068 67538 440096 67594
rect 439976 67510 440096 67538
rect 439976 58002 440004 67510
rect 439872 57996 439924 58002
rect 439872 57938 439924 57944
rect 439964 57996 440016 58002
rect 439964 57938 440016 57944
rect 439884 57866 439912 57938
rect 439872 57860 439924 57866
rect 439872 57802 439924 57808
rect 439964 48340 440016 48346
rect 439964 48282 440016 48288
rect 439976 41478 440004 48282
rect 439964 41472 440016 41478
rect 439964 41414 440016 41420
rect 439872 38684 439924 38690
rect 439872 38626 439924 38632
rect 439884 36582 439912 38626
rect 438860 36576 438912 36582
rect 438860 36518 438912 36524
rect 439872 36576 439924 36582
rect 439872 36518 439924 36524
rect 438124 7608 438176 7614
rect 438124 7550 438176 7556
rect 438872 3482 438900 36518
rect 440160 8974 440188 100642
rect 441540 60042 441568 102054
rect 441724 98666 441752 102068
rect 442566 102054 442856 102082
rect 441712 98660 441764 98666
rect 441712 98602 441764 98608
rect 441620 90364 441672 90370
rect 441620 90306 441672 90312
rect 441528 60036 441580 60042
rect 441528 59978 441580 59984
rect 440240 14476 440292 14482
rect 440240 14418 440292 14424
rect 440148 8968 440200 8974
rect 440148 8910 440200 8916
rect 440252 3482 440280 14418
rect 441632 3482 441660 90306
rect 442828 37942 442856 102054
rect 443380 99482 443408 102068
rect 444300 100706 444328 102068
rect 445142 102054 445708 102082
rect 444288 100700 444340 100706
rect 444288 100642 444340 100648
rect 445024 100700 445076 100706
rect 445024 100642 445076 100648
rect 443368 99476 443420 99482
rect 443368 99418 443420 99424
rect 443000 98728 443052 98734
rect 443000 98670 443052 98676
rect 442816 37936 442868 37942
rect 442816 37878 442868 37884
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 98670
rect 444380 39364 444432 39370
rect 444380 39306 444432 39312
rect 443092 15904 443144 15910
rect 443092 15846 443144 15852
rect 443104 3482 443132 15846
rect 444392 3482 444420 39306
rect 445036 29646 445064 100642
rect 445680 39370 445708 102054
rect 445956 100706 445984 102068
rect 446798 102054 447088 102082
rect 445944 100700 445996 100706
rect 445944 100642 445996 100648
rect 446956 100700 447008 100706
rect 446956 100642 447008 100648
rect 446968 61402 446996 100642
rect 446956 61396 447008 61402
rect 446956 61338 447008 61344
rect 445668 39364 445720 39370
rect 445668 39306 445720 39312
rect 445024 29640 445076 29646
rect 445024 29582 445076 29588
rect 447060 10334 447088 102054
rect 447704 100162 447732 102068
rect 448532 100706 448560 102068
rect 449374 102054 449848 102082
rect 448520 100700 448572 100706
rect 448520 100642 448572 100648
rect 449716 100700 449768 100706
rect 449716 100642 449768 100648
rect 447692 100156 447744 100162
rect 447692 100098 447744 100104
rect 448428 100156 448480 100162
rect 448428 100098 448480 100104
rect 447784 99476 447836 99482
rect 447784 99418 447836 99424
rect 447796 17270 447824 99418
rect 448440 42090 448468 100098
rect 449728 72486 449756 100642
rect 449716 72480 449768 72486
rect 449716 72422 449768 72428
rect 448428 42084 448480 42090
rect 448428 42026 448480 42032
rect 447140 17264 447192 17270
rect 447140 17206 447192 17212
rect 447784 17264 447836 17270
rect 447784 17206 447836 17212
rect 447048 10328 447100 10334
rect 447048 10270 447100 10276
rect 446588 4140 446640 4146
rect 446588 4082 446640 4088
rect 443104 3454 444236 3482
rect 444392 3454 445432 3482
rect 444208 480 444236 3454
rect 445404 480 445432 3454
rect 446600 480 446628 4082
rect 447152 3482 447180 17206
rect 448520 13116 448572 13122
rect 448520 13058 448572 13064
rect 448532 3482 448560 13058
rect 449820 11762 449848 102054
rect 450280 99822 450308 102068
rect 451016 102054 451122 102082
rect 451950 102054 452608 102082
rect 450268 99816 450320 99822
rect 450268 99758 450320 99764
rect 451016 96665 451044 102054
rect 451924 99816 451976 99822
rect 451924 99758 451976 99764
rect 451002 96656 451058 96665
rect 451002 96591 451058 96600
rect 451186 96656 451242 96665
rect 451186 96591 451242 96600
rect 451200 89758 451228 96591
rect 451004 89752 451056 89758
rect 451004 89694 451056 89700
rect 451188 89752 451240 89758
rect 451188 89694 451240 89700
rect 451016 71058 451044 89694
rect 451004 71052 451056 71058
rect 451004 70994 451056 71000
rect 451936 44878 451964 99758
rect 451924 44872 451976 44878
rect 451924 44814 451976 44820
rect 451280 40724 451332 40730
rect 451280 40666 451332 40672
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 450176 4004 450228 4010
rect 450176 3946 450228 3952
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 3946
rect 451292 3398 451320 40666
rect 451372 18624 451424 18630
rect 451372 18566 451424 18572
rect 451280 3392 451332 3398
rect 451280 3334 451332 3340
rect 451384 1442 451412 18566
rect 452580 13122 452608 102054
rect 452764 100706 452792 102068
rect 453698 102054 453988 102082
rect 452752 100700 452804 100706
rect 452752 100642 452804 100648
rect 453856 100700 453908 100706
rect 453856 100642 453908 100648
rect 453868 82142 453896 100642
rect 453856 82136 453908 82142
rect 453856 82078 453908 82084
rect 453960 62830 453988 102054
rect 454512 97306 454540 102068
rect 454500 97300 454552 97306
rect 454500 97242 454552 97248
rect 455340 80714 455368 102068
rect 456182 102054 456748 102082
rect 455328 80708 455380 80714
rect 455328 80650 455380 80656
rect 456720 65550 456748 102054
rect 457088 95946 457116 102068
rect 457930 102054 458128 102082
rect 457076 95940 457128 95946
rect 457076 95882 457128 95888
rect 456708 65544 456760 65550
rect 456708 65486 456760 65492
rect 453948 62824 454000 62830
rect 453948 62766 454000 62772
rect 455420 43444 455472 43450
rect 455420 43386 455472 43392
rect 454040 19984 454092 19990
rect 454040 19926 454092 19932
rect 452568 13116 452620 13122
rect 452568 13058 452620 13064
rect 453672 4072 453724 4078
rect 453672 4014 453724 4020
rect 452476 3392 452528 3398
rect 452476 3334 452528 3340
rect 451292 1414 451412 1442
rect 451292 480 451320 1414
rect 452488 480 452516 3334
rect 453684 480 453712 4014
rect 454052 3482 454080 19926
rect 455432 3482 455460 43386
rect 458100 19990 458128 102054
rect 458744 99414 458772 102068
rect 459664 99414 459692 102068
rect 460506 102054 460796 102082
rect 458732 99408 458784 99414
rect 458732 99350 458784 99356
rect 459468 99408 459520 99414
rect 459468 99350 459520 99356
rect 459652 99408 459704 99414
rect 459652 99350 459704 99356
rect 459480 69698 459508 99350
rect 460768 79354 460796 102054
rect 461320 99414 461348 102068
rect 462148 99498 462176 102068
rect 463082 102054 463648 102082
rect 462148 99470 462452 99498
rect 460848 99408 460900 99414
rect 460848 99350 460900 99356
rect 461308 99408 461360 99414
rect 461308 99350 461360 99356
rect 462228 99408 462280 99414
rect 462228 99350 462280 99356
rect 460756 79348 460808 79354
rect 460756 79290 460808 79296
rect 459468 69692 459520 69698
rect 459468 69634 459520 69640
rect 459652 46232 459704 46238
rect 459652 46174 459704 46180
rect 458180 21412 458232 21418
rect 458180 21354 458232 21360
rect 458088 19984 458140 19990
rect 458088 19926 458140 19932
rect 457260 3936 457312 3942
rect 457260 3878 457312 3884
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3878
rect 458192 3482 458220 21354
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 46174
rect 460860 14482 460888 99350
rect 462240 66910 462268 99350
rect 462424 94518 462452 99470
rect 462320 94512 462372 94518
rect 462320 94454 462372 94460
rect 462412 94512 462464 94518
rect 462412 94454 462464 94460
rect 462228 66904 462280 66910
rect 462228 66846 462280 66852
rect 460940 22772 460992 22778
rect 460940 22714 460992 22720
rect 460848 14476 460900 14482
rect 460848 14418 460900 14424
rect 460848 3868 460900 3874
rect 460848 3810 460900 3816
rect 460860 480 460888 3810
rect 460952 3482 460980 22714
rect 462332 3482 462360 94454
rect 463620 21418 463648 102054
rect 463896 99414 463924 102068
rect 464738 102054 465028 102082
rect 465658 102054 466408 102082
rect 463884 99408 463936 99414
rect 463884 99350 463936 99356
rect 464896 99408 464948 99414
rect 464896 99350 464948 99356
rect 464908 68338 464936 99350
rect 464896 68332 464948 68338
rect 464896 68274 464948 68280
rect 463608 21412 463660 21418
rect 463608 21354 463660 21360
rect 465000 15910 465028 102054
rect 466380 43450 466408 102054
rect 466472 100706 466500 102068
rect 467314 102054 467696 102082
rect 466460 100700 466512 100706
rect 466460 100642 466512 100648
rect 467668 93158 467696 102054
rect 468128 100706 468156 102068
rect 467748 100700 467800 100706
rect 467748 100642 467800 100648
rect 468116 100700 468168 100706
rect 468116 100642 468168 100648
rect 467656 93152 467708 93158
rect 467656 93094 467708 93100
rect 467760 50386 467788 100642
rect 468772 96694 468800 102190
rect 469890 102054 470548 102082
rect 469864 100700 469916 100706
rect 469864 100642 469916 100648
rect 468760 96688 468812 96694
rect 468760 96630 468812 96636
rect 468852 96688 468904 96694
rect 468852 96630 468904 96636
rect 468864 96558 468892 96630
rect 468852 96552 468904 96558
rect 468852 96494 468904 96500
rect 469036 89684 469088 89690
rect 469036 89626 469088 89632
rect 469048 85542 469076 89626
rect 469036 85536 469088 85542
rect 469036 85478 469088 85484
rect 468944 67652 468996 67658
rect 468944 67594 468996 67600
rect 468956 60738 468984 67594
rect 468956 60710 469168 60738
rect 469140 51746 469168 60710
rect 469128 51740 469180 51746
rect 469128 51682 469180 51688
rect 469220 50448 469272 50454
rect 469220 50390 469272 50396
rect 467748 50380 467800 50386
rect 467748 50322 467800 50328
rect 466460 49020 466512 49026
rect 466460 48962 466512 48968
rect 466368 43444 466420 43450
rect 466368 43386 466420 43392
rect 465080 24132 465132 24138
rect 465080 24074 465132 24080
rect 464988 15904 465040 15910
rect 464988 15846 465040 15852
rect 464436 3800 464488 3806
rect 464436 3742 464488 3748
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3742
rect 465092 3482 465120 24074
rect 466472 3482 466500 48962
rect 467932 25560 467984 25566
rect 467932 25502 467984 25508
rect 467840 3664 467892 3670
rect 467840 3606 467892 3612
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 3210 467880 3606
rect 467944 3398 467972 25502
rect 469232 3482 469260 50390
rect 469876 22778 469904 100642
rect 470520 24138 470548 102054
rect 470704 100638 470732 102068
rect 471546 102054 471836 102082
rect 470692 100632 470744 100638
rect 470692 100574 470744 100580
rect 471808 53106 471836 102054
rect 471888 100632 471940 100638
rect 471888 100574 471940 100580
rect 471796 53100 471848 53106
rect 471796 53042 471848 53048
rect 471900 25566 471928 100574
rect 472452 100094 472480 102068
rect 472440 100088 472492 100094
rect 472440 100030 472492 100036
rect 473280 46238 473308 102068
rect 474122 102054 474688 102082
rect 473360 51808 473412 51814
rect 473360 51750 473412 51756
rect 473268 46232 473320 46238
rect 473268 46174 473320 46180
rect 471980 26920 472032 26926
rect 471980 26862 472032 26868
rect 471888 25560 471940 25566
rect 471888 25502 471940 25508
rect 470508 24132 470560 24138
rect 470508 24074 470560 24080
rect 469864 22772 469916 22778
rect 469864 22714 469916 22720
rect 471520 3732 471572 3738
rect 471520 3674 471572 3680
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 3182 467972 3210
rect 467944 480 467972 3182
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3674
rect 471992 3346 472020 26862
rect 473372 3346 473400 51750
rect 474660 4146 474688 102054
rect 475028 100706 475056 102068
rect 475870 102054 476068 102082
rect 476698 102054 477448 102082
rect 475016 100700 475068 100706
rect 475016 100642 475068 100648
rect 475936 100700 475988 100706
rect 475936 100642 475988 100648
rect 475948 91798 475976 100642
rect 475936 91792 475988 91798
rect 475936 91734 475988 91740
rect 476040 28286 476068 102054
rect 476120 28348 476172 28354
rect 476120 28290 476172 28296
rect 476028 28280 476080 28286
rect 476028 28222 476080 28228
rect 474648 4140 474700 4146
rect 474648 4082 474700 4088
rect 475108 3528 475160 3534
rect 475108 3470 475160 3476
rect 471992 3318 472756 3346
rect 473372 3318 473952 3346
rect 472728 480 472756 3318
rect 473924 480 473952 3318
rect 475120 480 475148 3470
rect 476132 3346 476160 28290
rect 477420 4078 477448 102054
rect 477512 99414 477540 102068
rect 478446 102054 478736 102082
rect 477500 99408 477552 99414
rect 477500 99350 477552 99356
rect 478708 77994 478736 102054
rect 479260 99414 479288 102068
rect 478788 99408 478840 99414
rect 478788 99350 478840 99356
rect 479248 99408 479300 99414
rect 479248 99350 479300 99356
rect 478696 77988 478748 77994
rect 478696 77930 478748 77936
rect 477592 53168 477644 53174
rect 477592 53110 477644 53116
rect 477408 4072 477460 4078
rect 477408 4014 477460 4020
rect 477604 3482 477632 53110
rect 478800 18630 478828 99350
rect 480088 90370 480116 102068
rect 481022 102054 481588 102082
rect 480168 99408 480220 99414
rect 480168 99350 480220 99356
rect 480076 90364 480128 90370
rect 480076 90306 480128 90312
rect 478880 31068 478932 31074
rect 478880 31010 478932 31016
rect 478788 18624 478840 18630
rect 478788 18566 478840 18572
rect 478696 3596 478748 3602
rect 478696 3538 478748 3544
rect 477512 3454 477632 3482
rect 476132 3318 476344 3346
rect 476316 480 476344 3318
rect 477512 480 477540 3454
rect 478708 480 478736 3538
rect 478892 3346 478920 31010
rect 480180 4010 480208 99350
rect 480260 54528 480312 54534
rect 480260 54470 480312 54476
rect 480168 4004 480220 4010
rect 480168 3946 480220 3952
rect 480272 3346 480300 54470
rect 481560 31074 481588 102054
rect 481836 99414 481864 102068
rect 482678 102054 482876 102082
rect 481824 99408 481876 99414
rect 481824 99350 481876 99356
rect 482848 89010 482876 102054
rect 483492 99414 483520 102068
rect 483664 100020 483716 100026
rect 483664 99962 483716 99968
rect 482928 99408 482980 99414
rect 482928 99350 482980 99356
rect 483480 99408 483532 99414
rect 483480 99350 483532 99356
rect 482836 89004 482888 89010
rect 482836 88946 482888 88952
rect 481548 31068 481600 31074
rect 481548 31010 481600 31016
rect 482940 3942 482968 99350
rect 483480 4820 483532 4826
rect 483480 4762 483532 4768
rect 482928 3936 482980 3942
rect 482928 3878 482980 3884
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 478892 3318 479932 3346
rect 480272 3318 481128 3346
rect 479904 480 479932 3318
rect 481100 480 481128 3318
rect 482296 480 482324 3402
rect 483492 480 483520 4762
rect 483676 4214 483704 99962
rect 484412 99414 484440 102068
rect 485240 100162 485268 102068
rect 485228 100156 485280 100162
rect 485228 100098 485280 100104
rect 486068 99414 486096 102068
rect 486910 102054 487108 102082
rect 487830 102054 488488 102082
rect 484308 99408 484360 99414
rect 484308 99350 484360 99356
rect 484400 99408 484452 99414
rect 484400 99350 484452 99356
rect 485688 99408 485740 99414
rect 485688 99350 485740 99356
rect 486056 99408 486108 99414
rect 486056 99350 486108 99356
rect 486976 99408 487028 99414
rect 486976 99350 487028 99356
rect 484320 49026 484348 99350
rect 484308 49020 484360 49026
rect 484308 48962 484360 48968
rect 484400 32428 484452 32434
rect 484400 32370 484452 32376
rect 483664 4208 483716 4214
rect 483664 4150 483716 4156
rect 484412 3346 484440 32370
rect 485700 3874 485728 99350
rect 486988 75206 487016 99350
rect 486976 75200 487028 75206
rect 486976 75142 487028 75148
rect 485780 55888 485832 55894
rect 485780 55830 485832 55836
rect 485688 3868 485740 3874
rect 485688 3810 485740 3816
rect 484412 3318 484624 3346
rect 484596 480 484624 3318
rect 485792 480 485820 55830
rect 486976 4208 487028 4214
rect 486976 4150 487028 4156
rect 486988 480 487016 4150
rect 487080 3806 487108 102054
rect 487160 47592 487212 47598
rect 487160 47534 487212 47540
rect 487068 3800 487120 3806
rect 487068 3742 487120 3748
rect 487172 3346 487200 47534
rect 488460 26926 488488 102054
rect 488644 99414 488672 102068
rect 489486 102054 489868 102082
rect 488632 99408 488684 99414
rect 488632 99350 488684 99356
rect 489736 99408 489788 99414
rect 489736 99350 489788 99356
rect 488540 57248 488592 57254
rect 488540 57190 488592 57196
rect 488448 26920 488500 26926
rect 488448 26862 488500 26868
rect 488552 3346 488580 57190
rect 489748 32434 489776 99350
rect 489736 32428 489788 32434
rect 489736 32370 489788 32376
rect 489840 3738 489868 102054
rect 490392 99414 490420 102068
rect 490380 99408 490432 99414
rect 490380 99350 490432 99356
rect 491220 73846 491248 102068
rect 492062 102054 492628 102082
rect 491944 99408 491996 99414
rect 491944 99350 491996 99356
rect 491956 86290 491984 99350
rect 491944 86284 491996 86290
rect 491944 86226 491996 86232
rect 491208 73840 491260 73846
rect 491208 73782 491260 73788
rect 491300 33788 491352 33794
rect 491300 33730 491352 33736
rect 490564 6180 490616 6186
rect 490564 6122 490616 6128
rect 489828 3732 489880 3738
rect 489828 3674 489880 3680
rect 487172 3318 488212 3346
rect 488552 3318 489408 3346
rect 488184 480 488212 3318
rect 489380 480 489408 3318
rect 490576 480 490604 6122
rect 491312 3482 491340 33730
rect 492600 3670 492628 102054
rect 492876 99414 492904 102068
rect 493810 102054 494008 102082
rect 492864 99408 492916 99414
rect 492864 99350 492916 99356
rect 493876 99408 493928 99414
rect 493876 99350 493928 99356
rect 493888 84862 493916 99350
rect 493876 84856 493928 84862
rect 493876 84798 493928 84804
rect 492680 58676 492732 58682
rect 492680 58618 492732 58624
rect 492588 3664 492640 3670
rect 492588 3606 492640 3612
rect 492692 3482 492720 58618
rect 493980 33794 494008 102054
rect 494624 99414 494652 102068
rect 495452 99414 495480 102068
rect 496386 102054 496768 102082
rect 494612 99408 494664 99414
rect 494612 99350 494664 99356
rect 495348 99408 495400 99414
rect 495348 99350 495400 99356
rect 495440 99408 495492 99414
rect 495440 99350 495492 99356
rect 496636 99408 496688 99414
rect 496636 99350 496688 99356
rect 494060 35216 494112 35222
rect 494060 35158 494112 35164
rect 493968 33788 494020 33794
rect 493968 33730 494020 33736
rect 494072 3534 494100 35158
rect 494152 7608 494204 7614
rect 494152 7550 494204 7556
rect 494060 3528 494112 3534
rect 491312 3454 491800 3482
rect 492692 3454 492996 3482
rect 494060 3470 494112 3476
rect 491772 480 491800 3454
rect 492968 480 492996 3454
rect 494164 480 494192 7550
rect 495360 5250 495388 99350
rect 496648 83502 496676 99350
rect 495440 83496 495492 83502
rect 495440 83438 495492 83444
rect 496636 83496 496688 83502
rect 496636 83438 496688 83444
rect 495176 5222 495388 5250
rect 495176 3602 495204 5222
rect 495164 3596 495216 3602
rect 495164 3538 495216 3544
rect 495348 3528 495400 3534
rect 495348 3470 495400 3476
rect 495452 3482 495480 83438
rect 496740 7614 496768 102054
rect 497200 99414 497228 102068
rect 498028 100026 498056 102068
rect 498870 102054 499528 102082
rect 498016 100020 498068 100026
rect 498016 99962 498068 99968
rect 497188 99408 497240 99414
rect 497188 99350 497240 99356
rect 498108 99408 498160 99414
rect 498108 99350 498160 99356
rect 497740 8968 497792 8974
rect 497740 8910 497792 8916
rect 496728 7608 496780 7614
rect 496728 7550 496780 7556
rect 495360 480 495388 3470
rect 495452 3454 496584 3482
rect 496556 480 496584 3454
rect 497752 480 497780 8910
rect 498120 3534 498148 99350
rect 498200 36576 498252 36582
rect 498200 36518 498252 36524
rect 498108 3528 498160 3534
rect 498108 3470 498160 3476
rect 498212 3482 498240 36518
rect 499500 8974 499528 102054
rect 499776 99414 499804 102068
rect 502984 100156 503036 100162
rect 502984 100098 503036 100104
rect 499764 99408 499816 99414
rect 499764 99350 499816 99356
rect 500868 99408 500920 99414
rect 500868 99350 500920 99356
rect 499580 60036 499632 60042
rect 499580 59978 499632 59984
rect 499488 8968 499540 8974
rect 499488 8910 499540 8916
rect 498212 3454 498976 3482
rect 498948 480 498976 3454
rect 499592 3346 499620 59978
rect 500880 3466 500908 99350
rect 500960 98660 501012 98666
rect 500960 98602 501012 98608
rect 500868 3460 500920 3466
rect 500868 3402 500920 3408
rect 499592 3318 500172 3346
rect 500144 480 500172 3318
rect 500972 626 501000 98602
rect 502340 37936 502392 37942
rect 502340 37878 502392 37884
rect 502352 3482 502380 37878
rect 502432 17264 502484 17270
rect 502432 17206 502484 17212
rect 502444 4214 502472 17206
rect 502996 6186 503024 100098
rect 504376 30326 504404 118079
rect 504468 41410 504496 128959
rect 504560 77246 504588 150719
rect 504652 88330 504680 161599
rect 504744 111790 504772 172479
rect 504836 124166 504864 183359
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 505006 139904 505062 139913
rect 505006 139839 505062 139848
rect 505020 139466 505048 139839
rect 505008 139460 505060 139466
rect 505008 139402 505060 139408
rect 519544 139460 519596 139466
rect 519544 139402 519596 139408
rect 504824 124160 504876 124166
rect 504824 124102 504876 124108
rect 504732 111784 504784 111790
rect 504732 111726 504784 111732
rect 505742 107400 505798 107409
rect 505742 107335 505798 107344
rect 504640 88324 504692 88330
rect 504640 88266 504692 88272
rect 504548 77240 504600 77246
rect 504548 77182 504600 77188
rect 504456 41404 504508 41410
rect 504456 41346 504508 41352
rect 505100 39364 505152 39370
rect 505100 39306 505152 39312
rect 504364 30320 504416 30326
rect 504364 30262 504416 30268
rect 503720 29640 503772 29646
rect 503720 29582 503772 29588
rect 502984 6180 503036 6186
rect 502984 6122 503036 6128
rect 502432 4208 502484 4214
rect 502432 4150 502484 4156
rect 503628 4208 503680 4214
rect 503628 4150 503680 4156
rect 502352 3454 502472 3482
rect 500972 598 501276 626
rect 501248 480 501276 598
rect 502444 480 502472 3454
rect 503640 480 503668 4150
rect 503732 3346 503760 29582
rect 505112 3346 505140 39306
rect 505756 17950 505784 107335
rect 507124 100088 507176 100094
rect 507124 100030 507176 100036
rect 506480 61396 506532 61402
rect 506480 61338 506532 61344
rect 505744 17944 505796 17950
rect 505744 17886 505796 17892
rect 506492 3346 506520 61338
rect 507136 4826 507164 100030
rect 518900 97300 518952 97306
rect 518900 97242 518952 97248
rect 516140 82136 516192 82142
rect 516140 82078 516192 82084
rect 510620 72480 510672 72486
rect 510620 72422 510672 72428
rect 509240 42084 509292 42090
rect 509240 42026 509292 42032
rect 507860 10328 507912 10334
rect 507860 10270 507912 10276
rect 507124 4820 507176 4826
rect 507124 4762 507176 4768
rect 507872 3346 507900 10270
rect 509252 3482 509280 42026
rect 510632 3482 510660 72422
rect 513380 71052 513432 71058
rect 513380 70994 513432 71000
rect 512000 44872 512052 44878
rect 512000 44814 512052 44820
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 506492 3318 507256 3346
rect 507872 3318 508452 3346
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507228 480 507256 3318
rect 508424 480 508452 3318
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 3398 512040 44814
rect 512092 11756 512144 11762
rect 512092 11698 512144 11704
rect 512000 3392 512052 3398
rect 512000 3334 512052 3340
rect 512104 1442 512132 11698
rect 513392 3482 513420 70994
rect 514760 13116 514812 13122
rect 514760 13058 514812 13064
rect 514772 3482 514800 13058
rect 516152 3482 516180 82078
rect 517520 62824 517572 62830
rect 517520 62766 517572 62772
rect 517532 3482 517560 62766
rect 518912 3482 518940 97242
rect 519556 64870 519584 139402
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 545764 100020 545816 100026
rect 545764 99962 545816 99968
rect 521660 95940 521712 95946
rect 521660 95882 521712 95888
rect 520280 80708 520332 80714
rect 520280 80650 520332 80656
rect 519544 64864 519596 64870
rect 519544 64806 519596 64812
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 512012 1414 512132 1442
rect 512012 480 512040 1414
rect 513208 480 513236 3334
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520292 480 520320 80650
rect 520372 65544 520424 65550
rect 520372 65486 520424 65492
rect 520384 3482 520412 65486
rect 521672 3482 521700 95882
rect 528560 94512 528612 94518
rect 528560 94454 528612 94460
rect 527180 79348 527232 79354
rect 527180 79290 527232 79296
rect 524420 69692 524472 69698
rect 524420 69634 524472 69640
rect 523040 19984 523092 19990
rect 523040 19926 523092 19932
rect 523052 3482 523080 19926
rect 524432 3482 524460 69634
rect 525800 14476 525852 14482
rect 525800 14418 525852 14424
rect 525812 3482 525840 14418
rect 527192 3482 527220 79290
rect 520384 3454 521516 3482
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 525812 3454 526300 3482
rect 527192 3454 527496 3482
rect 521488 480 521516 3454
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 3454
rect 527468 480 527496 3454
rect 528572 3398 528600 94454
rect 536840 93152 536892 93158
rect 536840 93094 536892 93100
rect 531320 68332 531372 68338
rect 531320 68274 531372 68280
rect 528652 66904 528704 66910
rect 528652 66846 528704 66852
rect 528560 3392 528612 3398
rect 528560 3334 528612 3340
rect 528664 480 528692 66846
rect 529940 21412 529992 21418
rect 529940 21354 529992 21360
rect 529952 3482 529980 21354
rect 531332 3482 531360 68274
rect 535460 50380 535512 50386
rect 535460 50322 535512 50328
rect 534080 43444 534132 43450
rect 534080 43386 534132 43392
rect 532700 15904 532752 15910
rect 532700 15846 532752 15852
rect 532712 3482 532740 15846
rect 534092 3482 534120 43386
rect 535472 3482 535500 50322
rect 536852 3482 536880 93094
rect 542360 53100 542412 53106
rect 542360 53042 542412 53048
rect 538220 51740 538272 51746
rect 538220 51682 538272 51688
rect 536932 22772 536984 22778
rect 536932 22714 536984 22720
rect 536944 4214 536972 22714
rect 536932 4208 536984 4214
rect 536932 4150 536984 4156
rect 538128 4208 538180 4214
rect 538128 4150 538180 4156
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 529848 3392 529900 3398
rect 529848 3334 529900 3340
rect 529860 480 529888 3334
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 4150
rect 538232 3346 538260 51682
rect 540980 25560 541032 25566
rect 540980 25502 541032 25508
rect 539600 24132 539652 24138
rect 539600 24074 539652 24080
rect 539612 3346 539640 24074
rect 540992 3346 541020 25502
rect 542372 3346 542400 53042
rect 545120 46232 545172 46238
rect 545120 46174 545172 46180
rect 544108 4820 544160 4826
rect 544108 4762 544160 4768
rect 538232 3318 539364 3346
rect 539612 3318 540560 3346
rect 540992 3318 541756 3346
rect 542372 3318 542952 3346
rect 539336 480 539364 3318
rect 540532 480 540560 3318
rect 541728 480 541756 3318
rect 542924 480 542952 3318
rect 544120 480 544148 4762
rect 545132 3346 545160 46174
rect 545776 4826 545804 99962
rect 546592 91792 546644 91798
rect 546592 91734 546644 91740
rect 545764 4820 545816 4826
rect 545764 4762 545816 4768
rect 546500 4140 546552 4146
rect 546500 4082 546552 4088
rect 545132 3318 545344 3346
rect 545316 480 545344 3318
rect 546512 480 546540 4082
rect 546604 3346 546632 91734
rect 554780 90364 554832 90370
rect 554780 90306 554832 90312
rect 552020 77988 552072 77994
rect 552020 77930 552072 77936
rect 547880 28280 547932 28286
rect 547880 28222 547932 28228
rect 547892 3482 547920 28222
rect 550640 18624 550692 18630
rect 550640 18566 550692 18572
rect 550088 4072 550140 4078
rect 550088 4014 550140 4020
rect 547892 3454 548932 3482
rect 546604 3318 547736 3346
rect 547708 480 547736 3318
rect 548904 480 548932 3454
rect 550100 480 550128 4014
rect 550652 3482 550680 18566
rect 552032 3482 552060 77930
rect 553584 4004 553636 4010
rect 553584 3946 553636 3952
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3946
rect 554792 480 554820 90306
rect 557540 89004 557592 89010
rect 557540 88946 557592 88952
rect 554872 31068 554924 31074
rect 554872 31010 554924 31016
rect 554884 3482 554912 31010
rect 557172 3936 557224 3942
rect 557172 3878 557224 3884
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3878
rect 557552 3482 557580 88946
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 568580 86284 568632 86290
rect 568580 86226 568632 86232
rect 563152 75200 563204 75206
rect 563152 75142 563204 75148
rect 558920 49020 558972 49026
rect 558920 48962 558972 48968
rect 558932 3482 558960 48962
rect 561956 6180 562008 6186
rect 561956 6122 562008 6128
rect 560760 3868 560812 3874
rect 560760 3810 560812 3816
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3810
rect 561968 480 561996 6122
rect 563164 480 563192 75142
rect 565820 32428 565872 32434
rect 565820 32370 565872 32376
rect 564440 26920 564492 26926
rect 564440 26862 564492 26868
rect 564348 3800 564400 3806
rect 564348 3742 564400 3748
rect 564360 480 564388 3742
rect 564452 3482 564480 26862
rect 565832 3482 565860 32370
rect 567844 3732 567896 3738
rect 567844 3674 567896 3680
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3674
rect 568592 3482 568620 86226
rect 571432 84856 571484 84862
rect 571432 84798 571484 84804
rect 569960 73840 570012 73846
rect 569960 73782 570012 73788
rect 569972 3482 570000 73782
rect 571340 3664 571392 3670
rect 571340 3606 571392 3612
rect 571352 3482 571380 3606
rect 571444 3602 571472 84798
rect 574744 83496 574796 83502
rect 574744 83438 574796 83444
rect 572720 33788 572772 33794
rect 572720 33730 572772 33736
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 572628 3596 572680 3602
rect 572628 3538 572680 3544
rect 568592 3454 569080 3482
rect 569972 3454 570276 3482
rect 571352 3454 571472 3482
rect 569052 480 569080 3454
rect 570248 480 570276 3454
rect 571444 480 571472 3454
rect 572640 480 572668 3538
rect 572732 3482 572760 33730
rect 572732 3454 573864 3482
rect 573836 480 573864 3454
rect 574756 3330 574784 83438
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 575020 3392 575072 3398
rect 575020 3334 575072 3340
rect 574744 3324 574796 3330
rect 574744 3266 574796 3272
rect 575032 480 575060 3334
rect 576216 3324 576268 3330
rect 576216 3266 576268 3272
rect 576228 480 576256 3266
rect 577424 480 577452 7550
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 579816 480 579844 4762
rect 581012 480 581040 8910
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667936 3478 667992
rect 3054 653520 3110 653576
rect 3238 624824 3294 624880
rect 3330 595992 3386 596048
rect 3514 610408 3570 610464
rect 3422 567296 3478 567352
rect 3422 553016 3478 553072
rect 3514 538600 3570 538656
rect 3422 509904 3478 509960
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 78678 595992 78734 596048
rect 504362 585520 504418 585576
rect 78678 584432 78734 584488
rect 78678 572736 78734 572792
rect 78678 561176 78734 561232
rect 78678 549480 78734 549536
rect 505006 574640 505062 574696
rect 504362 563760 504418 563816
rect 503810 552880 503866 552936
rect 505006 542000 505062 542056
rect 79322 537920 79378 537976
rect 504362 531120 504418 531176
rect 78678 526224 78734 526280
rect 504638 520240 504694 520296
rect 78678 514700 78680 514720
rect 78680 514700 78732 514720
rect 78732 514700 78734 514720
rect 78678 514664 78734 514700
rect 505006 509360 505062 509416
rect 78678 502968 78734 503024
rect 3514 495488 3570 495544
rect 3422 481072 3478 481128
rect 78678 491408 78734 491464
rect 78678 479712 78734 479768
rect 503718 476856 503774 476912
rect 78678 468152 78734 468208
rect 78678 456456 78734 456512
rect 505006 498480 505062 498536
rect 505006 487600 505062 487656
rect 505006 465976 505062 466032
rect 504362 455096 504418 455152
rect 3422 452376 3478 452432
rect 79322 444896 79378 444952
rect 505006 444216 505062 444272
rect 3146 437960 3202 438016
rect 79322 433200 79378 433256
rect 3238 423680 3294 423736
rect 503718 422456 503774 422512
rect 79414 421640 79470 421696
rect 79322 398384 79378 398440
rect 3146 394984 3202 395040
rect 3238 380568 3294 380624
rect 79506 409944 79562 410000
rect 79414 386688 79470 386744
rect 3146 366152 3202 366208
rect 79322 363432 79378 363488
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 78678 316920 78734 316976
rect 3330 308760 3386 308816
rect 3422 294344 3478 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3146 265648 3202 265704
rect 504638 433336 504694 433392
rect 580170 697992 580226 698048
rect 580262 686296 580318 686352
rect 542358 683168 542414 683224
rect 542726 683168 542782 683224
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 579894 592456 579950 592512
rect 580170 580760 580226 580816
rect 580354 639376 580410 639432
rect 580170 557232 580226 557288
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 579986 510312 580042 510368
rect 580262 498616 580318 498672
rect 579894 486784 579950 486840
rect 580170 463392 580226 463448
rect 580354 451696 580410 451752
rect 580170 439864 580226 439920
rect 580446 416472 580502 416528
rect 505006 411576 505062 411632
rect 580262 404776 580318 404832
rect 504362 400696 504418 400752
rect 579894 392944 579950 393000
rect 505006 389816 505062 389872
rect 503902 378936 503958 378992
rect 79690 375128 79746 375184
rect 79598 351872 79654 351928
rect 79506 340176 79562 340232
rect 79414 328616 79470 328672
rect 79322 305360 79378 305416
rect 78678 282104 78734 282160
rect 3238 251232 3294 251288
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 3422 208120 3478 208176
rect 3146 193840 3202 193896
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3422 78920 3478 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 4066 7112 4122 7168
rect 78678 247152 78734 247208
rect 580262 369552 580318 369608
rect 505006 368056 505062 368112
rect 580354 357856 580410 357912
rect 505006 357348 505008 357368
rect 505008 357348 505060 357368
rect 505060 357348 505062 357368
rect 505006 357312 505062 357348
rect 505006 346432 505062 346488
rect 580262 346024 580318 346080
rect 504546 335552 504602 335608
rect 505006 324672 505062 324728
rect 580170 322632 580226 322688
rect 504086 313792 504142 313848
rect 580170 310800 580226 310856
rect 504546 302912 504602 302968
rect 579802 299104 579858 299160
rect 79598 293664 79654 293720
rect 79506 270408 79562 270464
rect 79414 258848 79470 258904
rect 79322 235592 79378 235648
rect 78678 223896 78734 223952
rect 78678 212336 78734 212392
rect 78678 189100 78734 189136
rect 78678 189080 78680 189100
rect 78680 189080 78732 189100
rect 78732 189080 78734 189100
rect 78678 177384 78734 177440
rect 504362 292032 504418 292088
rect 504454 281152 504510 281208
rect 504362 270272 504418 270328
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 504546 259392 504602 259448
rect 504454 248512 504510 248568
rect 504362 237632 504418 237688
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 504638 226888 504694 226944
rect 504546 216008 504602 216064
rect 504454 205128 504510 205184
rect 79690 200640 79746 200696
rect 79598 165824 79654 165880
rect 79506 154128 79562 154184
rect 78678 142568 78734 142624
rect 79414 130872 79470 130928
rect 79322 119312 79378 119368
rect 31482 9696 31538 9752
rect 31666 9696 31722 9752
rect 504362 194248 504418 194304
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 504822 183368 504878 183424
rect 504730 172488 504786 172544
rect 504638 161608 504694 161664
rect 504546 150728 504602 150784
rect 504454 128968 504510 129024
rect 504362 118088 504418 118144
rect 88522 96600 88578 96656
rect 89166 96600 89222 96656
rect 101586 96600 101642 96656
rect 101954 96600 102010 96656
rect 104070 96600 104126 96656
rect 104530 96600 104586 96656
rect 105542 96600 105598 96656
rect 106186 96600 106242 96656
rect 106646 96600 106702 96656
rect 107106 96600 107162 96656
rect 108302 96600 108358 96656
rect 108762 96600 108818 96656
rect 111798 38664 111854 38720
rect 111798 38528 111854 38584
rect 124402 96600 124458 96656
rect 124954 96600 125010 96656
rect 142342 96600 142398 96656
rect 142894 96600 142950 96656
rect 153382 96600 153438 96656
rect 154026 96600 154082 96656
rect 164330 67496 164386 67552
rect 164422 67360 164478 67416
rect 175370 48184 175426 48240
rect 175462 48048 175518 48104
rect 200026 96600 200082 96656
rect 200302 96600 200358 96656
rect 206558 96600 206614 96656
rect 206926 96600 206982 96656
rect 207294 96600 207350 96656
rect 207018 77288 207074 77344
rect 207202 77288 207258 77344
rect 207754 96600 207810 96656
rect 208858 96620 208914 96656
rect 208858 96600 208860 96620
rect 208860 96600 208912 96620
rect 208912 96600 208914 96620
rect 209502 96600 209558 96656
rect 213090 96600 213146 96656
rect 213734 96600 213790 96656
rect 226522 86944 226578 87000
rect 226982 86944 227038 87000
rect 229006 75792 229062 75848
rect 229006 66272 229062 66328
rect 229282 75792 229338 75848
rect 229282 66272 229338 66328
rect 230662 67632 230718 67688
rect 230846 67632 230902 67688
rect 248694 48184 248750 48240
rect 248970 48184 249026 48240
rect 255870 87080 255926 87136
rect 255410 86944 255466 87000
rect 261206 77288 261262 77344
rect 260838 77152 260894 77208
rect 272062 38664 272118 38720
rect 272246 38664 272302 38720
rect 271786 29008 271842 29064
rect 271970 29008 272026 29064
rect 310150 96600 310206 96656
rect 310334 96600 310390 96656
rect 321190 66272 321246 66328
rect 321374 66272 321430 66328
rect 321190 46824 321246 46880
rect 321190 37304 321246 37360
rect 328090 96600 328146 96656
rect 328274 96620 328330 96656
rect 328274 96600 328276 96620
rect 328276 96600 328328 96620
rect 328328 96600 328330 96620
rect 327998 86944 328054 87000
rect 328182 86944 328238 87000
rect 332322 96600 332378 96656
rect 332506 96600 332562 96656
rect 332414 67632 332470 67688
rect 332598 67632 332654 67688
rect 350262 86944 350318 87000
rect 350446 86944 350502 87000
rect 350354 54032 350410 54088
rect 350354 53896 350410 53952
rect 350354 53760 350410 53816
rect 350538 53760 350594 53816
rect 379242 96600 379298 96656
rect 379426 96600 379482 96656
rect 390190 77288 390246 77344
rect 390374 77288 390430 77344
rect 411074 87080 411130 87136
rect 410982 86944 411038 87000
rect 421930 96600 421986 96656
rect 422114 96600 422170 96656
rect 428646 85448 428702 85504
rect 428922 85448 428978 85504
rect 433062 96600 433118 96656
rect 433246 96600 433302 96656
rect 439870 96600 439926 96656
rect 440054 96600 440110 96656
rect 451002 96600 451058 96656
rect 451186 96600 451242 96656
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 505006 139848 505062 139904
rect 505742 107344 505798 107400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 542353 683226 542419 683229
rect 542721 683226 542787 683229
rect 542353 683224 542787 683226
rect 542353 683168 542358 683224
rect 542414 683168 542726 683224
rect 542782 683168 542787 683224
rect 542353 683166 542787 683168
rect 542353 683163 542419 683166
rect 542721 683163 542787 683166
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3233 624882 3299 624885
rect -960 624880 3299 624882
rect -960 624824 3238 624880
rect 3294 624824 3299 624880
rect -960 624822 3299 624824
rect -960 624732 480 624822
rect 3233 624819 3299 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3509 610466 3575 610469
rect -960 610464 3575 610466
rect -960 610408 3514 610464
rect 3570 610408 3575 610464
rect -960 610406 3575 610408
rect -960 610316 480 610406
rect 3509 610403 3575 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 78673 596050 78739 596053
rect 78673 596048 82156 596050
rect 78673 595992 78678 596048
rect 78734 595992 82156 596048
rect 78673 595990 82156 595992
rect 78673 595987 78739 595990
rect 579889 592514 579955 592517
rect 583520 592514 584960 592604
rect 579889 592512 584960 592514
rect 579889 592456 579894 592512
rect 579950 592456 584960 592512
rect 579889 592454 584960 592456
rect 579889 592451 579955 592454
rect 583520 592364 584960 592454
rect 504357 585578 504423 585581
rect 501860 585576 504423 585578
rect 501860 585520 504362 585576
rect 504418 585520 504423 585576
rect 501860 585518 504423 585520
rect 504357 585515 504423 585518
rect 78673 584490 78739 584493
rect 78673 584488 82156 584490
rect 78673 584432 78678 584488
rect 78734 584432 82156 584488
rect 78673 584430 82156 584432
rect 78673 584427 78739 584430
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 505001 574698 505067 574701
rect 501860 574696 505067 574698
rect 501860 574640 505006 574696
rect 505062 574640 505067 574696
rect 501860 574638 505067 574640
rect 505001 574635 505067 574638
rect 78673 572794 78739 572797
rect 78673 572792 82156 572794
rect 78673 572736 78678 572792
rect 78734 572736 82156 572792
rect 78673 572734 82156 572736
rect 78673 572731 78739 572734
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 504357 563818 504423 563821
rect 501860 563816 504423 563818
rect 501860 563760 504362 563816
rect 504418 563760 504423 563816
rect 501860 563758 504423 563760
rect 504357 563755 504423 563758
rect 78673 561234 78739 561237
rect 78673 561232 82156 561234
rect 78673 561176 78678 561232
rect 78734 561176 82156 561232
rect 78673 561174 82156 561176
rect 78673 561171 78739 561174
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 503805 552938 503871 552941
rect 501860 552936 503871 552938
rect 501860 552880 503810 552936
rect 503866 552880 503871 552936
rect 501860 552878 503871 552880
rect 503805 552875 503871 552878
rect 78673 549538 78739 549541
rect 78673 549536 82156 549538
rect 78673 549480 78678 549536
rect 78734 549480 82156 549536
rect 78673 549478 82156 549480
rect 78673 549475 78739 549478
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 505001 542058 505067 542061
rect 501860 542056 505067 542058
rect 501860 542000 505006 542056
rect 505062 542000 505067 542056
rect 501860 541998 505067 542000
rect 505001 541995 505067 541998
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 79317 537978 79383 537981
rect 79317 537976 82156 537978
rect 79317 537920 79322 537976
rect 79378 537920 82156 537976
rect 79317 537918 82156 537920
rect 79317 537915 79383 537918
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 504357 531178 504423 531181
rect 501860 531176 504423 531178
rect 501860 531120 504362 531176
rect 504418 531120 504423 531176
rect 501860 531118 504423 531120
rect 504357 531115 504423 531118
rect 78673 526282 78739 526285
rect 78673 526280 82156 526282
rect 78673 526224 78678 526280
rect 78734 526224 82156 526280
rect 78673 526222 82156 526224
rect 78673 526219 78739 526222
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 504633 520298 504699 520301
rect 501860 520296 504699 520298
rect 501860 520240 504638 520296
rect 504694 520240 504699 520296
rect 501860 520238 504699 520240
rect 504633 520235 504699 520238
rect 78673 514722 78739 514725
rect 78673 514720 82156 514722
rect 78673 514664 78678 514720
rect 78734 514664 82156 514720
rect 78673 514662 82156 514664
rect 78673 514659 78739 514662
rect 579981 510370 580047 510373
rect 583520 510370 584960 510460
rect 579981 510368 584960 510370
rect 579981 510312 579986 510368
rect 580042 510312 584960 510368
rect 579981 510310 584960 510312
rect 579981 510307 580047 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 505001 509418 505067 509421
rect 501860 509416 505067 509418
rect 501860 509360 505006 509416
rect 505062 509360 505067 509416
rect 501860 509358 505067 509360
rect 505001 509355 505067 509358
rect 78673 503026 78739 503029
rect 78673 503024 82156 503026
rect 78673 502968 78678 503024
rect 78734 502968 82156 503024
rect 78673 502966 82156 502968
rect 78673 502963 78739 502966
rect 580257 498674 580323 498677
rect 583520 498674 584960 498764
rect 580257 498672 584960 498674
rect 580257 498616 580262 498672
rect 580318 498616 584960 498672
rect 580257 498614 584960 498616
rect 580257 498611 580323 498614
rect 505001 498538 505067 498541
rect 501860 498536 505067 498538
rect 501860 498480 505006 498536
rect 505062 498480 505067 498536
rect 583520 498524 584960 498614
rect 501860 498478 505067 498480
rect 505001 498475 505067 498478
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 78673 491466 78739 491469
rect 78673 491464 82156 491466
rect 78673 491408 78678 491464
rect 78734 491408 82156 491464
rect 78673 491406 82156 491408
rect 78673 491403 78739 491406
rect 505001 487658 505067 487661
rect 501860 487656 505067 487658
rect 501860 487600 505006 487656
rect 505062 487600 505067 487656
rect 501860 487598 505067 487600
rect 505001 487595 505067 487598
rect 579889 486842 579955 486845
rect 583520 486842 584960 486932
rect 579889 486840 584960 486842
rect 579889 486784 579894 486840
rect 579950 486784 584960 486840
rect 579889 486782 584960 486784
rect 579889 486779 579955 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3417 481130 3483 481133
rect -960 481128 3483 481130
rect -960 481072 3422 481128
rect 3478 481072 3483 481128
rect -960 481070 3483 481072
rect -960 480980 480 481070
rect 3417 481067 3483 481070
rect 78673 479770 78739 479773
rect 78673 479768 82156 479770
rect 78673 479712 78678 479768
rect 78734 479712 82156 479768
rect 78673 479710 82156 479712
rect 78673 479707 78739 479710
rect 503713 476914 503779 476917
rect 501860 476912 503779 476914
rect 501860 476856 503718 476912
rect 503774 476856 503779 476912
rect 501860 476854 503779 476856
rect 503713 476851 503779 476854
rect 583520 474996 584960 475236
rect 78673 468210 78739 468213
rect 78673 468208 82156 468210
rect 78673 468152 78678 468208
rect 78734 468152 82156 468208
rect 78673 468150 82156 468152
rect 78673 468147 78739 468150
rect -960 466700 480 466940
rect 505001 466034 505067 466037
rect 501860 466032 505067 466034
rect 501860 465976 505006 466032
rect 505062 465976 505067 466032
rect 501860 465974 505067 465976
rect 505001 465971 505067 465974
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 78673 456514 78739 456517
rect 78673 456512 82156 456514
rect 78673 456456 78678 456512
rect 78734 456456 82156 456512
rect 78673 456454 82156 456456
rect 78673 456451 78739 456454
rect 504357 455154 504423 455157
rect 501860 455152 504423 455154
rect 501860 455096 504362 455152
rect 504418 455096 504423 455152
rect 501860 455094 504423 455096
rect 504357 455091 504423 455094
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580349 451754 580415 451757
rect 583520 451754 584960 451844
rect 580349 451752 584960 451754
rect 580349 451696 580354 451752
rect 580410 451696 584960 451752
rect 580349 451694 584960 451696
rect 580349 451691 580415 451694
rect 583520 451604 584960 451694
rect 79317 444954 79383 444957
rect 79317 444952 82156 444954
rect 79317 444896 79322 444952
rect 79378 444896 82156 444952
rect 79317 444894 82156 444896
rect 79317 444891 79383 444894
rect 505001 444274 505067 444277
rect 501860 444272 505067 444274
rect 501860 444216 505006 444272
rect 505062 444216 505067 444272
rect 501860 444214 505067 444216
rect 505001 444211 505067 444214
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 504633 433394 504699 433397
rect 501860 433392 504699 433394
rect 501860 433336 504638 433392
rect 504694 433336 504699 433392
rect 501860 433334 504699 433336
rect 504633 433331 504699 433334
rect 79317 433258 79383 433261
rect 79317 433256 82156 433258
rect 79317 433200 79322 433256
rect 79378 433200 82156 433256
rect 79317 433198 82156 433200
rect 79317 433195 79383 433198
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 503713 422514 503779 422517
rect 501860 422512 503779 422514
rect 501860 422456 503718 422512
rect 503774 422456 503779 422512
rect 501860 422454 503779 422456
rect 503713 422451 503779 422454
rect 79409 421698 79475 421701
rect 79409 421696 82156 421698
rect 79409 421640 79414 421696
rect 79470 421640 82156 421696
rect 79409 421638 82156 421640
rect 79409 421635 79475 421638
rect 580441 416530 580507 416533
rect 583520 416530 584960 416620
rect 580441 416528 584960 416530
rect 580441 416472 580446 416528
rect 580502 416472 584960 416528
rect 580441 416470 584960 416472
rect 580441 416467 580507 416470
rect 583520 416380 584960 416470
rect 505001 411634 505067 411637
rect 501860 411632 505067 411634
rect 501860 411576 505006 411632
rect 505062 411576 505067 411632
rect 501860 411574 505067 411576
rect 505001 411571 505067 411574
rect 79501 410002 79567 410005
rect 79501 410000 82156 410002
rect 79501 409944 79506 410000
rect 79562 409944 82156 410000
rect 79501 409942 82156 409944
rect 79501 409939 79567 409942
rect -960 409172 480 409412
rect 580257 404834 580323 404837
rect 583520 404834 584960 404924
rect 580257 404832 584960 404834
rect 580257 404776 580262 404832
rect 580318 404776 584960 404832
rect 580257 404774 584960 404776
rect 580257 404771 580323 404774
rect 583520 404684 584960 404774
rect 504357 400754 504423 400757
rect 501860 400752 504423 400754
rect 501860 400696 504362 400752
rect 504418 400696 504423 400752
rect 501860 400694 504423 400696
rect 504357 400691 504423 400694
rect 79317 398442 79383 398445
rect 79317 398440 82156 398442
rect 79317 398384 79322 398440
rect 79378 398384 82156 398440
rect 79317 398382 82156 398384
rect 79317 398379 79383 398382
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 579889 393002 579955 393005
rect 583520 393002 584960 393092
rect 579889 393000 584960 393002
rect 579889 392944 579894 393000
rect 579950 392944 584960 393000
rect 579889 392942 584960 392944
rect 579889 392939 579955 392942
rect 583520 392852 584960 392942
rect 505001 389874 505067 389877
rect 501860 389872 505067 389874
rect 501860 389816 505006 389872
rect 505062 389816 505067 389872
rect 501860 389814 505067 389816
rect 505001 389811 505067 389814
rect 79409 386746 79475 386749
rect 79409 386744 82156 386746
rect 79409 386688 79414 386744
rect 79470 386688 82156 386744
rect 79409 386686 82156 386688
rect 79409 386683 79475 386686
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 503897 378994 503963 378997
rect 501860 378992 503963 378994
rect 501860 378936 503902 378992
rect 503958 378936 503963 378992
rect 501860 378934 503963 378936
rect 503897 378931 503963 378934
rect 79685 375186 79751 375189
rect 79685 375184 82156 375186
rect 79685 375128 79690 375184
rect 79746 375128 82156 375184
rect 79685 375126 82156 375128
rect 79685 375123 79751 375126
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 583520 369460 584960 369550
rect 505001 368114 505067 368117
rect 501860 368112 505067 368114
rect 501860 368056 505006 368112
rect 505062 368056 505067 368112
rect 501860 368054 505067 368056
rect 505001 368051 505067 368054
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 79317 363490 79383 363493
rect 79317 363488 82156 363490
rect 79317 363432 79322 363488
rect 79378 363432 82156 363488
rect 79317 363430 82156 363432
rect 79317 363427 79383 363430
rect 580349 357914 580415 357917
rect 583520 357914 584960 358004
rect 580349 357912 584960 357914
rect 580349 357856 580354 357912
rect 580410 357856 584960 357912
rect 580349 357854 584960 357856
rect 580349 357851 580415 357854
rect 583520 357764 584960 357854
rect 505001 357370 505067 357373
rect 501860 357368 505067 357370
rect 501860 357312 505006 357368
rect 505062 357312 505067 357368
rect 501860 357310 505067 357312
rect 505001 357307 505067 357310
rect -960 351780 480 352020
rect 79593 351930 79659 351933
rect 79593 351928 82156 351930
rect 79593 351872 79598 351928
rect 79654 351872 82156 351928
rect 79593 351870 82156 351872
rect 79593 351867 79659 351870
rect 505001 346490 505067 346493
rect 501860 346488 505067 346490
rect 501860 346432 505006 346488
rect 505062 346432 505067 346488
rect 501860 346430 505067 346432
rect 505001 346427 505067 346430
rect 580257 346082 580323 346085
rect 583520 346082 584960 346172
rect 580257 346080 584960 346082
rect 580257 346024 580262 346080
rect 580318 346024 584960 346080
rect 580257 346022 584960 346024
rect 580257 346019 580323 346022
rect 583520 345932 584960 346022
rect 79501 340234 79567 340237
rect 79501 340232 82156 340234
rect 79501 340176 79506 340232
rect 79562 340176 82156 340232
rect 79501 340174 82156 340176
rect 79501 340171 79567 340174
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 504541 335610 504607 335613
rect 501860 335608 504607 335610
rect 501860 335552 504546 335608
rect 504602 335552 504607 335608
rect 501860 335550 504607 335552
rect 504541 335547 504607 335550
rect 583520 334236 584960 334476
rect 79409 328674 79475 328677
rect 79409 328672 82156 328674
rect 79409 328616 79414 328672
rect 79470 328616 82156 328672
rect 79409 328614 82156 328616
rect 79409 328611 79475 328614
rect 505001 324730 505067 324733
rect 501860 324728 505067 324730
rect 501860 324672 505006 324728
rect 505062 324672 505067 324728
rect 501860 324670 505067 324672
rect 505001 324667 505067 324670
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 78673 316978 78739 316981
rect 78673 316976 82156 316978
rect 78673 316920 78678 316976
rect 78734 316920 82156 316976
rect 78673 316918 82156 316920
rect 78673 316915 78739 316918
rect 504081 313850 504147 313853
rect 501860 313848 504147 313850
rect 501860 313792 504086 313848
rect 504142 313792 504147 313848
rect 501860 313790 504147 313792
rect 504081 313787 504147 313790
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 79317 305418 79383 305421
rect 79317 305416 82156 305418
rect 79317 305360 79322 305416
rect 79378 305360 82156 305416
rect 79317 305358 82156 305360
rect 79317 305355 79383 305358
rect 504541 302970 504607 302973
rect 501860 302968 504607 302970
rect 501860 302912 504546 302968
rect 504602 302912 504607 302968
rect 501860 302910 504607 302912
rect 504541 302907 504607 302910
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 79593 293722 79659 293725
rect 79593 293720 82156 293722
rect 79593 293664 79598 293720
rect 79654 293664 82156 293720
rect 79593 293662 82156 293664
rect 79593 293659 79659 293662
rect 504357 292090 504423 292093
rect 501860 292088 504423 292090
rect 501860 292032 504362 292088
rect 504418 292032 504423 292088
rect 501860 292030 504423 292032
rect 504357 292027 504423 292030
rect 583520 287316 584960 287556
rect 78673 282162 78739 282165
rect 78673 282160 82156 282162
rect 78673 282104 78678 282160
rect 78734 282104 82156 282160
rect 78673 282102 82156 282104
rect 78673 282099 78739 282102
rect 504449 281210 504515 281213
rect 501860 281208 504515 281210
rect 501860 281152 504454 281208
rect 504510 281152 504515 281208
rect 501860 281150 504515 281152
rect 504449 281147 504515 281150
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 79501 270466 79567 270469
rect 79501 270464 82156 270466
rect 79501 270408 79506 270464
rect 79562 270408 82156 270464
rect 79501 270406 82156 270408
rect 79501 270403 79567 270406
rect 504357 270330 504423 270333
rect 501860 270328 504423 270330
rect 501860 270272 504362 270328
rect 504418 270272 504423 270328
rect 501860 270270 504423 270272
rect 504357 270267 504423 270270
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 504541 259450 504607 259453
rect 501860 259448 504607 259450
rect 501860 259392 504546 259448
rect 504602 259392 504607 259448
rect 501860 259390 504607 259392
rect 504541 259387 504607 259390
rect 79409 258906 79475 258909
rect 79409 258904 82156 258906
rect 79409 258848 79414 258904
rect 79470 258848 82156 258904
rect 79409 258846 82156 258848
rect 79409 258843 79475 258846
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3233 251290 3299 251293
rect -960 251288 3299 251290
rect -960 251232 3238 251288
rect 3294 251232 3299 251288
rect -960 251230 3299 251232
rect -960 251140 480 251230
rect 3233 251227 3299 251230
rect 504449 248570 504515 248573
rect 501860 248568 504515 248570
rect 501860 248512 504454 248568
rect 504510 248512 504515 248568
rect 501860 248510 504515 248512
rect 504449 248507 504515 248510
rect 78673 247210 78739 247213
rect 78673 247208 82156 247210
rect 78673 247152 78678 247208
rect 78734 247152 82156 247208
rect 78673 247150 82156 247152
rect 78673 247147 78739 247150
rect 583520 240396 584960 240636
rect 504357 237690 504423 237693
rect 501860 237688 504423 237690
rect 501860 237632 504362 237688
rect 504418 237632 504423 237688
rect 501860 237630 504423 237632
rect 504357 237627 504423 237630
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 79317 235650 79383 235653
rect 79317 235648 82156 235650
rect 79317 235592 79322 235648
rect 79378 235592 82156 235648
rect 79317 235590 82156 235592
rect 79317 235587 79383 235590
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 504633 226946 504699 226949
rect 501860 226944 504699 226946
rect 501860 226888 504638 226944
rect 504694 226888 504699 226944
rect 501860 226886 504699 226888
rect 504633 226883 504699 226886
rect 78673 223954 78739 223957
rect 78673 223952 82156 223954
rect 78673 223896 78678 223952
rect 78734 223896 82156 223952
rect 78673 223894 82156 223896
rect 78673 223891 78739 223894
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 504541 216066 504607 216069
rect 501860 216064 504607 216066
rect 501860 216008 504546 216064
rect 504602 216008 504607 216064
rect 501860 216006 504607 216008
rect 504541 216003 504607 216006
rect 78673 212394 78739 212397
rect 78673 212392 82156 212394
rect 78673 212336 78678 212392
rect 78734 212336 82156 212392
rect 78673 212334 82156 212336
rect 78673 212331 78739 212334
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 504449 205186 504515 205189
rect 501860 205184 504515 205186
rect 501860 205128 504454 205184
rect 504510 205128 504515 205184
rect 583520 205172 584960 205262
rect 501860 205126 504515 205128
rect 504449 205123 504515 205126
rect 79685 200698 79751 200701
rect 79685 200696 82156 200698
rect 79685 200640 79690 200696
rect 79746 200640 82156 200696
rect 79685 200638 82156 200640
rect 79685 200635 79751 200638
rect 504357 194306 504423 194309
rect 501860 194304 504423 194306
rect 501860 194248 504362 194304
rect 504418 194248 504423 194304
rect 501860 194246 504423 194248
rect 504357 194243 504423 194246
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 78673 189138 78739 189141
rect 78673 189136 82156 189138
rect 78673 189080 78678 189136
rect 78734 189080 82156 189136
rect 78673 189078 82156 189080
rect 78673 189075 78739 189078
rect 504817 183426 504883 183429
rect 501860 183424 504883 183426
rect 501860 183368 504822 183424
rect 504878 183368 504883 183424
rect 501860 183366 504883 183368
rect 504817 183363 504883 183366
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 78673 177442 78739 177445
rect 78673 177440 82156 177442
rect 78673 177384 78678 177440
rect 78734 177384 82156 177440
rect 78673 177382 82156 177384
rect 78673 177379 78739 177382
rect 504725 172546 504791 172549
rect 501860 172544 504791 172546
rect 501860 172488 504730 172544
rect 504786 172488 504791 172544
rect 501860 172486 504791 172488
rect 504725 172483 504791 172486
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 79593 165882 79659 165885
rect 79593 165880 82156 165882
rect 79593 165824 79598 165880
rect 79654 165824 82156 165880
rect 79593 165822 82156 165824
rect 79593 165819 79659 165822
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 504633 161666 504699 161669
rect 501860 161664 504699 161666
rect 501860 161608 504638 161664
rect 504694 161608 504699 161664
rect 501860 161606 504699 161608
rect 504633 161603 504699 161606
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 79501 154186 79567 154189
rect 79501 154184 82156 154186
rect 79501 154128 79506 154184
rect 79562 154128 82156 154184
rect 79501 154126 82156 154128
rect 79501 154123 79567 154126
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect 504541 150786 504607 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect 501860 150784 504607 150786
rect 501860 150728 504546 150784
rect 504602 150728 504607 150784
rect 501860 150726 504607 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 504541 150723 504607 150726
rect 583520 146556 584960 146796
rect 78673 142626 78739 142629
rect 78673 142624 82156 142626
rect 78673 142568 78678 142624
rect 78734 142568 82156 142624
rect 78673 142566 82156 142568
rect 78673 142563 78739 142566
rect 505001 139906 505067 139909
rect 501860 139904 505067 139906
rect 501860 139848 505006 139904
rect 505062 139848 505067 139904
rect 501860 139846 505067 139848
rect 505001 139843 505067 139846
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 79409 130930 79475 130933
rect 79409 130928 82156 130930
rect 79409 130872 79414 130928
rect 79470 130872 82156 130928
rect 79409 130870 82156 130872
rect 79409 130867 79475 130870
rect 504449 129026 504515 129029
rect 501860 129024 504515 129026
rect 501860 128968 504454 129024
rect 504510 128968 504515 129024
rect 501860 128966 504515 128968
rect 504449 128963 504515 128966
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 79317 119370 79383 119373
rect 79317 119368 82156 119370
rect 79317 119312 79322 119368
rect 79378 119312 82156 119368
rect 79317 119310 82156 119312
rect 79317 119307 79383 119310
rect 504357 118146 504423 118149
rect 501860 118144 504423 118146
rect 501860 118088 504362 118144
rect 504418 118088 504423 118144
rect 501860 118086 504423 118088
rect 504357 118083 504423 118086
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 505737 107402 505803 107405
rect 501860 107400 505803 107402
rect 501860 107344 505742 107400
rect 505798 107344 505803 107400
rect 501860 107342 505803 107344
rect 505737 107339 505803 107342
rect 583520 99636 584960 99876
rect 88517 96658 88583 96661
rect 89161 96658 89227 96661
rect 88517 96656 89227 96658
rect 88517 96600 88522 96656
rect 88578 96600 89166 96656
rect 89222 96600 89227 96656
rect 88517 96598 89227 96600
rect 88517 96595 88583 96598
rect 89161 96595 89227 96598
rect 101581 96658 101647 96661
rect 101949 96658 102015 96661
rect 101581 96656 102015 96658
rect 101581 96600 101586 96656
rect 101642 96600 101954 96656
rect 102010 96600 102015 96656
rect 101581 96598 102015 96600
rect 101581 96595 101647 96598
rect 101949 96595 102015 96598
rect 104065 96658 104131 96661
rect 104525 96658 104591 96661
rect 104065 96656 104591 96658
rect 104065 96600 104070 96656
rect 104126 96600 104530 96656
rect 104586 96600 104591 96656
rect 104065 96598 104591 96600
rect 104065 96595 104131 96598
rect 104525 96595 104591 96598
rect 105537 96658 105603 96661
rect 106181 96658 106247 96661
rect 105537 96656 106247 96658
rect 105537 96600 105542 96656
rect 105598 96600 106186 96656
rect 106242 96600 106247 96656
rect 105537 96598 106247 96600
rect 105537 96595 105603 96598
rect 106181 96595 106247 96598
rect 106641 96658 106707 96661
rect 107101 96658 107167 96661
rect 106641 96656 107167 96658
rect 106641 96600 106646 96656
rect 106702 96600 107106 96656
rect 107162 96600 107167 96656
rect 106641 96598 107167 96600
rect 106641 96595 106707 96598
rect 107101 96595 107167 96598
rect 108297 96658 108363 96661
rect 108757 96658 108823 96661
rect 108297 96656 108823 96658
rect 108297 96600 108302 96656
rect 108358 96600 108762 96656
rect 108818 96600 108823 96656
rect 108297 96598 108823 96600
rect 108297 96595 108363 96598
rect 108757 96595 108823 96598
rect 124397 96658 124463 96661
rect 124949 96658 125015 96661
rect 124397 96656 125015 96658
rect 124397 96600 124402 96656
rect 124458 96600 124954 96656
rect 125010 96600 125015 96656
rect 124397 96598 125015 96600
rect 124397 96595 124463 96598
rect 124949 96595 125015 96598
rect 142337 96658 142403 96661
rect 142889 96658 142955 96661
rect 142337 96656 142955 96658
rect 142337 96600 142342 96656
rect 142398 96600 142894 96656
rect 142950 96600 142955 96656
rect 142337 96598 142955 96600
rect 142337 96595 142403 96598
rect 142889 96595 142955 96598
rect 153377 96658 153443 96661
rect 154021 96658 154087 96661
rect 153377 96656 154087 96658
rect 153377 96600 153382 96656
rect 153438 96600 154026 96656
rect 154082 96600 154087 96656
rect 153377 96598 154087 96600
rect 153377 96595 153443 96598
rect 154021 96595 154087 96598
rect 200021 96658 200087 96661
rect 200297 96658 200363 96661
rect 200021 96656 200363 96658
rect 200021 96600 200026 96656
rect 200082 96600 200302 96656
rect 200358 96600 200363 96656
rect 200021 96598 200363 96600
rect 200021 96595 200087 96598
rect 200297 96595 200363 96598
rect 206553 96658 206619 96661
rect 206921 96658 206987 96661
rect 206553 96656 206987 96658
rect 206553 96600 206558 96656
rect 206614 96600 206926 96656
rect 206982 96600 206987 96656
rect 206553 96598 206987 96600
rect 206553 96595 206619 96598
rect 206921 96595 206987 96598
rect 207289 96658 207355 96661
rect 207749 96658 207815 96661
rect 207289 96656 207815 96658
rect 207289 96600 207294 96656
rect 207350 96600 207754 96656
rect 207810 96600 207815 96656
rect 207289 96598 207815 96600
rect 207289 96595 207355 96598
rect 207749 96595 207815 96598
rect 208853 96658 208919 96661
rect 209497 96658 209563 96661
rect 208853 96656 209563 96658
rect 208853 96600 208858 96656
rect 208914 96600 209502 96656
rect 209558 96600 209563 96656
rect 208853 96598 209563 96600
rect 208853 96595 208919 96598
rect 209497 96595 209563 96598
rect 213085 96658 213151 96661
rect 213729 96658 213795 96661
rect 213085 96656 213795 96658
rect 213085 96600 213090 96656
rect 213146 96600 213734 96656
rect 213790 96600 213795 96656
rect 213085 96598 213795 96600
rect 213085 96595 213151 96598
rect 213729 96595 213795 96598
rect 310145 96658 310211 96661
rect 310329 96658 310395 96661
rect 310145 96656 310395 96658
rect 310145 96600 310150 96656
rect 310206 96600 310334 96656
rect 310390 96600 310395 96656
rect 310145 96598 310395 96600
rect 310145 96595 310211 96598
rect 310329 96595 310395 96598
rect 328085 96658 328151 96661
rect 328269 96658 328335 96661
rect 328085 96656 328335 96658
rect 328085 96600 328090 96656
rect 328146 96600 328274 96656
rect 328330 96600 328335 96656
rect 328085 96598 328335 96600
rect 328085 96595 328151 96598
rect 328269 96595 328335 96598
rect 332317 96658 332383 96661
rect 332501 96658 332567 96661
rect 332317 96656 332567 96658
rect 332317 96600 332322 96656
rect 332378 96600 332506 96656
rect 332562 96600 332567 96656
rect 332317 96598 332567 96600
rect 332317 96595 332383 96598
rect 332501 96595 332567 96598
rect 379237 96658 379303 96661
rect 379421 96658 379487 96661
rect 379237 96656 379487 96658
rect 379237 96600 379242 96656
rect 379298 96600 379426 96656
rect 379482 96600 379487 96656
rect 379237 96598 379487 96600
rect 379237 96595 379303 96598
rect 379421 96595 379487 96598
rect 421925 96658 421991 96661
rect 422109 96658 422175 96661
rect 421925 96656 422175 96658
rect 421925 96600 421930 96656
rect 421986 96600 422114 96656
rect 422170 96600 422175 96656
rect 421925 96598 422175 96600
rect 421925 96595 421991 96598
rect 422109 96595 422175 96598
rect 433057 96658 433123 96661
rect 433241 96658 433307 96661
rect 433057 96656 433307 96658
rect 433057 96600 433062 96656
rect 433118 96600 433246 96656
rect 433302 96600 433307 96656
rect 433057 96598 433307 96600
rect 433057 96595 433123 96598
rect 433241 96595 433307 96598
rect 439865 96658 439931 96661
rect 440049 96658 440115 96661
rect 439865 96656 440115 96658
rect 439865 96600 439870 96656
rect 439926 96600 440054 96656
rect 440110 96600 440115 96656
rect 439865 96598 440115 96600
rect 439865 96595 439931 96598
rect 440049 96595 440115 96598
rect 450997 96658 451063 96661
rect 451181 96658 451247 96661
rect 450997 96656 451247 96658
rect 450997 96600 451002 96656
rect 451058 96600 451186 96656
rect 451242 96600 451247 96656
rect 450997 96598 451247 96600
rect 450997 96595 451063 96598
rect 451181 96595 451247 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 255865 87138 255931 87141
rect 411069 87138 411135 87141
rect 255270 87136 255931 87138
rect 255270 87080 255870 87136
rect 255926 87080 255931 87136
rect 255270 87078 255931 87080
rect 226517 87002 226583 87005
rect 226977 87002 227043 87005
rect 226517 87000 227043 87002
rect 226517 86944 226522 87000
rect 226578 86944 226982 87000
rect 227038 86944 227043 87000
rect 226517 86942 227043 86944
rect 255270 87002 255330 87078
rect 255865 87075 255931 87078
rect 410934 87136 411135 87138
rect 410934 87080 411074 87136
rect 411130 87080 411135 87136
rect 410934 87078 411135 87080
rect 410934 87005 410994 87078
rect 411069 87075 411135 87078
rect 255405 87002 255471 87005
rect 255270 87000 255471 87002
rect 255270 86944 255410 87000
rect 255466 86944 255471 87000
rect 255270 86942 255471 86944
rect 226517 86939 226583 86942
rect 226977 86939 227043 86942
rect 255405 86939 255471 86942
rect 327993 87002 328059 87005
rect 328177 87002 328243 87005
rect 327993 87000 328243 87002
rect 327993 86944 327998 87000
rect 328054 86944 328182 87000
rect 328238 86944 328243 87000
rect 327993 86942 328243 86944
rect 327993 86939 328059 86942
rect 328177 86939 328243 86942
rect 350257 87002 350323 87005
rect 350441 87002 350507 87005
rect 350257 87000 350507 87002
rect 350257 86944 350262 87000
rect 350318 86944 350446 87000
rect 350502 86944 350507 87000
rect 350257 86942 350507 86944
rect 410934 87000 411043 87005
rect 410934 86944 410982 87000
rect 411038 86944 411043 87000
rect 410934 86942 411043 86944
rect 350257 86939 350323 86942
rect 350441 86939 350507 86942
rect 410977 86939 411043 86942
rect 428641 85506 428707 85509
rect 428917 85506 428983 85509
rect 428641 85504 428983 85506
rect 428641 85448 428646 85504
rect 428702 85448 428922 85504
rect 428978 85448 428983 85504
rect 428641 85446 428983 85448
rect 428641 85443 428707 85446
rect 428917 85443 428983 85446
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 207013 77346 207079 77349
rect 207197 77346 207263 77349
rect 261201 77346 261267 77349
rect 207013 77344 207263 77346
rect 207013 77288 207018 77344
rect 207074 77288 207202 77344
rect 207258 77288 207263 77344
rect 207013 77286 207263 77288
rect 207013 77283 207079 77286
rect 207197 77283 207263 77286
rect 260974 77344 261267 77346
rect 260974 77288 261206 77344
rect 261262 77288 261267 77344
rect 260974 77286 261267 77288
rect 260833 77210 260899 77213
rect 260974 77210 261034 77286
rect 261201 77283 261267 77286
rect 390185 77346 390251 77349
rect 390369 77346 390435 77349
rect 390185 77344 390435 77346
rect 390185 77288 390190 77344
rect 390246 77288 390374 77344
rect 390430 77288 390435 77344
rect 390185 77286 390435 77288
rect 390185 77283 390251 77286
rect 390369 77283 390435 77286
rect 260833 77208 261034 77210
rect 260833 77152 260838 77208
rect 260894 77152 261034 77208
rect 260833 77150 261034 77152
rect 260833 77147 260899 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 229001 75850 229067 75853
rect 229277 75850 229343 75853
rect 229001 75848 229343 75850
rect 229001 75792 229006 75848
rect 229062 75792 229282 75848
rect 229338 75792 229343 75848
rect 229001 75790 229343 75792
rect 229001 75787 229067 75790
rect 229277 75787 229343 75790
rect 230657 67690 230723 67693
rect 230841 67690 230907 67693
rect 230657 67688 230907 67690
rect 230657 67632 230662 67688
rect 230718 67632 230846 67688
rect 230902 67632 230907 67688
rect 230657 67630 230907 67632
rect 230657 67627 230723 67630
rect 230841 67627 230907 67630
rect 332409 67690 332475 67693
rect 332593 67690 332659 67693
rect 332409 67688 332659 67690
rect 332409 67632 332414 67688
rect 332470 67632 332598 67688
rect 332654 67632 332659 67688
rect 332409 67630 332659 67632
rect 332409 67627 332475 67630
rect 332593 67627 332659 67630
rect 164325 67554 164391 67557
rect 164190 67552 164391 67554
rect 164190 67496 164330 67552
rect 164386 67496 164391 67552
rect 164190 67494 164391 67496
rect 164190 67418 164250 67494
rect 164325 67491 164391 67494
rect 164417 67418 164483 67421
rect 164190 67416 164483 67418
rect 164190 67360 164422 67416
rect 164478 67360 164483 67416
rect 164190 67358 164483 67360
rect 164417 67355 164483 67358
rect 229001 66330 229067 66333
rect 229277 66330 229343 66333
rect 229001 66328 229343 66330
rect 229001 66272 229006 66328
rect 229062 66272 229282 66328
rect 229338 66272 229343 66328
rect 229001 66270 229343 66272
rect 229001 66267 229067 66270
rect 229277 66267 229343 66270
rect 321185 66330 321251 66333
rect 321369 66330 321435 66333
rect 321185 66328 321435 66330
rect 321185 66272 321190 66328
rect 321246 66272 321374 66328
rect 321430 66272 321435 66328
rect 321185 66270 321435 66272
rect 321185 66267 321251 66270
rect 321369 66267 321435 66270
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 350349 54090 350415 54093
rect 350214 54088 350415 54090
rect 350214 54032 350354 54088
rect 350410 54032 350415 54088
rect 350214 54030 350415 54032
rect 350214 53954 350274 54030
rect 350349 54027 350415 54030
rect 350349 53954 350415 53957
rect 350214 53952 350415 53954
rect 350214 53896 350354 53952
rect 350410 53896 350415 53952
rect 350214 53894 350415 53896
rect 350349 53891 350415 53894
rect 350349 53818 350415 53821
rect 350533 53818 350599 53821
rect 350349 53816 350599 53818
rect 350349 53760 350354 53816
rect 350410 53760 350538 53816
rect 350594 53760 350599 53816
rect 350349 53758 350599 53760
rect 350349 53755 350415 53758
rect 350533 53755 350599 53758
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 175365 48242 175431 48245
rect 175230 48240 175431 48242
rect 175230 48184 175370 48240
rect 175426 48184 175431 48240
rect 175230 48182 175431 48184
rect 175230 48106 175290 48182
rect 175365 48179 175431 48182
rect 248689 48242 248755 48245
rect 248965 48242 249031 48245
rect 248689 48240 249031 48242
rect 248689 48184 248694 48240
rect 248750 48184 248970 48240
rect 249026 48184 249031 48240
rect 248689 48182 249031 48184
rect 248689 48179 248755 48182
rect 248965 48179 249031 48182
rect 175457 48106 175523 48109
rect 175230 48104 175523 48106
rect 175230 48048 175462 48104
rect 175518 48048 175523 48104
rect 175230 48046 175523 48048
rect 175457 48043 175523 48046
rect 321185 46882 321251 46885
rect 321318 46882 321324 46884
rect 321185 46880 321324 46882
rect 321185 46824 321190 46880
rect 321246 46824 321324 46880
rect 321185 46822 321324 46824
rect 321185 46819 321251 46822
rect 321318 46820 321324 46822
rect 321388 46820 321394 46884
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 111793 38722 111859 38725
rect 272057 38722 272123 38725
rect 272241 38722 272307 38725
rect 111793 38720 111994 38722
rect 111793 38664 111798 38720
rect 111854 38664 111994 38720
rect 111793 38662 111994 38664
rect 111793 38659 111859 38662
rect 111793 38586 111859 38589
rect 111934 38586 111994 38662
rect 272057 38720 272307 38722
rect 272057 38664 272062 38720
rect 272118 38664 272246 38720
rect 272302 38664 272307 38720
rect 272057 38662 272307 38664
rect 272057 38659 272123 38662
rect 272241 38659 272307 38662
rect 111793 38584 111994 38586
rect 111793 38528 111798 38584
rect 111854 38528 111994 38584
rect 111793 38526 111994 38528
rect 111793 38523 111859 38526
rect 321185 37362 321251 37365
rect 321318 37362 321324 37364
rect 321185 37360 321324 37362
rect 321185 37304 321190 37360
rect 321246 37304 321324 37360
rect 321185 37302 321324 37304
rect 321185 37299 321251 37302
rect 321318 37300 321324 37302
rect 321388 37300 321394 37364
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 271781 29066 271847 29069
rect 271965 29066 272031 29069
rect 271781 29064 272031 29066
rect 271781 29008 271786 29064
rect 271842 29008 271970 29064
rect 272026 29008 272031 29064
rect 271781 29006 272031 29008
rect 271781 29003 271847 29006
rect 271965 29003 272031 29006
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 31477 9754 31543 9757
rect 31661 9754 31727 9757
rect 31477 9752 31727 9754
rect 31477 9696 31482 9752
rect 31538 9696 31666 9752
rect 31722 9696 31727 9752
rect 31477 9694 31727 9696
rect 31477 9691 31543 9694
rect 31661 9691 31727 9694
rect -960 7170 480 7260
rect 4061 7170 4127 7173
rect -960 7168 4127 7170
rect -960 7112 4066 7168
rect 4122 7112 4127 7168
rect -960 7110 4127 7112
rect -960 7020 480 7110
rect 4061 7107 4127 7110
rect 583520 5796 584960 6036
<< via3 >>
rect 321324 46820 321388 46884
rect 321324 37300 321388 37364
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 602000 84204 624698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 602000 91404 631898
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 602000 95004 635498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 602000 98604 603098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 602000 102204 606698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 602000 109404 613898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 602000 113004 617498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 602000 116604 621098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 602000 120204 624698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 602000 127404 631898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 602000 131004 635498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 602000 134604 603098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 602000 138204 606698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 602000 145404 613898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 602000 149004 617498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 602000 152604 621098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 602000 156204 624698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 602000 163404 631898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 602000 167004 635498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 602000 170604 603098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 602000 174204 606698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 602000 181404 613898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 602000 185004 617498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 602000 188604 621098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 602000 192204 624698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 602000 199404 631898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 602000 203004 635498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 602000 206604 603098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 602000 210204 606698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 602000 217404 613898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 602000 221004 617498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 602000 224604 621098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 602000 228204 624698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 602000 235404 631898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 602000 239004 635498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 602000 242604 603098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 602000 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 602000 253404 613898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 602000 257004 617498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 602000 260604 621098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 602000 264204 624698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 602000 271404 631898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 602000 275004 635498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 602000 278604 603098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 602000 282204 606698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 602000 289404 613898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 602000 293004 617498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 602000 296604 621098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 602000 300204 624698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 602000 307404 631898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 602000 311004 635498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 602000 314604 603098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 602000 318204 606698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 602000 325404 613898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 602000 329004 617498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 602000 332604 621098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 602000 336204 624698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 602000 343404 631898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 602000 347004 635498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 602000 350604 603098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 602000 354204 606698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 602000 361404 613898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 602000 365004 617498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 602000 368604 621098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 602000 372204 624698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 602000 379404 631898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 602000 383004 635498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 602000 386604 603098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 602000 390204 606698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 602000 397404 613898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 602000 401004 617498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 602000 404604 621098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 602000 408204 624698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 602000 415404 631898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 602000 419004 635498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 602000 422604 603098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 602000 426204 606698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 602000 433404 613898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 602000 437004 617498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 602000 440604 621098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 602000 444204 624698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 602000 451404 631898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 602000 455004 635498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 602000 458604 603098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 602000 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 602000 469404 613898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 602000 473004 617498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 602000 476604 621098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 602000 480204 624698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 602000 487404 631898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 602000 491004 635498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 602000 494604 603098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 602000 498204 606698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 85254 84204 102000
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 92454 91404 102000
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 96054 95004 102000
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 99654 98604 102000
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 67254 102204 102000
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 74454 109404 102000
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 78054 113004 102000
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 81654 116604 102000
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 85254 120204 102000
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 92454 127404 102000
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 96054 131004 102000
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 99654 134604 102000
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 67254 138204 102000
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 74454 145404 102000
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 78054 149004 102000
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 81654 152604 102000
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 85254 156204 102000
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 92454 163404 102000
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 96054 167004 102000
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 99654 170604 102000
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 67254 174204 102000
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 74454 181404 102000
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 78054 185004 102000
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 81654 188604 102000
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 85254 192204 102000
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 92454 199404 102000
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 96054 203004 102000
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 99654 206604 102000
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 67254 210204 102000
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 74454 217404 102000
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 78054 221004 102000
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 81654 224604 102000
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 85254 228204 102000
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 92454 235404 102000
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 96054 239004 102000
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 99654 242604 102000
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 67254 246204 102000
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 74454 253404 102000
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 78054 257004 102000
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 81654 260604 102000
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 85254 264204 102000
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 92454 271404 102000
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 96054 275004 102000
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 99654 278604 102000
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 67254 282204 102000
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 102000
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 78054 293004 102000
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 81654 296604 102000
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 85254 300204 102000
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 92454 307404 102000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 96054 311004 102000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 99654 314604 102000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 67254 318204 102000
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 324804 74454 325404 102000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 321323 46884 321389 46885
rect 321323 46820 321324 46884
rect 321388 46820 321389 46884
rect 321323 46819 321389 46820
rect 321326 37365 321386 46819
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 321323 37364 321389 37365
rect 321323 37300 321324 37364
rect 321388 37300 321389 37364
rect 321323 37299 321389 37300
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 78054 329004 102000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 81654 332604 102000
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 85254 336204 102000
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 92454 343404 102000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 96054 347004 102000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 99654 350604 102000
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 67254 354204 102000
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 74454 361404 102000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 78054 365004 102000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 81654 368604 102000
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 85254 372204 102000
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 92454 379404 102000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 96054 383004 102000
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 99654 386604 102000
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 67254 390204 102000
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 74454 397404 102000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 78054 401004 102000
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 81654 404604 102000
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 85254 408204 102000
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 92454 415404 102000
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 96054 419004 102000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 99654 422604 102000
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 67254 426204 102000
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 74454 433404 102000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 78054 437004 102000
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 81654 440604 102000
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 85254 444204 102000
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 92454 451404 102000
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 96054 455004 102000
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 99654 458604 102000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 67254 462204 102000
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 74454 469404 102000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 78054 473004 102000
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 81654 476604 102000
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 85254 480204 102000
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 92454 487404 102000
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 96054 491004 102000
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 99654 494604 102000
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 67254 498204 102000
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use Ibtida_top_dffram_cv  mprj
timestamp 1607488137
transform 1 0 82000 0 1 102000
box 0 0 420000 500000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
