VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM
  CLASS BLOCK ;
  FOREIGN DFFRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 1012.325 BY 1023.045 ;
  PIN A[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.090 1019.045 575.370 1023.045 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.170 1019.045 965.450 1023.045 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 1019.045 141.130 1023.045 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 697.720 1012.325 698.320 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 825.560 1012.325 826.160 ;
    END
  END A[7]
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 618.330 1019.045 618.610 1023.045 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.450 1019.045 835.730 1023.045 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.970 1019.045 358.250 1023.045 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 632.440 1012.325 633.040 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.570 1019.045 661.850 1023.045 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 119.720 1012.325 120.320 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1008.410 1019.045 1008.690 1023.045 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.210 1019.045 401.490 1023.045 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 889.480 1012.325 890.080 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 1019.045 54.650 1023.045 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 1019.045 97.890 1023.045 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.210 1019.045 792.490 1023.045 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 1019.045 184.370 1023.045 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 183.640 1012.325 184.240 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 1019.045 10.490 1023.045 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 704.810 1019.045 705.090 1023.045 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 568.520 1012.325 569.120 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 531.850 1019.045 532.130 1023.045 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 953.400 1012.325 954.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 504.600 1012.325 505.200 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 55.800 1012.325 56.400 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 1019.045 270.850 1023.045 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 440.680 1012.325 441.280 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 376.760 1012.325 377.360 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 487.690 1019.045 487.970 1023.045 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 921.930 1019.045 922.210 1023.045 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.050 1019.045 748.330 1023.045 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 247.560 1012.325 248.160 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 444.450 1019.045 444.730 1023.045 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1008.325 312.840 1012.325 313.440 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.730 1019.045 315.010 1023.045 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 878.690 1019.045 878.970 1023.045 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1008.325 761.640 1012.325 762.240 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 1019.045 227.610 1023.045 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1006.480 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1006.480 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1006.480 1011.925 ;
      LAYER met1 ;
        RECT 2.830 10.640 1008.710 1012.080 ;
      LAYER met2 ;
        RECT 2.860 1018.765 9.930 1019.050 ;
        RECT 10.770 1018.765 54.090 1019.050 ;
        RECT 54.930 1018.765 97.330 1019.050 ;
        RECT 98.170 1018.765 140.570 1019.050 ;
        RECT 141.410 1018.765 183.810 1019.050 ;
        RECT 184.650 1018.765 227.050 1019.050 ;
        RECT 227.890 1018.765 270.290 1019.050 ;
        RECT 271.130 1018.765 314.450 1019.050 ;
        RECT 315.290 1018.765 357.690 1019.050 ;
        RECT 358.530 1018.765 400.930 1019.050 ;
        RECT 401.770 1018.765 444.170 1019.050 ;
        RECT 445.010 1018.765 487.410 1019.050 ;
        RECT 488.250 1018.765 531.570 1019.050 ;
        RECT 532.410 1018.765 574.810 1019.050 ;
        RECT 575.650 1018.765 618.050 1019.050 ;
        RECT 618.890 1018.765 661.290 1019.050 ;
        RECT 662.130 1018.765 704.530 1019.050 ;
        RECT 705.370 1018.765 747.770 1019.050 ;
        RECT 748.610 1018.765 791.930 1019.050 ;
        RECT 792.770 1018.765 835.170 1019.050 ;
        RECT 836.010 1018.765 878.410 1019.050 ;
        RECT 879.250 1018.765 921.650 1019.050 ;
        RECT 922.490 1018.765 964.890 1019.050 ;
        RECT 965.730 1018.765 1008.130 1019.050 ;
        RECT 2.860 4.280 1008.680 1018.765 ;
        RECT 3.410 4.000 45.810 4.280 ;
        RECT 46.650 4.000 89.050 4.280 ;
        RECT 89.890 4.000 132.290 4.280 ;
        RECT 133.130 4.000 175.530 4.280 ;
        RECT 176.370 4.000 218.770 4.280 ;
        RECT 219.610 4.000 262.930 4.280 ;
        RECT 263.770 4.000 306.170 4.280 ;
        RECT 307.010 4.000 349.410 4.280 ;
        RECT 350.250 4.000 392.650 4.280 ;
        RECT 393.490 4.000 435.890 4.280 ;
        RECT 436.730 4.000 479.130 4.280 ;
        RECT 479.970 4.000 523.290 4.280 ;
        RECT 524.130 4.000 566.530 4.280 ;
        RECT 567.370 4.000 609.770 4.280 ;
        RECT 610.610 4.000 653.010 4.280 ;
        RECT 653.850 4.000 696.250 4.280 ;
        RECT 697.090 4.000 740.410 4.280 ;
        RECT 741.250 4.000 783.650 4.280 ;
        RECT 784.490 4.000 826.890 4.280 ;
        RECT 827.730 4.000 870.130 4.280 ;
        RECT 870.970 4.000 913.370 4.280 ;
        RECT 914.210 4.000 956.610 4.280 ;
        RECT 957.450 4.000 1000.770 4.280 ;
        RECT 1001.610 4.000 1008.680 4.280 ;
      LAYER met3 ;
        RECT 4.000 966.640 1008.325 1012.005 ;
        RECT 4.400 965.240 1008.325 966.640 ;
        RECT 4.000 954.400 1008.325 965.240 ;
        RECT 4.000 953.000 1007.925 954.400 ;
        RECT 4.000 902.720 1008.325 953.000 ;
        RECT 4.400 901.320 1008.325 902.720 ;
        RECT 4.000 890.480 1008.325 901.320 ;
        RECT 4.000 889.080 1007.925 890.480 ;
        RECT 4.000 838.800 1008.325 889.080 ;
        RECT 4.400 837.400 1008.325 838.800 ;
        RECT 4.000 826.560 1008.325 837.400 ;
        RECT 4.000 825.160 1007.925 826.560 ;
        RECT 4.000 774.880 1008.325 825.160 ;
        RECT 4.400 773.480 1008.325 774.880 ;
        RECT 4.000 762.640 1008.325 773.480 ;
        RECT 4.000 761.240 1007.925 762.640 ;
        RECT 4.000 709.600 1008.325 761.240 ;
        RECT 4.400 708.200 1008.325 709.600 ;
        RECT 4.000 698.720 1008.325 708.200 ;
        RECT 4.000 697.320 1007.925 698.720 ;
        RECT 4.000 645.680 1008.325 697.320 ;
        RECT 4.400 644.280 1008.325 645.680 ;
        RECT 4.000 633.440 1008.325 644.280 ;
        RECT 4.000 632.040 1007.925 633.440 ;
        RECT 4.000 581.760 1008.325 632.040 ;
        RECT 4.400 580.360 1008.325 581.760 ;
        RECT 4.000 569.520 1008.325 580.360 ;
        RECT 4.000 568.120 1007.925 569.520 ;
        RECT 4.000 517.840 1008.325 568.120 ;
        RECT 4.400 516.440 1008.325 517.840 ;
        RECT 4.000 505.600 1008.325 516.440 ;
        RECT 4.000 504.200 1007.925 505.600 ;
        RECT 4.000 453.920 1008.325 504.200 ;
        RECT 4.400 452.520 1008.325 453.920 ;
        RECT 4.000 441.680 1008.325 452.520 ;
        RECT 4.000 440.280 1007.925 441.680 ;
        RECT 4.000 390.000 1008.325 440.280 ;
        RECT 4.400 388.600 1008.325 390.000 ;
        RECT 4.000 377.760 1008.325 388.600 ;
        RECT 4.000 376.360 1007.925 377.760 ;
        RECT 4.000 324.720 1008.325 376.360 ;
        RECT 4.400 323.320 1008.325 324.720 ;
        RECT 4.000 313.840 1008.325 323.320 ;
        RECT 4.000 312.440 1007.925 313.840 ;
        RECT 4.000 260.800 1008.325 312.440 ;
        RECT 4.400 259.400 1008.325 260.800 ;
        RECT 4.000 248.560 1008.325 259.400 ;
        RECT 4.000 247.160 1007.925 248.560 ;
        RECT 4.000 196.880 1008.325 247.160 ;
        RECT 4.400 195.480 1008.325 196.880 ;
        RECT 4.000 184.640 1008.325 195.480 ;
        RECT 4.000 183.240 1007.925 184.640 ;
        RECT 4.000 132.960 1008.325 183.240 ;
        RECT 4.400 131.560 1008.325 132.960 ;
        RECT 4.000 120.720 1008.325 131.560 ;
        RECT 4.000 119.320 1007.925 120.720 ;
        RECT 4.000 69.040 1008.325 119.320 ;
        RECT 4.400 67.640 1008.325 69.040 ;
        RECT 4.000 56.800 1008.325 67.640 ;
        RECT 4.000 55.400 1007.925 56.800 ;
        RECT 4.000 10.715 1008.325 55.400 ;
      LAYER met4 ;
        RECT 21.040 10.640 944.240 1012.080 ;
      LAYER met5 ;
        RECT 5.520 179.670 1006.480 947.170 ;
  END
END DFFRAM
END LIBRARY

