VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Ibtida_top_dffram_cv
  CLASS BLOCK ;
  FOREIGN Ibtida_top_dffram_cv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2100.000 BY 2500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 2496.000 108.930 2500.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1015.960 2100.000 1016.560 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.570 2496.000 1627.850 2500.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1645.050 0.000 1645.330 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1391.320 4.000 1391.920 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 2496.000 232.210 2500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1232.890 2496.000 1233.170 2500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1967.050 0.000 1967.330 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.970 2496.000 887.250 2500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 650.120 2100.000 650.720 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.770 2496.000 1591.050 2500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 66.680 2100.000 67.280 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1947.560 2100.000 1948.160 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2359.640 4.000 2360.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.330 0.000 1929.610 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.090 2496.000 874.370 2500.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.450 2496.000 973.730 2500.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 2496.000 824.690 2500.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2001.960 2100.000 2002.560 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2035.130 2496.000 2035.410 2500.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1436.200 2100.000 1436.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2422.200 2100.000 2422.800 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 2496.000 1195.450 2500.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 182.250 2496.000 182.530 2500.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.570 2496.000 454.850 2500.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1417.160 2100.000 1417.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2203.240 2100.000 2203.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1161.480 2100.000 1162.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 478.490 2496.000 478.770 2500.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 340.040 2100.000 340.640 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1124.760 2100.000 1125.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1596.290 0.000 1596.570 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 564.970 2496.000 565.250 2500.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2166.520 2100.000 2167.120 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1504.290 2496.000 1504.570 2500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1657.930 0.000 1658.210 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2458.920 2100.000 2459.520 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1899.890 2496.000 1900.170 2500.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1990.970 0.000 1991.250 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 2496.000 1146.690 2500.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1200.690 0.000 1200.970 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.290 2496.000 170.570 2500.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2468.440 4.000 2469.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 4.000 1227.360 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 2496.000 71.210 2500.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1508.280 2100.000 1508.880 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1998.330 2496.000 1998.610 2500.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 639.490 2496.000 639.770 2500.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2096.770 2496.000 2097.050 2500.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.570 0.000 1052.850 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1702.090 2496.000 1702.370 2500.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 516.210 2496.000 516.490 2500.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.850 2496.000 417.130 2500.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1534.650 0.000 1534.930 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1608.250 0.000 1608.530 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1362.760 2100.000 1363.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2257.640 2100.000 2258.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2140.680 4.000 2141.280 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.650 2496.000 1281.930 2500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.490 0.000 1237.770 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1794.090 0.000 1794.370 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1564.040 2100.000 1564.640 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1848.280 4.000 1848.880 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 528.170 2496.000 528.450 2500.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.800 4.000 1246.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2348.760 2100.000 2349.360 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 948.610 2496.000 948.890 2500.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 522.280 2100.000 522.880 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.330 2496.000 1331.610 2500.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.130 2496.000 862.410 2500.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 2496.000 355.490 2500.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 632.440 2100.000 633.040 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2312.040 2100.000 2312.640 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1368.130 2496.000 1368.410 2500.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 924.840 2100.000 925.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1751.770 2496.000 1752.050 2500.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1225.530 0.000 1225.810 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.890 2496.000 244.170 2500.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 467.880 2100.000 468.480 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 121.080 2100.000 121.680 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.450 2496.000 651.730 2500.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1862.170 2496.000 1862.450 2500.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1405.850 2496.000 1406.130 2500.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1719.570 0.000 1719.850 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1044.520 4.000 1045.120 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 777.960 2100.000 778.560 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1986.370 2496.000 1986.650 2500.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1792.520 4.000 1793.120 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1830.890 0.000 1831.170 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1954.170 0.000 1954.450 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 676.290 2496.000 676.570 2500.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1565.930 2496.000 1566.210 2500.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2487.480 4.000 2488.080 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.840 4.000 2013.440 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1920.360 4.000 1920.960 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1070.360 2100.000 1070.960 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 29.960 2100.000 30.560 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1928.520 2100.000 1929.120 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 2496.000 59.250 2500.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2476.600 2100.000 2477.200 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 2496.000 812.730 2500.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.370 2496.000 491.650 2500.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2003.850 0.000 2004.130 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.890 2496.000 1739.170 2500.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 613.400 2100.000 614.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2275.320 2100.000 2275.920 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1308.360 2100.000 1308.960 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1672.840 2100.000 1673.440 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 701.130 2496.000 701.410 2500.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.160 4.000 1519.760 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 595.720 2100.000 596.320 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.650 2496.000 614.930 2500.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1701.400 4.000 1702.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2331.080 2100.000 2331.680 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1089.400 2100.000 1090.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1891.800 2100.000 1892.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.490 2496.000 1467.770 2500.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1993.800 4.000 1994.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2303.880 4.000 2304.480 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2056.360 2100.000 2056.960 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1783.000 2100.000 1783.600 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2048.200 4.000 2048.800 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.530 2496.000 1294.810 2500.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2268.520 4.000 2269.120 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 541.320 2100.000 541.920 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1319.370 2496.000 1319.650 2500.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2450.760 4.000 2451.360 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1744.410 0.000 1744.690 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.330 2496.000 1492.610 2500.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1837.400 2100.000 1838.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1271.640 2100.000 1272.240 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1553.970 2496.000 1554.250 2500.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2011.210 2496.000 2011.490 2500.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2220.920 2100.000 2221.520 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2294.360 2100.000 2294.960 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2077.450 0.000 2077.730 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1602.730 2496.000 1603.010 2500.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 194.520 2100.000 195.120 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1541.090 2496.000 1541.370 2500.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.490 0.000 1398.770 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1033.640 2100.000 1034.240 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2322.920 4.000 2323.520 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1885.000 4.000 1885.600 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2385.480 2100.000 2386.080 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1306.490 2496.000 1306.770 2500.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.370 0.000 1756.650 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 2496.000 132.850 2500.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.010 2496.000 392.290 2500.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 888.120 2100.000 888.720 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 322.360 2100.000 322.960 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1942.210 0.000 1942.490 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1490.600 2100.000 1491.200 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1731.530 0.000 1731.810 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 47.640 2100.000 48.240 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2239.960 2100.000 2240.560 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 960.570 2496.000 960.850 2500.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2158.360 4.000 2158.960 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1707.610 0.000 1707.890 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.330 2496.000 503.610 2500.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2053.530 0.000 2053.810 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.650 2496.000 775.930 2500.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1800.530 2496.000 1800.810 2500.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1354.600 4.000 1355.200 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.050 2496.000 380.330 2500.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 578.040 2100.000 578.640 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1976.120 4.000 1976.720 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1509.810 0.000 1510.090 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1545.000 2100.000 1545.600 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.720 4.000 1446.320 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.690 0.000 1039.970 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1979.010 0.000 1979.290 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 157.800 2100.000 158.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1217.240 2100.000 1217.840 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2103.960 4.000 2104.560 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2030.520 4.000 2031.120 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1948.650 2496.000 1948.930 2500.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1126.170 0.000 1126.450 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.170 2496.000 22.450 2500.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.010 0.000 1312.290 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1555.880 4.000 1556.480 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1850.210 2496.000 1850.490 2500.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2367.800 2100.000 2368.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1496.930 0.000 1497.210 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 905.800 2100.000 906.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1198.200 2100.000 1198.800 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1720.440 4.000 1721.040 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.490 2496.000 800.770 2500.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.610 2496.000 281.890 2500.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1442.650 2496.000 1442.930 2500.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 559.000 2100.000 559.600 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1842.850 0.000 1843.130 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1208.050 2496.000 1208.330 2500.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.970 2496.000 1393.250 2500.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 553.010 2496.000 553.290 2500.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1583.410 0.000 1583.690 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1874.120 2100.000 1874.720 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.050 2496.000 1047.330 2500.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2093.080 2100.000 2093.680 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.850 2496.000 578.130 2500.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1647.000 4.000 1647.600 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 814.680 2100.000 815.280 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2184.200 2100.000 2184.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1453.880 2100.000 1454.480 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1664.680 4.000 1665.280 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 996.920 2100.000 997.520 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 979.240 2100.000 979.840 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.720 4.000 1684.320 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1578.810 2496.000 1579.090 2500.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 102.040 2100.000 102.640 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 669.160 2100.000 669.760 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 413.480 2100.000 414.080 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1746.280 2100.000 1746.880 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 2496.000 219.330 2500.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2431.720 4.000 2432.320 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1652.410 2496.000 1652.690 2500.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1516.250 2496.000 1516.530 2500.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1472.920 2100.000 1473.520 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.970 2496.000 726.250 2500.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.930 2496.000 1060.210 2500.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2072.850 2496.000 2073.130 2500.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.530 2496.000 305.810 2500.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2231.800 4.000 2232.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2038.680 2100.000 2039.280 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1763.730 2496.000 1764.010 2500.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1356.170 2496.000 1356.450 2500.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 851.400 2100.000 852.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.930 0.000 991.210 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1910.840 2100.000 1911.440 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2040.650 0.000 2040.930 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1256.810 2496.000 1257.090 2500.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1252.600 2100.000 1253.200 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1615.610 2496.000 1615.890 2500.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1448.170 0.000 1448.450 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1484.970 0.000 1485.250 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1010.250 2496.000 1010.530 2500.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1289.320 2100.000 1289.920 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1892.530 0.000 1892.810 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 212.200 2100.000 212.800 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2028.690 0.000 2028.970 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.170 2496.000 689.450 2500.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2023.170 2496.000 2023.450 2500.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1769.250 0.000 1769.530 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 705.880 2100.000 706.480 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1361.690 0.000 1361.970 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1689.210 2496.000 1689.490 2500.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 4.000 1318.480 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1345.080 2100.000 1345.680 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1385.610 0.000 1385.890 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1939.400 4.000 1940.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2286.200 4.000 2286.800 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2396.360 4.000 2396.960 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1180.520 2100.000 1181.120 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 2496.000 738.210 2500.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1143.800 2100.000 1144.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2065.490 0.000 2065.770 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.570 2496.000 293.850 2500.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1961.530 2496.000 1961.810 2500.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.010 2496.000 1887.290 2500.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 2496.000 34.410 2500.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1902.680 4.000 1903.280 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1856.440 2100.000 1857.040 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.090 2496.000 1035.370 2500.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.930 0.000 830.210 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1399.480 2100.000 1400.080 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1052.680 2100.000 1053.280 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1965.240 2100.000 1965.840 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 923.770 2496.000 924.050 2500.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1600.760 2100.000 1601.360 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.730 2496.000 936.010 2500.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.450 2496.000 1479.730 2500.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1460.130 0.000 1460.410 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2249.480 4.000 2250.080 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.330 2496.000 664.610 2500.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.530 2496.000 1133.810 2500.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 723.560 2100.000 724.160 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.050 2496.000 541.330 2500.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1417.810 2496.000 1418.090 2500.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 248.920 2100.000 249.520 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 10.920 2100.000 11.520 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2403.160 2100.000 2403.760 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 431.160 2100.000 431.760 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1714.050 2496.000 1714.330 2500.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1806.050 0.000 1806.330 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 741.240 2100.000 741.840 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 833.720 2100.000 834.320 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1819.720 2100.000 1820.320 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1220.010 2496.000 1220.290 2500.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.760 4.000 1465.360 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1326.040 2100.000 1326.640 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.210 2496.000 1183.490 2500.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 504.600 2100.000 505.200 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1865.960 4.000 1866.560 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1728.600 2100.000 1729.200 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 175.480 2100.000 176.080 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.050 0.000 1139.330 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 376.760 2100.000 377.360 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.010 0.000 1151.290 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1521.770 0.000 1522.050 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1904.490 0.000 1904.770 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 84.360 2100.000 84.960 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.690 2496.000 441.970 2500.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.730 2496.000 269.010 2500.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 2496.000 46.370 2500.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.160 4.000 1281.760 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1763.960 2100.000 1764.560 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2112.120 2100.000 2112.720 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1838.250 2496.000 1838.530 2500.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1800.680 2100.000 1801.280 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2377.320 4.000 2377.920 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 285.640 2100.000 286.240 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.690 2496.000 1775.970 2500.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1655.160 2100.000 1655.760 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 869.080 2100.000 869.680 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.730 2496.000 1097.010 2500.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1244.850 2496.000 1245.130 2500.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.810 2496.000 751.090 2500.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1726.930 2496.000 1727.210 2500.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1527.320 2100.000 1527.920 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.090 2496.000 368.370 2500.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2048.010 2496.000 2048.290 2500.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 2496.000 330.650 2500.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1529.130 2496.000 1529.410 2500.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2067.240 4.000 2067.840 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2019.640 2100.000 2020.240 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 2496.000 405.170 2500.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2084.920 4.000 2085.520 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.370 2496.000 997.650 2500.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1188.730 0.000 1189.010 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 961.560 2100.000 962.160 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1669.890 0.000 1670.170 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.050 2496.000 1875.330 2500.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1573.560 4.000 1574.160 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2147.480 2100.000 2148.080 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2121.640 4.000 2122.240 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1454.610 2496.000 1454.890 2500.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1813.410 2496.000 1813.690 2500.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2212.760 4.000 2213.360 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 760.280 2100.000 760.880 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.530 2496.000 466.810 2500.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 2496.000 1084.130 2500.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1636.120 2100.000 1636.720 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.410 2496.000 318.690 2500.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2195.080 4.000 2195.680 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 2496.000 84.090 2500.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 485.560 2100.000 486.160 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.690 2496.000 1269.970 2500.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 797.000 2100.000 797.600 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1984.280 2100.000 1984.880 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2059.970 2496.000 2060.250 2500.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 303.320 2100.000 303.920 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1738.120 4.000 1738.720 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 229.880 2100.000 230.480 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.290 2496.000 837.570 2500.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 394.440 2100.000 395.040 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1665.290 2496.000 1665.570 2500.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.010 2496.000 1381.290 2500.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1818.010 0.000 1818.290 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 138.760 2100.000 139.360 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1610.280 4.000 1610.880 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.090 0.000 1472.370 4.000 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2414.040 4.000 2414.640 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 849.250 2496.000 849.530 2500.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1263.480 4.000 1264.080 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2129.800 2100.000 2130.400 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 4.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.130 2496.000 195.410 2500.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 2496.000 9.570 2500.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1121.570 2496.000 1121.850 2500.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 2496.000 120.890 2500.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.850 2496.000 1912.130 2500.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.770 2496.000 1430.050 2500.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 686.840 2100.000 687.440 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1153.320 4.000 1153.920 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1022.210 2496.000 1022.490 2500.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1973.490 2496.000 1973.770 2500.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1501.480 4.000 1502.080 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 266.600 2100.000 267.200 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1709.560 2100.000 1710.160 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.410 2496.000 985.690 2500.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.690 2496.000 602.970 2500.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1691.880 2100.000 1692.480 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.890 2496.000 1072.170 2500.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1781.210 0.000 1781.490 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 942.520 2100.000 943.120 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1373.650 0.000 1373.930 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.890 2496.000 911.170 2500.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.810 0.000 1349.090 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.090 0.000 1633.370 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 2496.000 257.050 2500.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.920 4.000 1337.520 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1936.690 2496.000 1936.970 2500.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1924.730 2496.000 1925.010 2500.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2439.880 2100.000 2440.480 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1677.250 2496.000 1677.530 2500.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.090 2496.000 207.370 2500.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1957.080 4.000 1957.680 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 2496.000 1158.650 2500.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1581.720 2100.000 1582.320 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1618.440 2100.000 1619.040 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 2496.000 145.730 2500.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 357.720 2100.000 358.320 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 450.200 2100.000 450.800 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1694.730 0.000 1695.010 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1380.440 2100.000 1381.040 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1855.730 0.000 1856.010 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.330 2496.000 1170.610 2500.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.610 2496.000 787.890 2500.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1788.570 2496.000 1788.850 2500.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.930 2496.000 899.210 2500.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.370 0.000 1917.650 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2090.330 0.000 2090.610 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.410 2496.000 157.690 2500.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.810 2496.000 2085.090 2500.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1825.370 2496.000 1825.650 2500.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.730 2496.000 430.010 2500.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.010 2496.000 714.290 2500.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1621.130 0.000 1621.410 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.160 4.000 1757.760 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.810 2496.000 590.090 2500.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1811.560 4.000 1812.160 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2075.400 2100.000 2076.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.770 2496.000 763.050 2500.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 2496.000 96.050 2500.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.530 2496.000 627.810 2500.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1640.450 2496.000 1640.730 2500.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1343.290 2496.000 1343.570 2500.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.250 2496.000 343.530 2500.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1175.850 0.000 1176.130 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2340.600 4.000 2341.200 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1234.920 2100.000 1235.520 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.690 2496.000 1108.970 2500.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1107.080 2100.000 1107.680 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2489.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2489.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2094.380 2488.885 ;
      LAYER met1 ;
        RECT 5.520 4.460 2097.070 2489.040 ;
      LAYER met2 ;
        RECT 8.840 2495.720 9.010 2496.010 ;
        RECT 9.850 2495.720 21.890 2496.010 ;
        RECT 22.730 2495.720 33.850 2496.010 ;
        RECT 34.690 2495.720 45.810 2496.010 ;
        RECT 46.650 2495.720 58.690 2496.010 ;
        RECT 59.530 2495.720 70.650 2496.010 ;
        RECT 71.490 2495.720 83.530 2496.010 ;
        RECT 84.370 2495.720 95.490 2496.010 ;
        RECT 96.330 2495.720 108.370 2496.010 ;
        RECT 109.210 2495.720 120.330 2496.010 ;
        RECT 121.170 2495.720 132.290 2496.010 ;
        RECT 133.130 2495.720 145.170 2496.010 ;
        RECT 146.010 2495.720 157.130 2496.010 ;
        RECT 157.970 2495.720 170.010 2496.010 ;
        RECT 170.850 2495.720 181.970 2496.010 ;
        RECT 182.810 2495.720 194.850 2496.010 ;
        RECT 195.690 2495.720 206.810 2496.010 ;
        RECT 207.650 2495.720 218.770 2496.010 ;
        RECT 219.610 2495.720 231.650 2496.010 ;
        RECT 232.490 2495.720 243.610 2496.010 ;
        RECT 244.450 2495.720 256.490 2496.010 ;
        RECT 257.330 2495.720 268.450 2496.010 ;
        RECT 269.290 2495.720 281.330 2496.010 ;
        RECT 282.170 2495.720 293.290 2496.010 ;
        RECT 294.130 2495.720 305.250 2496.010 ;
        RECT 306.090 2495.720 318.130 2496.010 ;
        RECT 318.970 2495.720 330.090 2496.010 ;
        RECT 330.930 2495.720 342.970 2496.010 ;
        RECT 343.810 2495.720 354.930 2496.010 ;
        RECT 355.770 2495.720 367.810 2496.010 ;
        RECT 368.650 2495.720 379.770 2496.010 ;
        RECT 380.610 2495.720 391.730 2496.010 ;
        RECT 392.570 2495.720 404.610 2496.010 ;
        RECT 405.450 2495.720 416.570 2496.010 ;
        RECT 417.410 2495.720 429.450 2496.010 ;
        RECT 430.290 2495.720 441.410 2496.010 ;
        RECT 442.250 2495.720 454.290 2496.010 ;
        RECT 455.130 2495.720 466.250 2496.010 ;
        RECT 467.090 2495.720 478.210 2496.010 ;
        RECT 479.050 2495.720 491.090 2496.010 ;
        RECT 491.930 2495.720 503.050 2496.010 ;
        RECT 503.890 2495.720 515.930 2496.010 ;
        RECT 516.770 2495.720 527.890 2496.010 ;
        RECT 528.730 2495.720 540.770 2496.010 ;
        RECT 541.610 2495.720 552.730 2496.010 ;
        RECT 553.570 2495.720 564.690 2496.010 ;
        RECT 565.530 2495.720 577.570 2496.010 ;
        RECT 578.410 2495.720 589.530 2496.010 ;
        RECT 590.370 2495.720 602.410 2496.010 ;
        RECT 603.250 2495.720 614.370 2496.010 ;
        RECT 615.210 2495.720 627.250 2496.010 ;
        RECT 628.090 2495.720 639.210 2496.010 ;
        RECT 640.050 2495.720 651.170 2496.010 ;
        RECT 652.010 2495.720 664.050 2496.010 ;
        RECT 664.890 2495.720 676.010 2496.010 ;
        RECT 676.850 2495.720 688.890 2496.010 ;
        RECT 689.730 2495.720 700.850 2496.010 ;
        RECT 701.690 2495.720 713.730 2496.010 ;
        RECT 714.570 2495.720 725.690 2496.010 ;
        RECT 726.530 2495.720 737.650 2496.010 ;
        RECT 738.490 2495.720 750.530 2496.010 ;
        RECT 751.370 2495.720 762.490 2496.010 ;
        RECT 763.330 2495.720 775.370 2496.010 ;
        RECT 776.210 2495.720 787.330 2496.010 ;
        RECT 788.170 2495.720 800.210 2496.010 ;
        RECT 801.050 2495.720 812.170 2496.010 ;
        RECT 813.010 2495.720 824.130 2496.010 ;
        RECT 824.970 2495.720 837.010 2496.010 ;
        RECT 837.850 2495.720 848.970 2496.010 ;
        RECT 849.810 2495.720 861.850 2496.010 ;
        RECT 862.690 2495.720 873.810 2496.010 ;
        RECT 874.650 2495.720 886.690 2496.010 ;
        RECT 887.530 2495.720 898.650 2496.010 ;
        RECT 899.490 2495.720 910.610 2496.010 ;
        RECT 911.450 2495.720 923.490 2496.010 ;
        RECT 924.330 2495.720 935.450 2496.010 ;
        RECT 936.290 2495.720 948.330 2496.010 ;
        RECT 949.170 2495.720 960.290 2496.010 ;
        RECT 961.130 2495.720 973.170 2496.010 ;
        RECT 974.010 2495.720 985.130 2496.010 ;
        RECT 985.970 2495.720 997.090 2496.010 ;
        RECT 997.930 2495.720 1009.970 2496.010 ;
        RECT 1010.810 2495.720 1021.930 2496.010 ;
        RECT 1022.770 2495.720 1034.810 2496.010 ;
        RECT 1035.650 2495.720 1046.770 2496.010 ;
        RECT 1047.610 2495.720 1059.650 2496.010 ;
        RECT 1060.490 2495.720 1071.610 2496.010 ;
        RECT 1072.450 2495.720 1083.570 2496.010 ;
        RECT 1084.410 2495.720 1096.450 2496.010 ;
        RECT 1097.290 2495.720 1108.410 2496.010 ;
        RECT 1109.250 2495.720 1121.290 2496.010 ;
        RECT 1122.130 2495.720 1133.250 2496.010 ;
        RECT 1134.090 2495.720 1146.130 2496.010 ;
        RECT 1146.970 2495.720 1158.090 2496.010 ;
        RECT 1158.930 2495.720 1170.050 2496.010 ;
        RECT 1170.890 2495.720 1182.930 2496.010 ;
        RECT 1183.770 2495.720 1194.890 2496.010 ;
        RECT 1195.730 2495.720 1207.770 2496.010 ;
        RECT 1208.610 2495.720 1219.730 2496.010 ;
        RECT 1220.570 2495.720 1232.610 2496.010 ;
        RECT 1233.450 2495.720 1244.570 2496.010 ;
        RECT 1245.410 2495.720 1256.530 2496.010 ;
        RECT 1257.370 2495.720 1269.410 2496.010 ;
        RECT 1270.250 2495.720 1281.370 2496.010 ;
        RECT 1282.210 2495.720 1294.250 2496.010 ;
        RECT 1295.090 2495.720 1306.210 2496.010 ;
        RECT 1307.050 2495.720 1319.090 2496.010 ;
        RECT 1319.930 2495.720 1331.050 2496.010 ;
        RECT 1331.890 2495.720 1343.010 2496.010 ;
        RECT 1343.850 2495.720 1355.890 2496.010 ;
        RECT 1356.730 2495.720 1367.850 2496.010 ;
        RECT 1368.690 2495.720 1380.730 2496.010 ;
        RECT 1381.570 2495.720 1392.690 2496.010 ;
        RECT 1393.530 2495.720 1405.570 2496.010 ;
        RECT 1406.410 2495.720 1417.530 2496.010 ;
        RECT 1418.370 2495.720 1429.490 2496.010 ;
        RECT 1430.330 2495.720 1442.370 2496.010 ;
        RECT 1443.210 2495.720 1454.330 2496.010 ;
        RECT 1455.170 2495.720 1467.210 2496.010 ;
        RECT 1468.050 2495.720 1479.170 2496.010 ;
        RECT 1480.010 2495.720 1492.050 2496.010 ;
        RECT 1492.890 2495.720 1504.010 2496.010 ;
        RECT 1504.850 2495.720 1515.970 2496.010 ;
        RECT 1516.810 2495.720 1528.850 2496.010 ;
        RECT 1529.690 2495.720 1540.810 2496.010 ;
        RECT 1541.650 2495.720 1553.690 2496.010 ;
        RECT 1554.530 2495.720 1565.650 2496.010 ;
        RECT 1566.490 2495.720 1578.530 2496.010 ;
        RECT 1579.370 2495.720 1590.490 2496.010 ;
        RECT 1591.330 2495.720 1602.450 2496.010 ;
        RECT 1603.290 2495.720 1615.330 2496.010 ;
        RECT 1616.170 2495.720 1627.290 2496.010 ;
        RECT 1628.130 2495.720 1640.170 2496.010 ;
        RECT 1641.010 2495.720 1652.130 2496.010 ;
        RECT 1652.970 2495.720 1665.010 2496.010 ;
        RECT 1665.850 2495.720 1676.970 2496.010 ;
        RECT 1677.810 2495.720 1688.930 2496.010 ;
        RECT 1689.770 2495.720 1701.810 2496.010 ;
        RECT 1702.650 2495.720 1713.770 2496.010 ;
        RECT 1714.610 2495.720 1726.650 2496.010 ;
        RECT 1727.490 2495.720 1738.610 2496.010 ;
        RECT 1739.450 2495.720 1751.490 2496.010 ;
        RECT 1752.330 2495.720 1763.450 2496.010 ;
        RECT 1764.290 2495.720 1775.410 2496.010 ;
        RECT 1776.250 2495.720 1788.290 2496.010 ;
        RECT 1789.130 2495.720 1800.250 2496.010 ;
        RECT 1801.090 2495.720 1813.130 2496.010 ;
        RECT 1813.970 2495.720 1825.090 2496.010 ;
        RECT 1825.930 2495.720 1837.970 2496.010 ;
        RECT 1838.810 2495.720 1849.930 2496.010 ;
        RECT 1850.770 2495.720 1861.890 2496.010 ;
        RECT 1862.730 2495.720 1874.770 2496.010 ;
        RECT 1875.610 2495.720 1886.730 2496.010 ;
        RECT 1887.570 2495.720 1899.610 2496.010 ;
        RECT 1900.450 2495.720 1911.570 2496.010 ;
        RECT 1912.410 2495.720 1924.450 2496.010 ;
        RECT 1925.290 2495.720 1936.410 2496.010 ;
        RECT 1937.250 2495.720 1948.370 2496.010 ;
        RECT 1949.210 2495.720 1961.250 2496.010 ;
        RECT 1962.090 2495.720 1973.210 2496.010 ;
        RECT 1974.050 2495.720 1986.090 2496.010 ;
        RECT 1986.930 2495.720 1998.050 2496.010 ;
        RECT 1998.890 2495.720 2010.930 2496.010 ;
        RECT 2011.770 2495.720 2022.890 2496.010 ;
        RECT 2023.730 2495.720 2034.850 2496.010 ;
        RECT 2035.690 2495.720 2047.730 2496.010 ;
        RECT 2048.570 2495.720 2059.690 2496.010 ;
        RECT 2060.530 2495.720 2072.570 2496.010 ;
        RECT 2073.410 2495.720 2084.530 2496.010 ;
        RECT 2085.370 2495.720 2096.490 2496.010 ;
        RECT 8.840 4.280 2097.040 2495.720 ;
        RECT 8.840 4.000 14.530 4.280 ;
        RECT 15.370 4.000 26.490 4.280 ;
        RECT 27.330 4.000 39.370 4.280 ;
        RECT 40.210 4.000 51.330 4.280 ;
        RECT 52.170 4.000 64.210 4.280 ;
        RECT 65.050 4.000 76.170 4.280 ;
        RECT 77.010 4.000 88.130 4.280 ;
        RECT 88.970 4.000 101.010 4.280 ;
        RECT 101.850 4.000 112.970 4.280 ;
        RECT 113.810 4.000 125.850 4.280 ;
        RECT 126.690 4.000 137.810 4.280 ;
        RECT 138.650 4.000 150.690 4.280 ;
        RECT 151.530 4.000 162.650 4.280 ;
        RECT 163.490 4.000 174.610 4.280 ;
        RECT 175.450 4.000 187.490 4.280 ;
        RECT 188.330 4.000 199.450 4.280 ;
        RECT 200.290 4.000 212.330 4.280 ;
        RECT 213.170 4.000 224.290 4.280 ;
        RECT 225.130 4.000 237.170 4.280 ;
        RECT 238.010 4.000 249.130 4.280 ;
        RECT 249.970 4.000 261.090 4.280 ;
        RECT 261.930 4.000 273.970 4.280 ;
        RECT 274.810 4.000 285.930 4.280 ;
        RECT 286.770 4.000 298.810 4.280 ;
        RECT 299.650 4.000 310.770 4.280 ;
        RECT 311.610 4.000 323.650 4.280 ;
        RECT 324.490 4.000 335.610 4.280 ;
        RECT 336.450 4.000 347.570 4.280 ;
        RECT 348.410 4.000 360.450 4.280 ;
        RECT 361.290 4.000 372.410 4.280 ;
        RECT 373.250 4.000 385.290 4.280 ;
        RECT 386.130 4.000 397.250 4.280 ;
        RECT 398.090 4.000 410.130 4.280 ;
        RECT 410.970 4.000 422.090 4.280 ;
        RECT 422.930 4.000 434.050 4.280 ;
        RECT 434.890 4.000 446.930 4.280 ;
        RECT 447.770 4.000 458.890 4.280 ;
        RECT 459.730 4.000 471.770 4.280 ;
        RECT 472.610 4.000 483.730 4.280 ;
        RECT 484.570 4.000 496.610 4.280 ;
        RECT 497.450 4.000 508.570 4.280 ;
        RECT 509.410 4.000 520.530 4.280 ;
        RECT 521.370 4.000 533.410 4.280 ;
        RECT 534.250 4.000 545.370 4.280 ;
        RECT 546.210 4.000 558.250 4.280 ;
        RECT 559.090 4.000 570.210 4.280 ;
        RECT 571.050 4.000 583.090 4.280 ;
        RECT 583.930 4.000 595.050 4.280 ;
        RECT 595.890 4.000 607.010 4.280 ;
        RECT 607.850 4.000 619.890 4.280 ;
        RECT 620.730 4.000 631.850 4.280 ;
        RECT 632.690 4.000 644.730 4.280 ;
        RECT 645.570 4.000 656.690 4.280 ;
        RECT 657.530 4.000 669.570 4.280 ;
        RECT 670.410 4.000 681.530 4.280 ;
        RECT 682.370 4.000 693.490 4.280 ;
        RECT 694.330 4.000 706.370 4.280 ;
        RECT 707.210 4.000 718.330 4.280 ;
        RECT 719.170 4.000 731.210 4.280 ;
        RECT 732.050 4.000 743.170 4.280 ;
        RECT 744.010 4.000 756.050 4.280 ;
        RECT 756.890 4.000 768.010 4.280 ;
        RECT 768.850 4.000 779.970 4.280 ;
        RECT 780.810 4.000 792.850 4.280 ;
        RECT 793.690 4.000 804.810 4.280 ;
        RECT 805.650 4.000 817.690 4.280 ;
        RECT 818.530 4.000 829.650 4.280 ;
        RECT 830.490 4.000 842.530 4.280 ;
        RECT 843.370 4.000 854.490 4.280 ;
        RECT 855.330 4.000 866.450 4.280 ;
        RECT 867.290 4.000 879.330 4.280 ;
        RECT 880.170 4.000 891.290 4.280 ;
        RECT 892.130 4.000 904.170 4.280 ;
        RECT 905.010 4.000 916.130 4.280 ;
        RECT 916.970 4.000 929.010 4.280 ;
        RECT 929.850 4.000 940.970 4.280 ;
        RECT 941.810 4.000 952.930 4.280 ;
        RECT 953.770 4.000 965.810 4.280 ;
        RECT 966.650 4.000 977.770 4.280 ;
        RECT 978.610 4.000 990.650 4.280 ;
        RECT 991.490 4.000 1002.610 4.280 ;
        RECT 1003.450 4.000 1015.490 4.280 ;
        RECT 1016.330 4.000 1027.450 4.280 ;
        RECT 1028.290 4.000 1039.410 4.280 ;
        RECT 1040.250 4.000 1052.290 4.280 ;
        RECT 1053.130 4.000 1064.250 4.280 ;
        RECT 1065.090 4.000 1077.130 4.280 ;
        RECT 1077.970 4.000 1089.090 4.280 ;
        RECT 1089.930 4.000 1101.970 4.280 ;
        RECT 1102.810 4.000 1113.930 4.280 ;
        RECT 1114.770 4.000 1125.890 4.280 ;
        RECT 1126.730 4.000 1138.770 4.280 ;
        RECT 1139.610 4.000 1150.730 4.280 ;
        RECT 1151.570 4.000 1163.610 4.280 ;
        RECT 1164.450 4.000 1175.570 4.280 ;
        RECT 1176.410 4.000 1188.450 4.280 ;
        RECT 1189.290 4.000 1200.410 4.280 ;
        RECT 1201.250 4.000 1212.370 4.280 ;
        RECT 1213.210 4.000 1225.250 4.280 ;
        RECT 1226.090 4.000 1237.210 4.280 ;
        RECT 1238.050 4.000 1250.090 4.280 ;
        RECT 1250.930 4.000 1262.050 4.280 ;
        RECT 1262.890 4.000 1274.930 4.280 ;
        RECT 1275.770 4.000 1286.890 4.280 ;
        RECT 1287.730 4.000 1298.850 4.280 ;
        RECT 1299.690 4.000 1311.730 4.280 ;
        RECT 1312.570 4.000 1323.690 4.280 ;
        RECT 1324.530 4.000 1336.570 4.280 ;
        RECT 1337.410 4.000 1348.530 4.280 ;
        RECT 1349.370 4.000 1361.410 4.280 ;
        RECT 1362.250 4.000 1373.370 4.280 ;
        RECT 1374.210 4.000 1385.330 4.280 ;
        RECT 1386.170 4.000 1398.210 4.280 ;
        RECT 1399.050 4.000 1410.170 4.280 ;
        RECT 1411.010 4.000 1423.050 4.280 ;
        RECT 1423.890 4.000 1435.010 4.280 ;
        RECT 1435.850 4.000 1447.890 4.280 ;
        RECT 1448.730 4.000 1459.850 4.280 ;
        RECT 1460.690 4.000 1471.810 4.280 ;
        RECT 1472.650 4.000 1484.690 4.280 ;
        RECT 1485.530 4.000 1496.650 4.280 ;
        RECT 1497.490 4.000 1509.530 4.280 ;
        RECT 1510.370 4.000 1521.490 4.280 ;
        RECT 1522.330 4.000 1534.370 4.280 ;
        RECT 1535.210 4.000 1546.330 4.280 ;
        RECT 1547.170 4.000 1558.290 4.280 ;
        RECT 1559.130 4.000 1571.170 4.280 ;
        RECT 1572.010 4.000 1583.130 4.280 ;
        RECT 1583.970 4.000 1596.010 4.280 ;
        RECT 1596.850 4.000 1607.970 4.280 ;
        RECT 1608.810 4.000 1620.850 4.280 ;
        RECT 1621.690 4.000 1632.810 4.280 ;
        RECT 1633.650 4.000 1644.770 4.280 ;
        RECT 1645.610 4.000 1657.650 4.280 ;
        RECT 1658.490 4.000 1669.610 4.280 ;
        RECT 1670.450 4.000 1682.490 4.280 ;
        RECT 1683.330 4.000 1694.450 4.280 ;
        RECT 1695.290 4.000 1707.330 4.280 ;
        RECT 1708.170 4.000 1719.290 4.280 ;
        RECT 1720.130 4.000 1731.250 4.280 ;
        RECT 1732.090 4.000 1744.130 4.280 ;
        RECT 1744.970 4.000 1756.090 4.280 ;
        RECT 1756.930 4.000 1768.970 4.280 ;
        RECT 1769.810 4.000 1780.930 4.280 ;
        RECT 1781.770 4.000 1793.810 4.280 ;
        RECT 1794.650 4.000 1805.770 4.280 ;
        RECT 1806.610 4.000 1817.730 4.280 ;
        RECT 1818.570 4.000 1830.610 4.280 ;
        RECT 1831.450 4.000 1842.570 4.280 ;
        RECT 1843.410 4.000 1855.450 4.280 ;
        RECT 1856.290 4.000 1867.410 4.280 ;
        RECT 1868.250 4.000 1880.290 4.280 ;
        RECT 1881.130 4.000 1892.250 4.280 ;
        RECT 1893.090 4.000 1904.210 4.280 ;
        RECT 1905.050 4.000 1917.090 4.280 ;
        RECT 1917.930 4.000 1929.050 4.280 ;
        RECT 1929.890 4.000 1941.930 4.280 ;
        RECT 1942.770 4.000 1953.890 4.280 ;
        RECT 1954.730 4.000 1966.770 4.280 ;
        RECT 1967.610 4.000 1978.730 4.280 ;
        RECT 1979.570 4.000 1990.690 4.280 ;
        RECT 1991.530 4.000 2003.570 4.280 ;
        RECT 2004.410 4.000 2015.530 4.280 ;
        RECT 2016.370 4.000 2028.410 4.280 ;
        RECT 2029.250 4.000 2040.370 4.280 ;
        RECT 2041.210 4.000 2053.250 4.280 ;
        RECT 2054.090 4.000 2065.210 4.280 ;
        RECT 2066.050 4.000 2077.170 4.280 ;
        RECT 2078.010 4.000 2090.050 4.280 ;
        RECT 2090.890 4.000 2097.040 4.280 ;
      LAYER met3 ;
        RECT 4.000 2488.480 2096.000 2488.965 ;
        RECT 4.400 2487.080 2096.000 2488.480 ;
        RECT 4.000 2477.600 2096.000 2487.080 ;
        RECT 4.000 2476.200 2095.600 2477.600 ;
        RECT 4.000 2469.440 2096.000 2476.200 ;
        RECT 4.400 2468.040 2096.000 2469.440 ;
        RECT 4.000 2459.920 2096.000 2468.040 ;
        RECT 4.000 2458.520 2095.600 2459.920 ;
        RECT 4.000 2451.760 2096.000 2458.520 ;
        RECT 4.400 2450.360 2096.000 2451.760 ;
        RECT 4.000 2440.880 2096.000 2450.360 ;
        RECT 4.000 2439.480 2095.600 2440.880 ;
        RECT 4.000 2432.720 2096.000 2439.480 ;
        RECT 4.400 2431.320 2096.000 2432.720 ;
        RECT 4.000 2423.200 2096.000 2431.320 ;
        RECT 4.000 2421.800 2095.600 2423.200 ;
        RECT 4.000 2415.040 2096.000 2421.800 ;
        RECT 4.400 2413.640 2096.000 2415.040 ;
        RECT 4.000 2404.160 2096.000 2413.640 ;
        RECT 4.000 2402.760 2095.600 2404.160 ;
        RECT 4.000 2397.360 2096.000 2402.760 ;
        RECT 4.400 2395.960 2096.000 2397.360 ;
        RECT 4.000 2386.480 2096.000 2395.960 ;
        RECT 4.000 2385.080 2095.600 2386.480 ;
        RECT 4.000 2378.320 2096.000 2385.080 ;
        RECT 4.400 2376.920 2096.000 2378.320 ;
        RECT 4.000 2368.800 2096.000 2376.920 ;
        RECT 4.000 2367.400 2095.600 2368.800 ;
        RECT 4.000 2360.640 2096.000 2367.400 ;
        RECT 4.400 2359.240 2096.000 2360.640 ;
        RECT 4.000 2349.760 2096.000 2359.240 ;
        RECT 4.000 2348.360 2095.600 2349.760 ;
        RECT 4.000 2341.600 2096.000 2348.360 ;
        RECT 4.400 2340.200 2096.000 2341.600 ;
        RECT 4.000 2332.080 2096.000 2340.200 ;
        RECT 4.000 2330.680 2095.600 2332.080 ;
        RECT 4.000 2323.920 2096.000 2330.680 ;
        RECT 4.400 2322.520 2096.000 2323.920 ;
        RECT 4.000 2313.040 2096.000 2322.520 ;
        RECT 4.000 2311.640 2095.600 2313.040 ;
        RECT 4.000 2304.880 2096.000 2311.640 ;
        RECT 4.400 2303.480 2096.000 2304.880 ;
        RECT 4.000 2295.360 2096.000 2303.480 ;
        RECT 4.000 2293.960 2095.600 2295.360 ;
        RECT 4.000 2287.200 2096.000 2293.960 ;
        RECT 4.400 2285.800 2096.000 2287.200 ;
        RECT 4.000 2276.320 2096.000 2285.800 ;
        RECT 4.000 2274.920 2095.600 2276.320 ;
        RECT 4.000 2269.520 2096.000 2274.920 ;
        RECT 4.400 2268.120 2096.000 2269.520 ;
        RECT 4.000 2258.640 2096.000 2268.120 ;
        RECT 4.000 2257.240 2095.600 2258.640 ;
        RECT 4.000 2250.480 2096.000 2257.240 ;
        RECT 4.400 2249.080 2096.000 2250.480 ;
        RECT 4.000 2240.960 2096.000 2249.080 ;
        RECT 4.000 2239.560 2095.600 2240.960 ;
        RECT 4.000 2232.800 2096.000 2239.560 ;
        RECT 4.400 2231.400 2096.000 2232.800 ;
        RECT 4.000 2221.920 2096.000 2231.400 ;
        RECT 4.000 2220.520 2095.600 2221.920 ;
        RECT 4.000 2213.760 2096.000 2220.520 ;
        RECT 4.400 2212.360 2096.000 2213.760 ;
        RECT 4.000 2204.240 2096.000 2212.360 ;
        RECT 4.000 2202.840 2095.600 2204.240 ;
        RECT 4.000 2196.080 2096.000 2202.840 ;
        RECT 4.400 2194.680 2096.000 2196.080 ;
        RECT 4.000 2185.200 2096.000 2194.680 ;
        RECT 4.000 2183.800 2095.600 2185.200 ;
        RECT 4.000 2177.040 2096.000 2183.800 ;
        RECT 4.400 2175.640 2096.000 2177.040 ;
        RECT 4.000 2167.520 2096.000 2175.640 ;
        RECT 4.000 2166.120 2095.600 2167.520 ;
        RECT 4.000 2159.360 2096.000 2166.120 ;
        RECT 4.400 2157.960 2096.000 2159.360 ;
        RECT 4.000 2148.480 2096.000 2157.960 ;
        RECT 4.000 2147.080 2095.600 2148.480 ;
        RECT 4.000 2141.680 2096.000 2147.080 ;
        RECT 4.400 2140.280 2096.000 2141.680 ;
        RECT 4.000 2130.800 2096.000 2140.280 ;
        RECT 4.000 2129.400 2095.600 2130.800 ;
        RECT 4.000 2122.640 2096.000 2129.400 ;
        RECT 4.400 2121.240 2096.000 2122.640 ;
        RECT 4.000 2113.120 2096.000 2121.240 ;
        RECT 4.000 2111.720 2095.600 2113.120 ;
        RECT 4.000 2104.960 2096.000 2111.720 ;
        RECT 4.400 2103.560 2096.000 2104.960 ;
        RECT 4.000 2094.080 2096.000 2103.560 ;
        RECT 4.000 2092.680 2095.600 2094.080 ;
        RECT 4.000 2085.920 2096.000 2092.680 ;
        RECT 4.400 2084.520 2096.000 2085.920 ;
        RECT 4.000 2076.400 2096.000 2084.520 ;
        RECT 4.000 2075.000 2095.600 2076.400 ;
        RECT 4.000 2068.240 2096.000 2075.000 ;
        RECT 4.400 2066.840 2096.000 2068.240 ;
        RECT 4.000 2057.360 2096.000 2066.840 ;
        RECT 4.000 2055.960 2095.600 2057.360 ;
        RECT 4.000 2049.200 2096.000 2055.960 ;
        RECT 4.400 2047.800 2096.000 2049.200 ;
        RECT 4.000 2039.680 2096.000 2047.800 ;
        RECT 4.000 2038.280 2095.600 2039.680 ;
        RECT 4.000 2031.520 2096.000 2038.280 ;
        RECT 4.400 2030.120 2096.000 2031.520 ;
        RECT 4.000 2020.640 2096.000 2030.120 ;
        RECT 4.000 2019.240 2095.600 2020.640 ;
        RECT 4.000 2013.840 2096.000 2019.240 ;
        RECT 4.400 2012.440 2096.000 2013.840 ;
        RECT 4.000 2002.960 2096.000 2012.440 ;
        RECT 4.000 2001.560 2095.600 2002.960 ;
        RECT 4.000 1994.800 2096.000 2001.560 ;
        RECT 4.400 1993.400 2096.000 1994.800 ;
        RECT 4.000 1985.280 2096.000 1993.400 ;
        RECT 4.000 1983.880 2095.600 1985.280 ;
        RECT 4.000 1977.120 2096.000 1983.880 ;
        RECT 4.400 1975.720 2096.000 1977.120 ;
        RECT 4.000 1966.240 2096.000 1975.720 ;
        RECT 4.000 1964.840 2095.600 1966.240 ;
        RECT 4.000 1958.080 2096.000 1964.840 ;
        RECT 4.400 1956.680 2096.000 1958.080 ;
        RECT 4.000 1948.560 2096.000 1956.680 ;
        RECT 4.000 1947.160 2095.600 1948.560 ;
        RECT 4.000 1940.400 2096.000 1947.160 ;
        RECT 4.400 1939.000 2096.000 1940.400 ;
        RECT 4.000 1929.520 2096.000 1939.000 ;
        RECT 4.000 1928.120 2095.600 1929.520 ;
        RECT 4.000 1921.360 2096.000 1928.120 ;
        RECT 4.400 1919.960 2096.000 1921.360 ;
        RECT 4.000 1911.840 2096.000 1919.960 ;
        RECT 4.000 1910.440 2095.600 1911.840 ;
        RECT 4.000 1903.680 2096.000 1910.440 ;
        RECT 4.400 1902.280 2096.000 1903.680 ;
        RECT 4.000 1892.800 2096.000 1902.280 ;
        RECT 4.000 1891.400 2095.600 1892.800 ;
        RECT 4.000 1886.000 2096.000 1891.400 ;
        RECT 4.400 1884.600 2096.000 1886.000 ;
        RECT 4.000 1875.120 2096.000 1884.600 ;
        RECT 4.000 1873.720 2095.600 1875.120 ;
        RECT 4.000 1866.960 2096.000 1873.720 ;
        RECT 4.400 1865.560 2096.000 1866.960 ;
        RECT 4.000 1857.440 2096.000 1865.560 ;
        RECT 4.000 1856.040 2095.600 1857.440 ;
        RECT 4.000 1849.280 2096.000 1856.040 ;
        RECT 4.400 1847.880 2096.000 1849.280 ;
        RECT 4.000 1838.400 2096.000 1847.880 ;
        RECT 4.000 1837.000 2095.600 1838.400 ;
        RECT 4.000 1830.240 2096.000 1837.000 ;
        RECT 4.400 1828.840 2096.000 1830.240 ;
        RECT 4.000 1820.720 2096.000 1828.840 ;
        RECT 4.000 1819.320 2095.600 1820.720 ;
        RECT 4.000 1812.560 2096.000 1819.320 ;
        RECT 4.400 1811.160 2096.000 1812.560 ;
        RECT 4.000 1801.680 2096.000 1811.160 ;
        RECT 4.000 1800.280 2095.600 1801.680 ;
        RECT 4.000 1793.520 2096.000 1800.280 ;
        RECT 4.400 1792.120 2096.000 1793.520 ;
        RECT 4.000 1784.000 2096.000 1792.120 ;
        RECT 4.000 1782.600 2095.600 1784.000 ;
        RECT 4.000 1775.840 2096.000 1782.600 ;
        RECT 4.400 1774.440 2096.000 1775.840 ;
        RECT 4.000 1764.960 2096.000 1774.440 ;
        RECT 4.000 1763.560 2095.600 1764.960 ;
        RECT 4.000 1758.160 2096.000 1763.560 ;
        RECT 4.400 1756.760 2096.000 1758.160 ;
        RECT 4.000 1747.280 2096.000 1756.760 ;
        RECT 4.000 1745.880 2095.600 1747.280 ;
        RECT 4.000 1739.120 2096.000 1745.880 ;
        RECT 4.400 1737.720 2096.000 1739.120 ;
        RECT 4.000 1729.600 2096.000 1737.720 ;
        RECT 4.000 1728.200 2095.600 1729.600 ;
        RECT 4.000 1721.440 2096.000 1728.200 ;
        RECT 4.400 1720.040 2096.000 1721.440 ;
        RECT 4.000 1710.560 2096.000 1720.040 ;
        RECT 4.000 1709.160 2095.600 1710.560 ;
        RECT 4.000 1702.400 2096.000 1709.160 ;
        RECT 4.400 1701.000 2096.000 1702.400 ;
        RECT 4.000 1692.880 2096.000 1701.000 ;
        RECT 4.000 1691.480 2095.600 1692.880 ;
        RECT 4.000 1684.720 2096.000 1691.480 ;
        RECT 4.400 1683.320 2096.000 1684.720 ;
        RECT 4.000 1673.840 2096.000 1683.320 ;
        RECT 4.000 1672.440 2095.600 1673.840 ;
        RECT 4.000 1665.680 2096.000 1672.440 ;
        RECT 4.400 1664.280 2096.000 1665.680 ;
        RECT 4.000 1656.160 2096.000 1664.280 ;
        RECT 4.000 1654.760 2095.600 1656.160 ;
        RECT 4.000 1648.000 2096.000 1654.760 ;
        RECT 4.400 1646.600 2096.000 1648.000 ;
        RECT 4.000 1637.120 2096.000 1646.600 ;
        RECT 4.000 1635.720 2095.600 1637.120 ;
        RECT 4.000 1630.320 2096.000 1635.720 ;
        RECT 4.400 1628.920 2096.000 1630.320 ;
        RECT 4.000 1619.440 2096.000 1628.920 ;
        RECT 4.000 1618.040 2095.600 1619.440 ;
        RECT 4.000 1611.280 2096.000 1618.040 ;
        RECT 4.400 1609.880 2096.000 1611.280 ;
        RECT 4.000 1601.760 2096.000 1609.880 ;
        RECT 4.000 1600.360 2095.600 1601.760 ;
        RECT 4.000 1593.600 2096.000 1600.360 ;
        RECT 4.400 1592.200 2096.000 1593.600 ;
        RECT 4.000 1582.720 2096.000 1592.200 ;
        RECT 4.000 1581.320 2095.600 1582.720 ;
        RECT 4.000 1574.560 2096.000 1581.320 ;
        RECT 4.400 1573.160 2096.000 1574.560 ;
        RECT 4.000 1565.040 2096.000 1573.160 ;
        RECT 4.000 1563.640 2095.600 1565.040 ;
        RECT 4.000 1556.880 2096.000 1563.640 ;
        RECT 4.400 1555.480 2096.000 1556.880 ;
        RECT 4.000 1546.000 2096.000 1555.480 ;
        RECT 4.000 1544.600 2095.600 1546.000 ;
        RECT 4.000 1537.840 2096.000 1544.600 ;
        RECT 4.400 1536.440 2096.000 1537.840 ;
        RECT 4.000 1528.320 2096.000 1536.440 ;
        RECT 4.000 1526.920 2095.600 1528.320 ;
        RECT 4.000 1520.160 2096.000 1526.920 ;
        RECT 4.400 1518.760 2096.000 1520.160 ;
        RECT 4.000 1509.280 2096.000 1518.760 ;
        RECT 4.000 1507.880 2095.600 1509.280 ;
        RECT 4.000 1502.480 2096.000 1507.880 ;
        RECT 4.400 1501.080 2096.000 1502.480 ;
        RECT 4.000 1491.600 2096.000 1501.080 ;
        RECT 4.000 1490.200 2095.600 1491.600 ;
        RECT 4.000 1483.440 2096.000 1490.200 ;
        RECT 4.400 1482.040 2096.000 1483.440 ;
        RECT 4.000 1473.920 2096.000 1482.040 ;
        RECT 4.000 1472.520 2095.600 1473.920 ;
        RECT 4.000 1465.760 2096.000 1472.520 ;
        RECT 4.400 1464.360 2096.000 1465.760 ;
        RECT 4.000 1454.880 2096.000 1464.360 ;
        RECT 4.000 1453.480 2095.600 1454.880 ;
        RECT 4.000 1446.720 2096.000 1453.480 ;
        RECT 4.400 1445.320 2096.000 1446.720 ;
        RECT 4.000 1437.200 2096.000 1445.320 ;
        RECT 4.000 1435.800 2095.600 1437.200 ;
        RECT 4.000 1429.040 2096.000 1435.800 ;
        RECT 4.400 1427.640 2096.000 1429.040 ;
        RECT 4.000 1418.160 2096.000 1427.640 ;
        RECT 4.000 1416.760 2095.600 1418.160 ;
        RECT 4.000 1410.000 2096.000 1416.760 ;
        RECT 4.400 1408.600 2096.000 1410.000 ;
        RECT 4.000 1400.480 2096.000 1408.600 ;
        RECT 4.000 1399.080 2095.600 1400.480 ;
        RECT 4.000 1392.320 2096.000 1399.080 ;
        RECT 4.400 1390.920 2096.000 1392.320 ;
        RECT 4.000 1381.440 2096.000 1390.920 ;
        RECT 4.000 1380.040 2095.600 1381.440 ;
        RECT 4.000 1374.640 2096.000 1380.040 ;
        RECT 4.400 1373.240 2096.000 1374.640 ;
        RECT 4.000 1363.760 2096.000 1373.240 ;
        RECT 4.000 1362.360 2095.600 1363.760 ;
        RECT 4.000 1355.600 2096.000 1362.360 ;
        RECT 4.400 1354.200 2096.000 1355.600 ;
        RECT 4.000 1346.080 2096.000 1354.200 ;
        RECT 4.000 1344.680 2095.600 1346.080 ;
        RECT 4.000 1337.920 2096.000 1344.680 ;
        RECT 4.400 1336.520 2096.000 1337.920 ;
        RECT 4.000 1327.040 2096.000 1336.520 ;
        RECT 4.000 1325.640 2095.600 1327.040 ;
        RECT 4.000 1318.880 2096.000 1325.640 ;
        RECT 4.400 1317.480 2096.000 1318.880 ;
        RECT 4.000 1309.360 2096.000 1317.480 ;
        RECT 4.000 1307.960 2095.600 1309.360 ;
        RECT 4.000 1301.200 2096.000 1307.960 ;
        RECT 4.400 1299.800 2096.000 1301.200 ;
        RECT 4.000 1290.320 2096.000 1299.800 ;
        RECT 4.000 1288.920 2095.600 1290.320 ;
        RECT 4.000 1282.160 2096.000 1288.920 ;
        RECT 4.400 1280.760 2096.000 1282.160 ;
        RECT 4.000 1272.640 2096.000 1280.760 ;
        RECT 4.000 1271.240 2095.600 1272.640 ;
        RECT 4.000 1264.480 2096.000 1271.240 ;
        RECT 4.400 1263.080 2096.000 1264.480 ;
        RECT 4.000 1253.600 2096.000 1263.080 ;
        RECT 4.000 1252.200 2095.600 1253.600 ;
        RECT 4.000 1246.800 2096.000 1252.200 ;
        RECT 4.400 1245.400 2096.000 1246.800 ;
        RECT 4.000 1235.920 2096.000 1245.400 ;
        RECT 4.000 1234.520 2095.600 1235.920 ;
        RECT 4.000 1227.760 2096.000 1234.520 ;
        RECT 4.400 1226.360 2096.000 1227.760 ;
        RECT 4.000 1218.240 2096.000 1226.360 ;
        RECT 4.000 1216.840 2095.600 1218.240 ;
        RECT 4.000 1210.080 2096.000 1216.840 ;
        RECT 4.400 1208.680 2096.000 1210.080 ;
        RECT 4.000 1199.200 2096.000 1208.680 ;
        RECT 4.000 1197.800 2095.600 1199.200 ;
        RECT 4.000 1191.040 2096.000 1197.800 ;
        RECT 4.400 1189.640 2096.000 1191.040 ;
        RECT 4.000 1181.520 2096.000 1189.640 ;
        RECT 4.000 1180.120 2095.600 1181.520 ;
        RECT 4.000 1173.360 2096.000 1180.120 ;
        RECT 4.400 1171.960 2096.000 1173.360 ;
        RECT 4.000 1162.480 2096.000 1171.960 ;
        RECT 4.000 1161.080 2095.600 1162.480 ;
        RECT 4.000 1154.320 2096.000 1161.080 ;
        RECT 4.400 1152.920 2096.000 1154.320 ;
        RECT 4.000 1144.800 2096.000 1152.920 ;
        RECT 4.000 1143.400 2095.600 1144.800 ;
        RECT 4.000 1136.640 2096.000 1143.400 ;
        RECT 4.400 1135.240 2096.000 1136.640 ;
        RECT 4.000 1125.760 2096.000 1135.240 ;
        RECT 4.000 1124.360 2095.600 1125.760 ;
        RECT 4.000 1118.960 2096.000 1124.360 ;
        RECT 4.400 1117.560 2096.000 1118.960 ;
        RECT 4.000 1108.080 2096.000 1117.560 ;
        RECT 4.000 1106.680 2095.600 1108.080 ;
        RECT 4.000 1099.920 2096.000 1106.680 ;
        RECT 4.400 1098.520 2096.000 1099.920 ;
        RECT 4.000 1090.400 2096.000 1098.520 ;
        RECT 4.000 1089.000 2095.600 1090.400 ;
        RECT 4.000 1082.240 2096.000 1089.000 ;
        RECT 4.400 1080.840 2096.000 1082.240 ;
        RECT 4.000 1071.360 2096.000 1080.840 ;
        RECT 4.000 1069.960 2095.600 1071.360 ;
        RECT 4.000 1063.200 2096.000 1069.960 ;
        RECT 4.400 1061.800 2096.000 1063.200 ;
        RECT 4.000 1053.680 2096.000 1061.800 ;
        RECT 4.000 1052.280 2095.600 1053.680 ;
        RECT 4.000 1045.520 2096.000 1052.280 ;
        RECT 4.400 1044.120 2096.000 1045.520 ;
        RECT 4.000 1034.640 2096.000 1044.120 ;
        RECT 4.000 1033.240 2095.600 1034.640 ;
        RECT 4.000 1026.480 2096.000 1033.240 ;
        RECT 4.400 1025.080 2096.000 1026.480 ;
        RECT 4.000 1016.960 2096.000 1025.080 ;
        RECT 4.000 1015.560 2095.600 1016.960 ;
        RECT 4.000 1008.800 2096.000 1015.560 ;
        RECT 4.400 1007.400 2096.000 1008.800 ;
        RECT 4.000 997.920 2096.000 1007.400 ;
        RECT 4.000 996.520 2095.600 997.920 ;
        RECT 4.000 991.120 2096.000 996.520 ;
        RECT 4.400 989.720 2096.000 991.120 ;
        RECT 4.000 980.240 2096.000 989.720 ;
        RECT 4.000 978.840 2095.600 980.240 ;
        RECT 4.000 972.080 2096.000 978.840 ;
        RECT 4.400 970.680 2096.000 972.080 ;
        RECT 4.000 962.560 2096.000 970.680 ;
        RECT 4.000 961.160 2095.600 962.560 ;
        RECT 4.000 954.400 2096.000 961.160 ;
        RECT 4.400 953.000 2096.000 954.400 ;
        RECT 4.000 943.520 2096.000 953.000 ;
        RECT 4.000 942.120 2095.600 943.520 ;
        RECT 4.000 935.360 2096.000 942.120 ;
        RECT 4.400 933.960 2096.000 935.360 ;
        RECT 4.000 925.840 2096.000 933.960 ;
        RECT 4.000 924.440 2095.600 925.840 ;
        RECT 4.000 917.680 2096.000 924.440 ;
        RECT 4.400 916.280 2096.000 917.680 ;
        RECT 4.000 906.800 2096.000 916.280 ;
        RECT 4.000 905.400 2095.600 906.800 ;
        RECT 4.000 898.640 2096.000 905.400 ;
        RECT 4.400 897.240 2096.000 898.640 ;
        RECT 4.000 889.120 2096.000 897.240 ;
        RECT 4.000 887.720 2095.600 889.120 ;
        RECT 4.000 880.960 2096.000 887.720 ;
        RECT 4.400 879.560 2096.000 880.960 ;
        RECT 4.000 870.080 2096.000 879.560 ;
        RECT 4.000 868.680 2095.600 870.080 ;
        RECT 4.000 863.280 2096.000 868.680 ;
        RECT 4.400 861.880 2096.000 863.280 ;
        RECT 4.000 852.400 2096.000 861.880 ;
        RECT 4.000 851.000 2095.600 852.400 ;
        RECT 4.000 844.240 2096.000 851.000 ;
        RECT 4.400 842.840 2096.000 844.240 ;
        RECT 4.000 834.720 2096.000 842.840 ;
        RECT 4.000 833.320 2095.600 834.720 ;
        RECT 4.000 826.560 2096.000 833.320 ;
        RECT 4.400 825.160 2096.000 826.560 ;
        RECT 4.000 815.680 2096.000 825.160 ;
        RECT 4.000 814.280 2095.600 815.680 ;
        RECT 4.000 807.520 2096.000 814.280 ;
        RECT 4.400 806.120 2096.000 807.520 ;
        RECT 4.000 798.000 2096.000 806.120 ;
        RECT 4.000 796.600 2095.600 798.000 ;
        RECT 4.000 789.840 2096.000 796.600 ;
        RECT 4.400 788.440 2096.000 789.840 ;
        RECT 4.000 778.960 2096.000 788.440 ;
        RECT 4.000 777.560 2095.600 778.960 ;
        RECT 4.000 770.800 2096.000 777.560 ;
        RECT 4.400 769.400 2096.000 770.800 ;
        RECT 4.000 761.280 2096.000 769.400 ;
        RECT 4.000 759.880 2095.600 761.280 ;
        RECT 4.000 753.120 2096.000 759.880 ;
        RECT 4.400 751.720 2096.000 753.120 ;
        RECT 4.000 742.240 2096.000 751.720 ;
        RECT 4.000 740.840 2095.600 742.240 ;
        RECT 4.000 735.440 2096.000 740.840 ;
        RECT 4.400 734.040 2096.000 735.440 ;
        RECT 4.000 724.560 2096.000 734.040 ;
        RECT 4.000 723.160 2095.600 724.560 ;
        RECT 4.000 716.400 2096.000 723.160 ;
        RECT 4.400 715.000 2096.000 716.400 ;
        RECT 4.000 706.880 2096.000 715.000 ;
        RECT 4.000 705.480 2095.600 706.880 ;
        RECT 4.000 698.720 2096.000 705.480 ;
        RECT 4.400 697.320 2096.000 698.720 ;
        RECT 4.000 687.840 2096.000 697.320 ;
        RECT 4.000 686.440 2095.600 687.840 ;
        RECT 4.000 679.680 2096.000 686.440 ;
        RECT 4.400 678.280 2096.000 679.680 ;
        RECT 4.000 670.160 2096.000 678.280 ;
        RECT 4.000 668.760 2095.600 670.160 ;
        RECT 4.000 662.000 2096.000 668.760 ;
        RECT 4.400 660.600 2096.000 662.000 ;
        RECT 4.000 651.120 2096.000 660.600 ;
        RECT 4.000 649.720 2095.600 651.120 ;
        RECT 4.000 642.960 2096.000 649.720 ;
        RECT 4.400 641.560 2096.000 642.960 ;
        RECT 4.000 633.440 2096.000 641.560 ;
        RECT 4.000 632.040 2095.600 633.440 ;
        RECT 4.000 625.280 2096.000 632.040 ;
        RECT 4.400 623.880 2096.000 625.280 ;
        RECT 4.000 614.400 2096.000 623.880 ;
        RECT 4.000 613.000 2095.600 614.400 ;
        RECT 4.000 607.600 2096.000 613.000 ;
        RECT 4.400 606.200 2096.000 607.600 ;
        RECT 4.000 596.720 2096.000 606.200 ;
        RECT 4.000 595.320 2095.600 596.720 ;
        RECT 4.000 588.560 2096.000 595.320 ;
        RECT 4.400 587.160 2096.000 588.560 ;
        RECT 4.000 579.040 2096.000 587.160 ;
        RECT 4.000 577.640 2095.600 579.040 ;
        RECT 4.000 570.880 2096.000 577.640 ;
        RECT 4.400 569.480 2096.000 570.880 ;
        RECT 4.000 560.000 2096.000 569.480 ;
        RECT 4.000 558.600 2095.600 560.000 ;
        RECT 4.000 551.840 2096.000 558.600 ;
        RECT 4.400 550.440 2096.000 551.840 ;
        RECT 4.000 542.320 2096.000 550.440 ;
        RECT 4.000 540.920 2095.600 542.320 ;
        RECT 4.000 534.160 2096.000 540.920 ;
        RECT 4.400 532.760 2096.000 534.160 ;
        RECT 4.000 523.280 2096.000 532.760 ;
        RECT 4.000 521.880 2095.600 523.280 ;
        RECT 4.000 515.120 2096.000 521.880 ;
        RECT 4.400 513.720 2096.000 515.120 ;
        RECT 4.000 505.600 2096.000 513.720 ;
        RECT 4.000 504.200 2095.600 505.600 ;
        RECT 4.000 497.440 2096.000 504.200 ;
        RECT 4.400 496.040 2096.000 497.440 ;
        RECT 4.000 486.560 2096.000 496.040 ;
        RECT 4.000 485.160 2095.600 486.560 ;
        RECT 4.000 479.760 2096.000 485.160 ;
        RECT 4.400 478.360 2096.000 479.760 ;
        RECT 4.000 468.880 2096.000 478.360 ;
        RECT 4.000 467.480 2095.600 468.880 ;
        RECT 4.000 460.720 2096.000 467.480 ;
        RECT 4.400 459.320 2096.000 460.720 ;
        RECT 4.000 451.200 2096.000 459.320 ;
        RECT 4.000 449.800 2095.600 451.200 ;
        RECT 4.000 443.040 2096.000 449.800 ;
        RECT 4.400 441.640 2096.000 443.040 ;
        RECT 4.000 432.160 2096.000 441.640 ;
        RECT 4.000 430.760 2095.600 432.160 ;
        RECT 4.000 424.000 2096.000 430.760 ;
        RECT 4.400 422.600 2096.000 424.000 ;
        RECT 4.000 414.480 2096.000 422.600 ;
        RECT 4.000 413.080 2095.600 414.480 ;
        RECT 4.000 406.320 2096.000 413.080 ;
        RECT 4.400 404.920 2096.000 406.320 ;
        RECT 4.000 395.440 2096.000 404.920 ;
        RECT 4.000 394.040 2095.600 395.440 ;
        RECT 4.000 387.280 2096.000 394.040 ;
        RECT 4.400 385.880 2096.000 387.280 ;
        RECT 4.000 377.760 2096.000 385.880 ;
        RECT 4.000 376.360 2095.600 377.760 ;
        RECT 4.000 369.600 2096.000 376.360 ;
        RECT 4.400 368.200 2096.000 369.600 ;
        RECT 4.000 358.720 2096.000 368.200 ;
        RECT 4.000 357.320 2095.600 358.720 ;
        RECT 4.000 351.920 2096.000 357.320 ;
        RECT 4.400 350.520 2096.000 351.920 ;
        RECT 4.000 341.040 2096.000 350.520 ;
        RECT 4.000 339.640 2095.600 341.040 ;
        RECT 4.000 332.880 2096.000 339.640 ;
        RECT 4.400 331.480 2096.000 332.880 ;
        RECT 4.000 323.360 2096.000 331.480 ;
        RECT 4.000 321.960 2095.600 323.360 ;
        RECT 4.000 315.200 2096.000 321.960 ;
        RECT 4.400 313.800 2096.000 315.200 ;
        RECT 4.000 304.320 2096.000 313.800 ;
        RECT 4.000 302.920 2095.600 304.320 ;
        RECT 4.000 296.160 2096.000 302.920 ;
        RECT 4.400 294.760 2096.000 296.160 ;
        RECT 4.000 286.640 2096.000 294.760 ;
        RECT 4.000 285.240 2095.600 286.640 ;
        RECT 4.000 278.480 2096.000 285.240 ;
        RECT 4.400 277.080 2096.000 278.480 ;
        RECT 4.000 267.600 2096.000 277.080 ;
        RECT 4.000 266.200 2095.600 267.600 ;
        RECT 4.000 259.440 2096.000 266.200 ;
        RECT 4.400 258.040 2096.000 259.440 ;
        RECT 4.000 249.920 2096.000 258.040 ;
        RECT 4.000 248.520 2095.600 249.920 ;
        RECT 4.000 241.760 2096.000 248.520 ;
        RECT 4.400 240.360 2096.000 241.760 ;
        RECT 4.000 230.880 2096.000 240.360 ;
        RECT 4.000 229.480 2095.600 230.880 ;
        RECT 4.000 224.080 2096.000 229.480 ;
        RECT 4.400 222.680 2096.000 224.080 ;
        RECT 4.000 213.200 2096.000 222.680 ;
        RECT 4.000 211.800 2095.600 213.200 ;
        RECT 4.000 205.040 2096.000 211.800 ;
        RECT 4.400 203.640 2096.000 205.040 ;
        RECT 4.000 195.520 2096.000 203.640 ;
        RECT 4.000 194.120 2095.600 195.520 ;
        RECT 4.000 187.360 2096.000 194.120 ;
        RECT 4.400 185.960 2096.000 187.360 ;
        RECT 4.000 176.480 2096.000 185.960 ;
        RECT 4.000 175.080 2095.600 176.480 ;
        RECT 4.000 168.320 2096.000 175.080 ;
        RECT 4.400 166.920 2096.000 168.320 ;
        RECT 4.000 158.800 2096.000 166.920 ;
        RECT 4.000 157.400 2095.600 158.800 ;
        RECT 4.000 150.640 2096.000 157.400 ;
        RECT 4.400 149.240 2096.000 150.640 ;
        RECT 4.000 139.760 2096.000 149.240 ;
        RECT 4.000 138.360 2095.600 139.760 ;
        RECT 4.000 131.600 2096.000 138.360 ;
        RECT 4.400 130.200 2096.000 131.600 ;
        RECT 4.000 122.080 2096.000 130.200 ;
        RECT 4.000 120.680 2095.600 122.080 ;
        RECT 4.000 113.920 2096.000 120.680 ;
        RECT 4.400 112.520 2096.000 113.920 ;
        RECT 4.000 103.040 2096.000 112.520 ;
        RECT 4.000 101.640 2095.600 103.040 ;
        RECT 4.000 96.240 2096.000 101.640 ;
        RECT 4.400 94.840 2096.000 96.240 ;
        RECT 4.000 85.360 2096.000 94.840 ;
        RECT 4.000 83.960 2095.600 85.360 ;
        RECT 4.000 77.200 2096.000 83.960 ;
        RECT 4.400 75.800 2096.000 77.200 ;
        RECT 4.000 67.680 2096.000 75.800 ;
        RECT 4.000 66.280 2095.600 67.680 ;
        RECT 4.000 59.520 2096.000 66.280 ;
        RECT 4.400 58.120 2096.000 59.520 ;
        RECT 4.000 48.640 2096.000 58.120 ;
        RECT 4.000 47.240 2095.600 48.640 ;
        RECT 4.000 40.480 2096.000 47.240 ;
        RECT 4.400 39.080 2096.000 40.480 ;
        RECT 4.000 30.960 2096.000 39.080 ;
        RECT 4.000 29.560 2095.600 30.960 ;
        RECT 4.000 22.800 2096.000 29.560 ;
        RECT 4.400 21.400 2096.000 22.800 ;
        RECT 4.000 11.920 2096.000 21.400 ;
        RECT 4.000 10.520 2095.600 11.920 ;
        RECT 4.000 4.255 2096.000 10.520 ;
      LAYER met4 ;
        RECT 12.255 10.640 20.640 2489.040 ;
        RECT 23.040 10.640 97.440 2489.040 ;
        RECT 99.840 10.640 2019.440 2489.040 ;
  END
END Ibtida_top_dffram_cv
END LIBRARY

