VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2528.690 89.660 2529.010 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2528.690 89.520 2899.310 89.660 ;
        RECT 2528.690 89.460 2529.010 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2528.720 89.460 2528.980 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2528.710 536.675 2528.990 537.045 ;
        RECT 2528.780 89.750 2528.920 536.675 ;
        RECT 2528.720 89.430 2528.980 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2528.710 536.720 2528.990 537.000 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2506.000 537.010 2510.000 537.160 ;
        RECT 2528.685 537.010 2529.015 537.025 ;
        RECT 2506.000 536.710 2529.015 537.010 ;
        RECT 2506.000 536.560 2510.000 536.710 ;
        RECT 2528.685 536.695 2529.015 536.710 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.090 2429.200 2570.410 2429.260 ;
        RECT 2899.450 2429.200 2899.770 2429.260 ;
        RECT 2570.090 2429.060 2899.770 2429.200 ;
        RECT 2570.090 2429.000 2570.410 2429.060 ;
        RECT 2899.450 2429.000 2899.770 2429.060 ;
        RECT 2523.170 2173.520 2523.490 2173.580 ;
        RECT 2570.090 2173.520 2570.410 2173.580 ;
        RECT 2523.170 2173.380 2570.410 2173.520 ;
        RECT 2523.170 2173.320 2523.490 2173.380 ;
        RECT 2570.090 2173.320 2570.410 2173.380 ;
      LAYER via ;
        RECT 2570.120 2429.000 2570.380 2429.260 ;
        RECT 2899.480 2429.000 2899.740 2429.260 ;
        RECT 2523.200 2173.320 2523.460 2173.580 ;
        RECT 2570.120 2173.320 2570.380 2173.580 ;
      LAYER met2 ;
        RECT 2899.470 2433.875 2899.750 2434.245 ;
        RECT 2899.540 2429.290 2899.680 2433.875 ;
        RECT 2570.120 2428.970 2570.380 2429.290 ;
        RECT 2899.480 2428.970 2899.740 2429.290 ;
        RECT 2570.180 2173.610 2570.320 2428.970 ;
        RECT 2523.200 2173.290 2523.460 2173.610 ;
        RECT 2570.120 2173.290 2570.380 2173.610 ;
        RECT 2523.260 2167.005 2523.400 2173.290 ;
        RECT 2523.190 2166.635 2523.470 2167.005 ;
      LAYER via2 ;
        RECT 2899.470 2433.920 2899.750 2434.200 ;
        RECT 2523.190 2166.680 2523.470 2166.960 ;
      LAYER met3 ;
        RECT 2899.445 2434.210 2899.775 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2899.445 2433.910 2924.800 2434.210 ;
        RECT 2899.445 2433.895 2899.775 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2506.000 2166.970 2510.000 2167.120 ;
        RECT 2523.165 2166.970 2523.495 2166.985 ;
        RECT 2506.000 2166.670 2523.495 2166.970 ;
        RECT 2506.000 2166.520 2510.000 2166.670 ;
        RECT 2523.165 2166.655 2523.495 2166.670 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2597.690 2663.800 2598.010 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2597.690 2663.660 2901.150 2663.800 ;
        RECT 2597.690 2663.600 2598.010 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2525.010 2331.960 2525.330 2332.020 ;
        RECT 2597.690 2331.960 2598.010 2332.020 ;
        RECT 2525.010 2331.820 2598.010 2331.960 ;
        RECT 2525.010 2331.760 2525.330 2331.820 ;
        RECT 2597.690 2331.760 2598.010 2331.820 ;
      LAYER via ;
        RECT 2597.720 2663.600 2597.980 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2525.040 2331.760 2525.300 2332.020 ;
        RECT 2597.720 2331.760 2597.980 2332.020 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2597.720 2663.570 2597.980 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2597.780 2332.050 2597.920 2663.570 ;
        RECT 2525.040 2331.730 2525.300 2332.050 ;
        RECT 2597.720 2331.730 2597.980 2332.050 ;
        RECT 2525.100 2330.205 2525.240 2331.730 ;
        RECT 2525.030 2329.835 2525.310 2330.205 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2525.030 2329.880 2525.310 2330.160 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2506.000 2330.170 2510.000 2330.320 ;
        RECT 2525.005 2330.170 2525.335 2330.185 ;
        RECT 2506.000 2329.870 2525.335 2330.170 ;
        RECT 2506.000 2329.720 2510.000 2329.870 ;
        RECT 2525.005 2329.855 2525.335 2329.870 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.090 2898.400 2570.410 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2570.090 2898.260 2901.150 2898.400 ;
        RECT 2570.090 2898.200 2570.410 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2525.010 2497.540 2525.330 2497.600 ;
        RECT 2570.090 2497.540 2570.410 2497.600 ;
        RECT 2525.010 2497.400 2570.410 2497.540 ;
        RECT 2525.010 2497.340 2525.330 2497.400 ;
        RECT 2570.090 2497.340 2570.410 2497.400 ;
      LAYER via ;
        RECT 2570.120 2898.200 2570.380 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2525.040 2497.340 2525.300 2497.600 ;
        RECT 2570.120 2497.340 2570.380 2497.600 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2570.120 2898.170 2570.380 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2570.180 2497.630 2570.320 2898.170 ;
        RECT 2525.040 2497.310 2525.300 2497.630 ;
        RECT 2570.120 2497.310 2570.380 2497.630 ;
        RECT 2525.100 2492.725 2525.240 2497.310 ;
        RECT 2525.030 2492.355 2525.310 2492.725 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2525.030 2492.400 2525.310 2492.680 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2506.000 2492.690 2510.000 2492.840 ;
        RECT 2525.005 2492.690 2525.335 2492.705 ;
        RECT 2506.000 2492.390 2525.335 2492.690 ;
        RECT 2506.000 2492.240 2510.000 2492.390 ;
        RECT 2525.005 2492.375 2525.335 2492.390 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2597.690 3133.000 2598.010 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2597.690 3132.860 2901.150 3133.000 ;
        RECT 2597.690 3132.800 2598.010 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2521.790 2687.600 2522.110 2687.660 ;
        RECT 2597.690 2687.600 2598.010 2687.660 ;
        RECT 2521.790 2687.460 2598.010 2687.600 ;
        RECT 2521.790 2687.400 2522.110 2687.460 ;
        RECT 2597.690 2687.400 2598.010 2687.460 ;
      LAYER via ;
        RECT 2597.720 3132.800 2597.980 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2521.820 2687.400 2522.080 2687.660 ;
        RECT 2597.720 2687.400 2597.980 2687.660 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2597.720 3132.770 2597.980 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2597.780 2687.690 2597.920 3132.770 ;
        RECT 2521.820 2687.370 2522.080 2687.690 ;
        RECT 2597.720 2687.370 2597.980 2687.690 ;
        RECT 2521.880 2655.925 2522.020 2687.370 ;
        RECT 2521.810 2655.555 2522.090 2655.925 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2521.810 2655.600 2522.090 2655.880 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2506.000 2655.890 2510.000 2656.040 ;
        RECT 2521.785 2655.890 2522.115 2655.905 ;
        RECT 2506.000 2655.590 2522.115 2655.890 ;
        RECT 2506.000 2655.440 2510.000 2655.590 ;
        RECT 2521.785 2655.575 2522.115 2655.590 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.090 3367.600 2570.410 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2570.090 3367.460 2901.150 3367.600 ;
        RECT 2570.090 3367.400 2570.410 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2521.790 2908.260 2522.110 2908.320 ;
        RECT 2570.090 2908.260 2570.410 2908.320 ;
        RECT 2521.790 2908.120 2570.410 2908.260 ;
        RECT 2521.790 2908.060 2522.110 2908.120 ;
        RECT 2570.090 2908.060 2570.410 2908.120 ;
      LAYER via ;
        RECT 2570.120 3367.400 2570.380 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2521.820 2908.060 2522.080 2908.320 ;
        RECT 2570.120 2908.060 2570.380 2908.320 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2570.120 3367.370 2570.380 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2570.180 2908.350 2570.320 3367.370 ;
        RECT 2521.820 2908.030 2522.080 2908.350 ;
        RECT 2570.120 2908.030 2570.380 2908.350 ;
        RECT 2521.880 2819.125 2522.020 2908.030 ;
        RECT 2521.810 2818.755 2522.090 2819.125 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2521.810 2818.800 2522.090 2819.080 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2506.000 2819.090 2510.000 2819.240 ;
        RECT 2521.785 2819.090 2522.115 2819.105 ;
        RECT 2506.000 2818.790 2522.115 2819.090 ;
        RECT 2506.000 2818.640 2510.000 2818.790 ;
        RECT 2521.785 2818.775 2522.115 2818.790 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3415.555 ;
      LAYER mcon ;
        RECT 2796.485 3415.385 2796.655 3415.555 ;
      LAYER met1 ;
        RECT 2794.570 3422.340 2794.890 3422.400 ;
        RECT 2798.250 3422.340 2798.570 3422.400 ;
        RECT 2794.570 3422.200 2798.570 3422.340 ;
        RECT 2794.570 3422.140 2794.890 3422.200 ;
        RECT 2798.250 3422.140 2798.570 3422.200 ;
        RECT 2794.570 3415.540 2794.890 3415.600 ;
        RECT 2796.425 3415.540 2796.715 3415.585 ;
        RECT 2794.570 3415.400 2796.715 3415.540 ;
        RECT 2794.570 3415.340 2794.890 3415.400 ;
        RECT 2796.425 3415.355 2796.715 3415.400 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2475.330 3018.760 2475.650 3018.820 ;
        RECT 2795.030 3018.760 2795.350 3018.820 ;
        RECT 2475.330 3018.620 2795.350 3018.760 ;
        RECT 2475.330 3018.560 2475.650 3018.620 ;
        RECT 2795.030 3018.560 2795.350 3018.620 ;
      LAYER via ;
        RECT 2794.600 3422.140 2794.860 3422.400 ;
        RECT 2798.280 3422.140 2798.540 3422.400 ;
        RECT 2794.600 3415.340 2794.860 3415.600 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2475.360 3018.560 2475.620 3018.820 ;
        RECT 2795.060 3018.560 2795.320 3018.820 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.430 2798.480 3517.600 ;
        RECT 2794.600 3422.110 2794.860 3422.430 ;
        RECT 2798.280 3422.110 2798.540 3422.430 ;
        RECT 2794.660 3415.630 2794.800 3422.110 ;
        RECT 2794.600 3415.310 2794.860 3415.630 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3018.850 2795.260 3056.610 ;
        RECT 2475.360 3018.530 2475.620 3018.850 ;
        RECT 2795.060 3018.530 2795.320 3018.850 ;
        RECT 2475.420 3010.000 2475.560 3018.530 ;
        RECT 2475.420 3009.340 2475.770 3010.000 ;
        RECT 2475.490 3006.000 2475.770 3009.340 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2470.270 3464.160 2470.590 3464.220 ;
        RECT 2474.410 3464.160 2474.730 3464.220 ;
        RECT 2470.270 3464.020 2474.730 3464.160 ;
        RECT 2470.270 3463.960 2470.590 3464.020 ;
        RECT 2474.410 3463.960 2474.730 3464.020 ;
        RECT 2470.270 3367.600 2470.590 3367.660 ;
        RECT 2471.190 3367.600 2471.510 3367.660 ;
        RECT 2470.270 3367.460 2471.510 3367.600 ;
        RECT 2470.270 3367.400 2470.590 3367.460 ;
        RECT 2471.190 3367.400 2471.510 3367.460 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2272.010 3018.760 2272.330 3018.820 ;
        RECT 2471.190 3018.760 2471.510 3018.820 ;
        RECT 2272.010 3018.620 2471.510 3018.760 ;
        RECT 2272.010 3018.560 2272.330 3018.620 ;
        RECT 2471.190 3018.560 2471.510 3018.620 ;
      LAYER via ;
        RECT 2470.300 3463.960 2470.560 3464.220 ;
        RECT 2474.440 3463.960 2474.700 3464.220 ;
        RECT 2470.300 3367.400 2470.560 3367.660 ;
        RECT 2471.220 3367.400 2471.480 3367.660 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2272.040 3018.560 2272.300 3018.820 ;
        RECT 2471.220 3018.560 2471.480 3018.820 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3464.250 2474.640 3517.230 ;
        RECT 2470.300 3463.930 2470.560 3464.250 ;
        RECT 2474.440 3463.930 2474.700 3464.250 ;
        RECT 2470.360 3415.370 2470.500 3463.930 ;
        RECT 2470.360 3415.230 2471.420 3415.370 ;
        RECT 2471.280 3367.690 2471.420 3415.230 ;
        RECT 2470.300 3367.370 2470.560 3367.690 ;
        RECT 2471.220 3367.370 2471.480 3367.690 ;
        RECT 2470.360 3318.810 2470.500 3367.370 ;
        RECT 2470.360 3318.670 2471.420 3318.810 ;
        RECT 2471.280 3270.790 2471.420 3318.670 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 3018.850 2471.420 3028.990 ;
        RECT 2272.040 3018.530 2272.300 3018.850 ;
        RECT 2471.220 3018.530 2471.480 3018.850 ;
        RECT 2272.100 3010.000 2272.240 3018.530 ;
        RECT 2272.100 3009.340 2272.450 3010.000 ;
        RECT 2272.170 3006.000 2272.450 3009.340 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3415.555 ;
      LAYER mcon ;
        RECT 2147.885 3415.385 2148.055 3415.555 ;
      LAYER met1 ;
        RECT 2145.970 3422.340 2146.290 3422.400 ;
        RECT 2149.190 3422.340 2149.510 3422.400 ;
        RECT 2145.970 3422.200 2149.510 3422.340 ;
        RECT 2145.970 3422.140 2146.290 3422.200 ;
        RECT 2149.190 3422.140 2149.510 3422.200 ;
        RECT 2145.970 3415.540 2146.290 3415.600 ;
        RECT 2147.825 3415.540 2148.115 3415.585 ;
        RECT 2145.970 3415.400 2148.115 3415.540 ;
        RECT 2145.970 3415.340 2146.290 3415.400 ;
        RECT 2147.825 3415.355 2148.115 3415.400 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2069.150 3018.760 2069.470 3018.820 ;
        RECT 2146.430 3018.760 2146.750 3018.820 ;
        RECT 2069.150 3018.620 2146.750 3018.760 ;
        RECT 2069.150 3018.560 2069.470 3018.620 ;
        RECT 2146.430 3018.560 2146.750 3018.620 ;
      LAYER via ;
        RECT 2146.000 3422.140 2146.260 3422.400 ;
        RECT 2149.220 3422.140 2149.480 3422.400 ;
        RECT 2146.000 3415.340 2146.260 3415.600 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2069.180 3018.560 2069.440 3018.820 ;
        RECT 2146.460 3018.560 2146.720 3018.820 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3422.430 2149.420 3517.600 ;
        RECT 2146.000 3422.110 2146.260 3422.430 ;
        RECT 2149.220 3422.110 2149.480 3422.430 ;
        RECT 2146.060 3415.630 2146.200 3422.110 ;
        RECT 2146.000 3415.310 2146.260 3415.630 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3018.850 2146.660 3056.610 ;
        RECT 2069.180 3018.530 2069.440 3018.850 ;
        RECT 2146.460 3018.530 2146.720 3018.850 ;
        RECT 2069.240 3010.000 2069.380 3018.530 ;
        RECT 2069.240 3009.340 2069.590 3010.000 ;
        RECT 2069.310 3006.000 2069.590 3009.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
        RECT 1828.110 3016.380 1828.430 3016.440 ;
        RECT 1865.830 3016.380 1866.150 3016.440 ;
        RECT 1828.110 3016.240 1866.150 3016.380 ;
        RECT 1828.110 3016.180 1828.430 3016.240 ;
        RECT 1865.830 3016.180 1866.150 3016.240 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
        RECT 1828.140 3016.180 1828.400 3016.440 ;
        RECT 1865.860 3016.180 1866.120 3016.440 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3016.470 1828.340 3498.270 ;
        RECT 1828.140 3016.150 1828.400 3016.470 ;
        RECT 1865.860 3016.150 1866.120 3016.470 ;
        RECT 1865.920 3010.000 1866.060 3016.150 ;
        RECT 1865.920 3009.340 1866.270 3010.000 ;
        RECT 1865.990 3006.000 1866.270 3009.340 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3019.440 1504.130 3019.500 ;
        RECT 1662.510 3019.440 1662.830 3019.500 ;
        RECT 1503.810 3019.300 1662.830 3019.440 ;
        RECT 1503.810 3019.240 1504.130 3019.300 ;
        RECT 1662.510 3019.240 1662.830 3019.300 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3019.240 1504.100 3019.500 ;
        RECT 1662.540 3019.240 1662.800 3019.500 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3019.530 1504.040 3498.270 ;
        RECT 1503.840 3019.210 1504.100 3019.530 ;
        RECT 1662.540 3019.210 1662.800 3019.530 ;
        RECT 1662.600 3010.000 1662.740 3019.210 ;
        RECT 1662.600 3009.340 1662.950 3010.000 ;
        RECT 1662.670 3006.000 1662.950 3009.340 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 697.240 2525.330 697.300 ;
        RECT 2597.690 697.240 2598.010 697.300 ;
        RECT 2525.010 697.100 2598.010 697.240 ;
        RECT 2525.010 697.040 2525.330 697.100 ;
        RECT 2597.690 697.040 2598.010 697.100 ;
        RECT 2597.690 324.260 2598.010 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2597.690 324.120 2899.310 324.260 ;
        RECT 2597.690 324.060 2598.010 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2525.040 697.040 2525.300 697.300 ;
        RECT 2597.720 697.040 2597.980 697.300 ;
        RECT 2597.720 324.060 2597.980 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2525.030 699.195 2525.310 699.565 ;
        RECT 2525.100 697.330 2525.240 699.195 ;
        RECT 2525.040 697.010 2525.300 697.330 ;
        RECT 2597.720 697.010 2597.980 697.330 ;
        RECT 2597.780 324.350 2597.920 697.010 ;
        RECT 2597.720 324.030 2597.980 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2525.030 699.240 2525.310 699.520 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2506.000 699.530 2510.000 699.680 ;
        RECT 2525.005 699.530 2525.335 699.545 ;
        RECT 2506.000 699.230 2525.335 699.530 ;
        RECT 2506.000 699.080 2510.000 699.230 ;
        RECT 2525.005 699.215 2525.335 699.230 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3020.120 1179.830 3020.180 ;
        RECT 1459.190 3020.120 1459.510 3020.180 ;
        RECT 1179.510 3019.980 1459.510 3020.120 ;
        RECT 1179.510 3019.920 1179.830 3019.980 ;
        RECT 1459.190 3019.920 1459.510 3019.980 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3019.920 1179.800 3020.180 ;
        RECT 1459.220 3019.920 1459.480 3020.180 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3020.210 1179.740 3498.270 ;
        RECT 1179.540 3019.890 1179.800 3020.210 ;
        RECT 1459.220 3019.890 1459.480 3020.210 ;
        RECT 1459.280 3010.000 1459.420 3019.890 ;
        RECT 1459.280 3009.340 1459.630 3010.000 ;
        RECT 1459.350 3006.000 1459.630 3009.340 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 3019.100 855.530 3019.160 ;
        RECT 1256.330 3019.100 1256.650 3019.160 ;
        RECT 855.210 3018.960 1256.650 3019.100 ;
        RECT 855.210 3018.900 855.530 3018.960 ;
        RECT 1256.330 3018.900 1256.650 3018.960 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 3018.900 855.500 3019.160 ;
        RECT 1256.360 3018.900 1256.620 3019.160 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 3019.190 855.440 3500.990 ;
        RECT 855.240 3018.870 855.500 3019.190 ;
        RECT 1256.360 3018.870 1256.620 3019.190 ;
        RECT 1256.420 3010.000 1256.560 3018.870 ;
        RECT 1256.420 3009.340 1256.770 3010.000 ;
        RECT 1256.490 3006.000 1256.770 3009.340 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 3020.460 531.230 3020.520 ;
        RECT 1053.010 3020.460 1053.330 3020.520 ;
        RECT 530.910 3020.320 1053.330 3020.460 ;
        RECT 530.910 3020.260 531.230 3020.320 ;
        RECT 1053.010 3020.260 1053.330 3020.320 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 3020.260 531.200 3020.520 ;
        RECT 1053.040 3020.260 1053.300 3020.520 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3020.550 531.140 3498.270 ;
        RECT 530.940 3020.230 531.200 3020.550 ;
        RECT 1053.040 3020.230 1053.300 3020.550 ;
        RECT 1053.100 3010.000 1053.240 3020.230 ;
        RECT 1053.100 3009.340 1053.450 3010.000 ;
        RECT 1053.170 3006.000 1053.450 3009.340 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 3019.440 206.930 3019.500 ;
        RECT 849.690 3019.440 850.010 3019.500 ;
        RECT 206.610 3019.300 850.010 3019.440 ;
        RECT 206.610 3019.240 206.930 3019.300 ;
        RECT 849.690 3019.240 850.010 3019.300 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 3019.240 206.900 3019.500 ;
        RECT 849.720 3019.240 849.980 3019.500 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 3019.530 206.840 3501.670 ;
        RECT 206.640 3019.210 206.900 3019.530 ;
        RECT 849.720 3019.210 849.980 3019.530 ;
        RECT 849.780 3010.000 849.920 3019.210 ;
        RECT 849.780 3009.340 850.130 3010.000 ;
        RECT 849.850 3006.000 850.130 3009.340 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 44.690 3408.740 45.010 3408.800 ;
        RECT 17.550 3408.600 45.010 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 44.690 3408.540 45.010 3408.600 ;
        RECT 44.690 2980.680 45.010 2980.740 ;
        RECT 393.370 2980.680 393.690 2980.740 ;
        RECT 44.690 2980.540 393.690 2980.680 ;
        RECT 44.690 2980.480 45.010 2980.540 ;
        RECT 393.370 2980.480 393.690 2980.540 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 44.720 3408.540 44.980 3408.800 ;
        RECT 44.720 2980.480 44.980 2980.740 ;
        RECT 393.400 2980.480 393.660 2980.740 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 44.720 3408.510 44.980 3408.830 ;
        RECT 44.780 2980.770 44.920 3408.510 ;
        RECT 44.720 2980.450 44.980 2980.770 ;
        RECT 393.400 2980.450 393.660 2980.770 ;
        RECT 393.460 2980.285 393.600 2980.450 ;
        RECT 393.390 2979.915 393.670 2980.285 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 393.390 2979.960 393.670 2980.240 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 393.365 2980.250 393.695 2980.265 ;
        RECT 410.000 2980.250 414.000 2980.400 ;
        RECT 393.365 2979.950 414.000 2980.250 ;
        RECT 393.365 2979.935 393.695 2979.950 ;
        RECT 410.000 2979.800 414.000 2979.950 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 51.590 3119.060 51.910 3119.120 ;
        RECT 16.170 3118.920 51.910 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 51.590 3118.860 51.910 3118.920 ;
        RECT 51.590 2808.300 51.910 2808.360 ;
        RECT 393.370 2808.300 393.690 2808.360 ;
        RECT 51.590 2808.160 393.690 2808.300 ;
        RECT 51.590 2808.100 51.910 2808.160 ;
        RECT 393.370 2808.100 393.690 2808.160 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 51.620 3118.860 51.880 3119.120 ;
        RECT 51.620 2808.100 51.880 2808.360 ;
        RECT 393.400 2808.100 393.660 2808.360 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 51.620 3118.830 51.880 3119.150 ;
        RECT 51.680 2808.390 51.820 3118.830 ;
        RECT 51.620 2808.070 51.880 2808.390 ;
        RECT 393.400 2808.070 393.660 2808.390 ;
        RECT 393.460 2806.205 393.600 2808.070 ;
        RECT 393.390 2805.835 393.670 2806.205 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
        RECT 393.390 2805.880 393.670 2806.160 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
        RECT 393.365 2806.170 393.695 2806.185 ;
        RECT 410.000 2806.170 414.000 2806.320 ;
        RECT 393.365 2805.870 414.000 2806.170 ;
        RECT 393.365 2805.855 393.695 2805.870 ;
        RECT 410.000 2805.720 414.000 2805.870 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 44.690 2836.180 45.010 2836.240 ;
        RECT 17.090 2836.040 45.010 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 44.690 2835.980 45.010 2836.040 ;
        RECT 44.690 2635.580 45.010 2635.640 ;
        RECT 393.370 2635.580 393.690 2635.640 ;
        RECT 44.690 2635.440 393.690 2635.580 ;
        RECT 44.690 2635.380 45.010 2635.440 ;
        RECT 393.370 2635.380 393.690 2635.440 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 44.720 2835.980 44.980 2836.240 ;
        RECT 44.720 2635.380 44.980 2635.640 ;
        RECT 393.400 2635.380 393.660 2635.640 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 44.720 2835.950 44.980 2836.270 ;
        RECT 44.780 2635.670 44.920 2835.950 ;
        RECT 44.720 2635.350 44.980 2635.670 ;
        RECT 393.400 2635.350 393.660 2635.670 ;
        RECT 393.460 2631.445 393.600 2635.350 ;
        RECT 393.390 2631.075 393.670 2631.445 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 393.390 2631.120 393.670 2631.400 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 393.365 2631.410 393.695 2631.425 ;
        RECT 410.000 2631.410 414.000 2631.560 ;
        RECT 393.365 2631.110 414.000 2631.410 ;
        RECT 393.365 2631.095 393.695 2631.110 ;
        RECT 410.000 2630.960 414.000 2631.110 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2463.200 17.410 2463.260 ;
        RECT 393.370 2463.200 393.690 2463.260 ;
        RECT 17.090 2463.060 393.690 2463.200 ;
        RECT 17.090 2463.000 17.410 2463.060 ;
        RECT 393.370 2463.000 393.690 2463.060 ;
      LAYER via ;
        RECT 17.120 2463.000 17.380 2463.260 ;
        RECT 393.400 2463.000 393.660 2463.260 ;
      LAYER met2 ;
        RECT 17.110 2549.475 17.390 2549.845 ;
        RECT 17.180 2463.290 17.320 2549.475 ;
        RECT 17.120 2462.970 17.380 2463.290 ;
        RECT 393.400 2462.970 393.660 2463.290 ;
        RECT 393.460 2457.365 393.600 2462.970 ;
        RECT 393.390 2456.995 393.670 2457.365 ;
      LAYER via2 ;
        RECT 17.110 2549.520 17.390 2549.800 ;
        RECT 393.390 2457.040 393.670 2457.320 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 17.085 2549.810 17.415 2549.825 ;
        RECT -4.800 2549.510 17.415 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 17.085 2549.495 17.415 2549.510 ;
        RECT 393.365 2457.330 393.695 2457.345 ;
        RECT 410.000 2457.330 414.000 2457.480 ;
        RECT 393.365 2457.030 414.000 2457.330 ;
        RECT 393.365 2457.015 393.695 2457.030 ;
        RECT 410.000 2456.880 414.000 2457.030 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 393.370 2262.940 393.690 2263.000 ;
        RECT 17.090 2262.800 393.690 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 393.370 2262.740 393.690 2262.800 ;
      LAYER via ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 393.400 2262.740 393.660 2263.000 ;
      LAYER met2 ;
        RECT 393.390 2282.235 393.670 2282.605 ;
        RECT 393.460 2263.030 393.600 2282.235 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 393.400 2262.710 393.660 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 393.390 2282.280 393.670 2282.560 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT 393.365 2282.570 393.695 2282.585 ;
        RECT 410.000 2282.570 414.000 2282.720 ;
        RECT 393.365 2282.270 414.000 2282.570 ;
        RECT 393.365 2282.255 393.695 2282.270 ;
        RECT 410.000 2282.120 414.000 2282.270 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 397.050 1980.060 397.370 1980.120 ;
        RECT 15.710 1979.920 397.370 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 397.050 1979.860 397.370 1979.920 ;
      LAYER via ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 397.080 1979.860 397.340 1980.120 ;
      LAYER met2 ;
        RECT 397.070 2108.155 397.350 2108.525 ;
        RECT 397.140 1980.150 397.280 2108.155 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 397.080 1979.830 397.340 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 397.070 2108.200 397.350 2108.480 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 397.045 2108.490 397.375 2108.505 ;
        RECT 410.000 2108.490 414.000 2108.640 ;
        RECT 397.045 2108.190 414.000 2108.490 ;
        RECT 397.045 2108.175 397.375 2108.190 ;
        RECT 410.000 2108.040 414.000 2108.190 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2523.630 558.860 2523.950 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2523.630 558.720 2899.310 558.860 ;
        RECT 2523.630 558.660 2523.950 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2523.660 558.660 2523.920 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2523.650 862.395 2523.930 862.765 ;
        RECT 2523.720 558.950 2523.860 862.395 ;
        RECT 2523.660 558.630 2523.920 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2523.650 862.440 2523.930 862.720 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2506.000 862.730 2510.000 862.880 ;
        RECT 2523.625 862.730 2523.955 862.745 ;
        RECT 2506.000 862.430 2523.955 862.730 ;
        RECT 2506.000 862.280 2510.000 862.430 ;
        RECT 2523.625 862.415 2523.955 862.430 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 397.050 1690.380 397.370 1690.440 ;
        RECT 17.090 1690.240 397.370 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 397.050 1690.180 397.370 1690.240 ;
      LAYER via ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 397.080 1690.180 397.340 1690.440 ;
      LAYER met2 ;
        RECT 397.070 1933.395 397.350 1933.765 ;
        RECT 397.140 1690.470 397.280 1933.395 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 397.080 1690.150 397.340 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 397.070 1933.440 397.350 1933.720 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 397.045 1933.730 397.375 1933.745 ;
        RECT 410.000 1933.730 414.000 1933.880 ;
        RECT 397.045 1933.430 414.000 1933.730 ;
        RECT 397.045 1933.415 397.375 1933.430 ;
        RECT 410.000 1933.280 414.000 1933.430 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 397.970 1476.520 398.290 1476.580 ;
        RECT 17.090 1476.380 398.290 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 397.970 1476.320 398.290 1476.380 ;
      LAYER via ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 398.000 1476.320 398.260 1476.580 ;
      LAYER met2 ;
        RECT 397.990 1759.315 398.270 1759.685 ;
        RECT 398.060 1476.610 398.200 1759.315 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 398.000 1476.290 398.260 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 397.990 1759.360 398.270 1759.640 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 397.965 1759.650 398.295 1759.665 ;
        RECT 410.000 1759.650 414.000 1759.800 ;
        RECT 397.965 1759.350 414.000 1759.650 ;
        RECT 397.965 1759.335 398.295 1759.350 ;
        RECT 410.000 1759.200 414.000 1759.350 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 1580.220 45.010 1580.280 ;
        RECT 393.370 1580.220 393.690 1580.280 ;
        RECT 44.690 1580.080 393.690 1580.220 ;
        RECT 44.690 1580.020 45.010 1580.080 ;
        RECT 393.370 1580.020 393.690 1580.080 ;
        RECT 16.170 1262.320 16.490 1262.380 ;
        RECT 44.690 1262.320 45.010 1262.380 ;
        RECT 16.170 1262.180 45.010 1262.320 ;
        RECT 16.170 1262.120 16.490 1262.180 ;
        RECT 44.690 1262.120 45.010 1262.180 ;
      LAYER via ;
        RECT 44.720 1580.020 44.980 1580.280 ;
        RECT 393.400 1580.020 393.660 1580.280 ;
        RECT 16.200 1262.120 16.460 1262.380 ;
        RECT 44.720 1262.120 44.980 1262.380 ;
      LAYER met2 ;
        RECT 393.390 1584.555 393.670 1584.925 ;
        RECT 393.460 1580.310 393.600 1584.555 ;
        RECT 44.720 1579.990 44.980 1580.310 ;
        RECT 393.400 1579.990 393.660 1580.310 ;
        RECT 44.780 1262.410 44.920 1579.990 ;
        RECT 16.200 1262.090 16.460 1262.410 ;
        RECT 44.720 1262.090 44.980 1262.410 ;
        RECT 16.260 1256.485 16.400 1262.090 ;
        RECT 16.190 1256.115 16.470 1256.485 ;
      LAYER via2 ;
        RECT 393.390 1584.600 393.670 1584.880 ;
        RECT 16.190 1256.160 16.470 1256.440 ;
      LAYER met3 ;
        RECT 393.365 1584.890 393.695 1584.905 ;
        RECT 410.000 1584.890 414.000 1585.040 ;
        RECT 393.365 1584.590 414.000 1584.890 ;
        RECT 393.365 1584.575 393.695 1584.590 ;
        RECT 410.000 1584.440 414.000 1584.590 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 16.165 1256.450 16.495 1256.465 ;
        RECT -4.800 1256.150 16.495 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 16.165 1256.135 16.495 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 1407.840 86.410 1407.900 ;
        RECT 393.370 1407.840 393.690 1407.900 ;
        RECT 86.090 1407.700 393.690 1407.840 ;
        RECT 86.090 1407.640 86.410 1407.700 ;
        RECT 393.370 1407.640 393.690 1407.700 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 86.090 1041.660 86.410 1041.720 ;
        RECT 17.090 1041.520 86.410 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 86.090 1041.460 86.410 1041.520 ;
      LAYER via ;
        RECT 86.120 1407.640 86.380 1407.900 ;
        RECT 393.400 1407.640 393.660 1407.900 ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 86.120 1041.460 86.380 1041.720 ;
      LAYER met2 ;
        RECT 393.390 1410.475 393.670 1410.845 ;
        RECT 393.460 1407.930 393.600 1410.475 ;
        RECT 86.120 1407.610 86.380 1407.930 ;
        RECT 393.400 1407.610 393.660 1407.930 ;
        RECT 86.180 1041.750 86.320 1407.610 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 86.120 1041.430 86.380 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 393.390 1410.520 393.670 1410.800 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 393.365 1410.810 393.695 1410.825 ;
        RECT 410.000 1410.810 414.000 1410.960 ;
        RECT 393.365 1410.510 414.000 1410.810 ;
        RECT 393.365 1410.495 393.695 1410.510 ;
        RECT 410.000 1410.360 414.000 1410.510 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 1235.460 141.610 1235.520 ;
        RECT 393.370 1235.460 393.690 1235.520 ;
        RECT 141.290 1235.320 393.690 1235.460 ;
        RECT 141.290 1235.260 141.610 1235.320 ;
        RECT 393.370 1235.260 393.690 1235.320 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 141.290 827.800 141.610 827.860 ;
        RECT 17.550 827.660 141.610 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 141.290 827.600 141.610 827.660 ;
      LAYER via ;
        RECT 141.320 1235.260 141.580 1235.520 ;
        RECT 393.400 1235.260 393.660 1235.520 ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 141.320 827.600 141.580 827.860 ;
      LAYER met2 ;
        RECT 393.390 1235.715 393.670 1236.085 ;
        RECT 393.460 1235.550 393.600 1235.715 ;
        RECT 141.320 1235.230 141.580 1235.550 ;
        RECT 393.400 1235.230 393.660 1235.550 ;
        RECT 141.380 827.890 141.520 1235.230 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 141.320 827.570 141.580 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 393.390 1235.760 393.670 1236.040 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT 393.365 1236.050 393.695 1236.065 ;
        RECT 410.000 1236.050 414.000 1236.200 ;
        RECT 393.365 1235.750 414.000 1236.050 ;
        RECT 393.365 1235.735 393.695 1235.750 ;
        RECT 410.000 1235.600 414.000 1235.750 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 1055.940 45.010 1056.000 ;
        RECT 393.370 1055.940 393.690 1056.000 ;
        RECT 44.690 1055.800 393.690 1055.940 ;
        RECT 44.690 1055.740 45.010 1055.800 ;
        RECT 393.370 1055.740 393.690 1055.800 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 44.690 613.940 45.010 614.000 ;
        RECT 17.090 613.800 45.010 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 44.690 613.740 45.010 613.800 ;
      LAYER via ;
        RECT 44.720 1055.740 44.980 1056.000 ;
        RECT 393.400 1055.740 393.660 1056.000 ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 44.720 613.740 44.980 614.000 ;
      LAYER met2 ;
        RECT 393.390 1061.635 393.670 1062.005 ;
        RECT 393.460 1056.030 393.600 1061.635 ;
        RECT 44.720 1055.710 44.980 1056.030 ;
        RECT 393.400 1055.710 393.660 1056.030 ;
        RECT 44.780 614.030 44.920 1055.710 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 44.720 613.710 44.980 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 393.390 1061.680 393.670 1061.960 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 393.365 1061.970 393.695 1061.985 ;
        RECT 410.000 1061.970 414.000 1062.120 ;
        RECT 393.365 1061.670 414.000 1061.970 ;
        RECT 393.365 1061.655 393.695 1061.670 ;
        RECT 410.000 1061.520 414.000 1061.670 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 883.560 86.410 883.620 ;
        RECT 393.370 883.560 393.690 883.620 ;
        RECT 86.090 883.420 393.690 883.560 ;
        RECT 86.090 883.360 86.410 883.420 ;
        RECT 393.370 883.360 393.690 883.420 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 86.090 400.080 86.410 400.140 ;
        RECT 17.090 399.940 86.410 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 86.090 399.880 86.410 399.940 ;
      LAYER via ;
        RECT 86.120 883.360 86.380 883.620 ;
        RECT 393.400 883.360 393.660 883.620 ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 86.120 399.880 86.380 400.140 ;
      LAYER met2 ;
        RECT 393.390 886.875 393.670 887.245 ;
        RECT 393.460 883.650 393.600 886.875 ;
        RECT 86.120 883.330 86.380 883.650 ;
        RECT 393.400 883.330 393.660 883.650 ;
        RECT 86.180 400.170 86.320 883.330 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 86.120 399.850 86.380 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 393.390 886.920 393.670 887.200 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 393.365 887.210 393.695 887.225 ;
        RECT 410.000 887.210 414.000 887.360 ;
        RECT 393.365 886.910 414.000 887.210 ;
        RECT 393.365 886.895 393.695 886.910 ;
        RECT 410.000 886.760 414.000 886.910 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 710.840 51.910 710.900 ;
        RECT 393.370 710.840 393.690 710.900 ;
        RECT 51.590 710.700 393.690 710.840 ;
        RECT 51.590 710.640 51.910 710.700 ;
        RECT 393.370 710.640 393.690 710.700 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 51.590 179.420 51.910 179.480 ;
        RECT 17.090 179.280 51.910 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 51.590 179.220 51.910 179.280 ;
      LAYER via ;
        RECT 51.620 710.640 51.880 710.900 ;
        RECT 393.400 710.640 393.660 710.900 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 51.620 179.220 51.880 179.480 ;
      LAYER met2 ;
        RECT 393.390 712.795 393.670 713.165 ;
        RECT 393.460 710.930 393.600 712.795 ;
        RECT 51.620 710.610 51.880 710.930 ;
        RECT 393.400 710.610 393.660 710.930 ;
        RECT 51.680 179.510 51.820 710.610 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 51.620 179.190 51.880 179.510 ;
      LAYER via2 ;
        RECT 393.390 712.840 393.670 713.120 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 393.365 713.130 393.695 713.145 ;
        RECT 410.000 713.130 414.000 713.280 ;
        RECT 393.365 712.830 414.000 713.130 ;
        RECT 393.365 712.815 393.695 712.830 ;
        RECT 410.000 712.680 414.000 712.830 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.250 793.460 2522.570 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2522.250 793.320 2899.310 793.460 ;
        RECT 2522.250 793.260 2522.570 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2522.280 793.260 2522.540 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2522.270 1025.595 2522.550 1025.965 ;
        RECT 2522.340 793.550 2522.480 1025.595 ;
        RECT 2522.280 793.230 2522.540 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2522.270 1025.640 2522.550 1025.920 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2506.000 1025.930 2510.000 1026.080 ;
        RECT 2522.245 1025.930 2522.575 1025.945 ;
        RECT 2506.000 1025.630 2522.575 1025.930 ;
        RECT 2506.000 1025.480 2510.000 1025.630 ;
        RECT 2522.245 1025.615 2522.575 1025.630 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1028.060 2522.110 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2521.790 1027.920 2899.310 1028.060 ;
        RECT 2521.790 1027.860 2522.110 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2521.820 1027.860 2522.080 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2521.810 1188.115 2522.090 1188.485 ;
        RECT 2521.880 1028.150 2522.020 1188.115 ;
        RECT 2521.820 1027.830 2522.080 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2521.810 1188.160 2522.090 1188.440 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2506.000 1188.450 2510.000 1188.600 ;
        RECT 2521.785 1188.450 2522.115 1188.465 ;
        RECT 2506.000 1188.150 2522.115 1188.450 ;
        RECT 2506.000 1188.000 2510.000 1188.150 ;
        RECT 2521.785 1188.135 2522.115 1188.150 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1262.660 2522.110 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2521.790 1262.520 2899.310 1262.660 ;
        RECT 2521.790 1262.460 2522.110 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2521.820 1262.460 2522.080 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2521.810 1351.315 2522.090 1351.685 ;
        RECT 2521.880 1262.750 2522.020 1351.315 ;
        RECT 2521.820 1262.430 2522.080 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2521.810 1351.360 2522.090 1351.640 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2506.000 1351.650 2510.000 1351.800 ;
        RECT 2521.785 1351.650 2522.115 1351.665 ;
        RECT 2506.000 1351.350 2522.115 1351.650 ;
        RECT 2506.000 1351.200 2510.000 1351.350 ;
        RECT 2521.785 1351.335 2522.115 1351.350 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.710 1497.260 2523.030 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 2522.710 1497.120 2899.310 1497.260 ;
        RECT 2522.710 1497.060 2523.030 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 2522.740 1497.060 2523.000 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 2522.730 1514.515 2523.010 1514.885 ;
        RECT 2522.800 1497.350 2522.940 1514.515 ;
        RECT 2522.740 1497.030 2523.000 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2522.730 1514.560 2523.010 1514.840 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2506.000 1514.850 2510.000 1515.000 ;
        RECT 2522.705 1514.850 2523.035 1514.865 ;
        RECT 2506.000 1514.550 2523.035 1514.850 ;
        RECT 2506.000 1514.400 2510.000 1514.550 ;
        RECT 2522.705 1514.535 2523.035 1514.550 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.710 1683.580 2523.030 1683.640 ;
        RECT 2901.290 1683.580 2901.610 1683.640 ;
        RECT 2522.710 1683.440 2901.610 1683.580 ;
        RECT 2522.710 1683.380 2523.030 1683.440 ;
        RECT 2901.290 1683.380 2901.610 1683.440 ;
      LAYER via ;
        RECT 2522.740 1683.380 2523.000 1683.640 ;
        RECT 2901.320 1683.380 2901.580 1683.640 ;
      LAYER met2 ;
        RECT 2901.310 1730.075 2901.590 1730.445 ;
        RECT 2901.380 1683.670 2901.520 1730.075 ;
        RECT 2522.740 1683.350 2523.000 1683.670 ;
        RECT 2901.320 1683.350 2901.580 1683.670 ;
        RECT 2522.800 1678.085 2522.940 1683.350 ;
        RECT 2522.730 1677.715 2523.010 1678.085 ;
      LAYER via2 ;
        RECT 2901.310 1730.120 2901.590 1730.400 ;
        RECT 2522.730 1677.760 2523.010 1678.040 ;
      LAYER met3 ;
        RECT 2901.285 1730.410 2901.615 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2901.285 1730.110 2924.800 1730.410 ;
        RECT 2901.285 1730.095 2901.615 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2506.000 1678.050 2510.000 1678.200 ;
        RECT 2522.705 1678.050 2523.035 1678.065 ;
        RECT 2506.000 1677.750 2523.035 1678.050 ;
        RECT 2506.000 1677.600 2510.000 1677.750 ;
        RECT 2522.705 1677.735 2523.035 1677.750 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.090 1960.000 2570.410 1960.060 ;
        RECT 2899.450 1960.000 2899.770 1960.060 ;
        RECT 2570.090 1959.860 2899.770 1960.000 ;
        RECT 2570.090 1959.800 2570.410 1959.860 ;
        RECT 2899.450 1959.800 2899.770 1959.860 ;
        RECT 2525.010 1842.360 2525.330 1842.420 ;
        RECT 2570.090 1842.360 2570.410 1842.420 ;
        RECT 2525.010 1842.220 2570.410 1842.360 ;
        RECT 2525.010 1842.160 2525.330 1842.220 ;
        RECT 2570.090 1842.160 2570.410 1842.220 ;
      LAYER via ;
        RECT 2570.120 1959.800 2570.380 1960.060 ;
        RECT 2899.480 1959.800 2899.740 1960.060 ;
        RECT 2525.040 1842.160 2525.300 1842.420 ;
        RECT 2570.120 1842.160 2570.380 1842.420 ;
      LAYER met2 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
        RECT 2899.540 1960.090 2899.680 1964.675 ;
        RECT 2570.120 1959.770 2570.380 1960.090 ;
        RECT 2899.480 1959.770 2899.740 1960.090 ;
        RECT 2570.180 1842.450 2570.320 1959.770 ;
        RECT 2525.040 1842.130 2525.300 1842.450 ;
        RECT 2570.120 1842.130 2570.380 1842.450 ;
        RECT 2525.100 1840.605 2525.240 1842.130 ;
        RECT 2525.030 1840.235 2525.310 1840.605 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
        RECT 2525.030 1840.280 2525.310 1840.560 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.445 1964.710 2924.800 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2506.000 1840.570 2510.000 1840.720 ;
        RECT 2525.005 1840.570 2525.335 1840.585 ;
        RECT 2506.000 1840.270 2525.335 1840.570 ;
        RECT 2506.000 1840.120 2510.000 1840.270 ;
        RECT 2525.005 1840.255 2525.335 1840.270 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.790 2194.600 2522.110 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2521.790 2194.460 2901.150 2194.600 ;
        RECT 2521.790 2194.400 2522.110 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2521.820 2194.400 2522.080 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2521.820 2194.370 2522.080 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2521.880 2003.805 2522.020 2194.370 ;
        RECT 2521.810 2003.435 2522.090 2003.805 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2521.810 2003.480 2522.090 2003.760 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2506.000 2003.770 2510.000 2003.920 ;
        RECT 2521.785 2003.770 2522.115 2003.785 ;
        RECT 2506.000 2003.470 2522.115 2003.770 ;
        RECT 2506.000 2003.320 2510.000 2003.470 ;
        RECT 2521.785 2003.455 2522.115 2003.470 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 206.960 2522.570 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2522.250 206.820 2901.150 206.960 ;
        RECT 2522.250 206.760 2522.570 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2522.280 206.760 2522.540 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2522.270 644.795 2522.550 645.165 ;
        RECT 2522.340 207.050 2522.480 644.795 ;
        RECT 2522.280 206.730 2522.540 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2522.270 644.840 2522.550 645.120 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2506.000 645.130 2510.000 645.280 ;
        RECT 2522.245 645.130 2522.575 645.145 ;
        RECT 2506.000 644.830 2522.575 645.130 ;
        RECT 2506.000 644.680 2510.000 644.830 ;
        RECT 2522.245 644.815 2522.575 644.830 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2891.170 2548.200 2891.490 2548.260 ;
        RECT 2899.910 2548.200 2900.230 2548.260 ;
        RECT 2891.170 2548.060 2900.230 2548.200 ;
        RECT 2891.170 2548.000 2891.490 2548.060 ;
        RECT 2899.910 2548.000 2900.230 2548.060 ;
        RECT 2521.790 2542.760 2522.110 2542.820 ;
        RECT 2891.170 2542.760 2891.490 2542.820 ;
        RECT 2521.790 2542.620 2891.490 2542.760 ;
        RECT 2521.790 2542.560 2522.110 2542.620 ;
        RECT 2891.170 2542.560 2891.490 2542.620 ;
      LAYER via ;
        RECT 2891.200 2548.000 2891.460 2548.260 ;
        RECT 2899.940 2548.000 2900.200 2548.260 ;
        RECT 2521.820 2542.560 2522.080 2542.820 ;
        RECT 2891.200 2542.560 2891.460 2542.820 ;
      LAYER met2 ;
        RECT 2899.930 2551.515 2900.210 2551.885 ;
        RECT 2900.000 2548.290 2900.140 2551.515 ;
        RECT 2891.200 2547.970 2891.460 2548.290 ;
        RECT 2899.940 2547.970 2900.200 2548.290 ;
        RECT 2891.260 2542.850 2891.400 2547.970 ;
        RECT 2521.820 2542.530 2522.080 2542.850 ;
        RECT 2891.200 2542.530 2891.460 2542.850 ;
        RECT 2521.880 2275.805 2522.020 2542.530 ;
        RECT 2521.810 2275.435 2522.090 2275.805 ;
      LAYER via2 ;
        RECT 2899.930 2551.560 2900.210 2551.840 ;
        RECT 2521.810 2275.480 2522.090 2275.760 ;
      LAYER met3 ;
        RECT 2899.905 2551.850 2900.235 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2899.905 2551.550 2924.800 2551.850 ;
        RECT 2899.905 2551.535 2900.235 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2506.000 2275.770 2510.000 2275.920 ;
        RECT 2521.785 2275.770 2522.115 2275.785 ;
        RECT 2506.000 2275.470 2522.115 2275.770 ;
        RECT 2506.000 2275.320 2510.000 2275.470 ;
        RECT 2521.785 2275.455 2522.115 2275.470 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2549.390 2781.100 2549.710 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2549.390 2780.960 2901.150 2781.100 ;
        RECT 2549.390 2780.900 2549.710 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2525.010 2437.360 2525.330 2437.420 ;
        RECT 2549.390 2437.360 2549.710 2437.420 ;
        RECT 2525.010 2437.220 2549.710 2437.360 ;
        RECT 2525.010 2437.160 2525.330 2437.220 ;
        RECT 2549.390 2437.160 2549.710 2437.220 ;
      LAYER via ;
        RECT 2549.420 2780.900 2549.680 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2525.040 2437.160 2525.300 2437.420 ;
        RECT 2549.420 2437.160 2549.680 2437.420 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2549.420 2780.870 2549.680 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2525.030 2437.955 2525.310 2438.325 ;
        RECT 2525.100 2437.450 2525.240 2437.955 ;
        RECT 2549.480 2437.450 2549.620 2780.870 ;
        RECT 2525.040 2437.130 2525.300 2437.450 ;
        RECT 2549.420 2437.130 2549.680 2437.450 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2525.030 2438.000 2525.310 2438.280 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2506.000 2438.290 2510.000 2438.440 ;
        RECT 2525.005 2438.290 2525.335 2438.305 ;
        RECT 2506.000 2437.990 2525.335 2438.290 ;
        RECT 2506.000 2437.840 2510.000 2437.990 ;
        RECT 2525.005 2437.975 2525.335 2437.990 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2804.690 3015.700 2805.010 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2804.690 3015.560 2901.150 3015.700 ;
        RECT 2804.690 3015.500 2805.010 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2523.170 2608.040 2523.490 2608.100 ;
        RECT 2804.690 2608.040 2805.010 2608.100 ;
        RECT 2523.170 2607.900 2805.010 2608.040 ;
        RECT 2523.170 2607.840 2523.490 2607.900 ;
        RECT 2804.690 2607.840 2805.010 2607.900 ;
      LAYER via ;
        RECT 2804.720 3015.500 2804.980 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2523.200 2607.840 2523.460 2608.100 ;
        RECT 2804.720 2607.840 2804.980 2608.100 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2804.720 3015.470 2804.980 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2804.780 2608.130 2804.920 3015.470 ;
        RECT 2523.200 2607.810 2523.460 2608.130 ;
        RECT 2804.720 2607.810 2804.980 2608.130 ;
        RECT 2523.260 2601.525 2523.400 2607.810 ;
        RECT 2523.190 2601.155 2523.470 2601.525 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2523.190 2601.200 2523.470 2601.480 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2506.000 2601.490 2510.000 2601.640 ;
        RECT 2523.165 2601.490 2523.495 2601.505 ;
        RECT 2506.000 2601.190 2523.495 2601.490 ;
        RECT 2506.000 2601.040 2510.000 2601.190 ;
        RECT 2523.165 2601.175 2523.495 2601.190 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2625.290 3250.300 2625.610 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2625.290 3250.160 2901.150 3250.300 ;
        RECT 2625.290 3250.100 2625.610 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2519.030 2766.820 2519.350 2766.880 ;
        RECT 2625.290 2766.820 2625.610 2766.880 ;
        RECT 2519.030 2766.680 2625.610 2766.820 ;
        RECT 2519.030 2766.620 2519.350 2766.680 ;
        RECT 2625.290 2766.620 2625.610 2766.680 ;
      LAYER via ;
        RECT 2625.320 3250.100 2625.580 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2519.060 2766.620 2519.320 2766.880 ;
        RECT 2625.320 2766.620 2625.580 2766.880 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2625.320 3250.070 2625.580 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2625.380 2766.910 2625.520 3250.070 ;
        RECT 2519.060 2766.590 2519.320 2766.910 ;
        RECT 2625.320 2766.590 2625.580 2766.910 ;
        RECT 2519.120 2764.725 2519.260 2766.590 ;
        RECT 2519.050 2764.355 2519.330 2764.725 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2519.050 2764.400 2519.330 2764.680 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2506.000 2764.690 2510.000 2764.840 ;
        RECT 2519.025 2764.690 2519.355 2764.705 ;
        RECT 2506.000 2764.390 2519.355 2764.690 ;
        RECT 2506.000 2764.240 2510.000 2764.390 ;
        RECT 2519.025 2764.375 2519.355 2764.390 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 3484.900 2522.110 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2521.790 3484.760 2901.150 3484.900 ;
        RECT 2521.790 3484.700 2522.110 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 2521.820 3484.700 2522.080 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2521.820 3484.670 2522.080 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2521.880 2927.925 2522.020 3484.670 ;
        RECT 2521.810 2927.555 2522.090 2927.925 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2521.810 2927.600 2522.090 2927.880 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2506.000 2927.890 2510.000 2928.040 ;
        RECT 2521.785 2927.890 2522.115 2927.905 ;
        RECT 2506.000 2927.590 2522.115 2927.890 ;
        RECT 2506.000 2927.440 2510.000 2927.590 ;
        RECT 2521.785 2927.575 2522.115 2927.590 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2340.090 3019.440 2340.410 3019.500 ;
        RECT 2635.870 3019.440 2636.190 3019.500 ;
        RECT 2340.090 3019.300 2636.190 3019.440 ;
        RECT 2340.090 3019.240 2340.410 3019.300 ;
        RECT 2635.870 3019.240 2636.190 3019.300 ;
      LAYER via ;
        RECT 2340.120 3019.240 2340.380 3019.500 ;
        RECT 2635.900 3019.240 2636.160 3019.500 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3019.530 2636.100 3517.600 ;
        RECT 2340.120 3019.210 2340.380 3019.530 ;
        RECT 2635.900 3019.210 2636.160 3019.530 ;
        RECT 2340.180 3010.000 2340.320 3019.210 ;
        RECT 2340.180 3009.340 2340.530 3010.000 ;
        RECT 2340.250 3006.000 2340.530 3009.340 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2136.770 3019.440 2137.090 3019.500 ;
        RECT 2311.570 3019.440 2311.890 3019.500 ;
        RECT 2136.770 3019.300 2311.890 3019.440 ;
        RECT 2136.770 3019.240 2137.090 3019.300 ;
        RECT 2311.570 3019.240 2311.890 3019.300 ;
      LAYER via ;
        RECT 2136.800 3019.240 2137.060 3019.500 ;
        RECT 2311.600 3019.240 2311.860 3019.500 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3019.530 2311.800 3517.600 ;
        RECT 2136.800 3019.210 2137.060 3019.530 ;
        RECT 2311.600 3019.210 2311.860 3019.530 ;
        RECT 2136.860 3010.000 2137.000 3019.210 ;
        RECT 2136.860 3009.340 2137.210 3010.000 ;
        RECT 2136.930 3006.000 2137.210 3009.340 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1933.450 3018.760 1933.770 3018.820 ;
        RECT 1987.270 3018.760 1987.590 3018.820 ;
        RECT 1933.450 3018.620 1987.590 3018.760 ;
        RECT 1933.450 3018.560 1933.770 3018.620 ;
        RECT 1987.270 3018.560 1987.590 3018.620 ;
      LAYER via ;
        RECT 1933.480 3018.560 1933.740 3018.820 ;
        RECT 1987.300 3018.560 1987.560 3018.820 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3018.850 1987.500 3517.600 ;
        RECT 1933.480 3018.530 1933.740 3018.850 ;
        RECT 1987.300 3018.530 1987.560 3018.850 ;
        RECT 1933.540 3010.000 1933.680 3018.530 ;
        RECT 1933.540 3009.340 1933.890 3010.000 ;
        RECT 1933.610 3006.000 1933.890 3009.340 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1661.590 3018.760 1661.910 3018.820 ;
        RECT 1730.130 3018.760 1730.450 3018.820 ;
        RECT 1661.590 3018.620 1730.450 3018.760 ;
        RECT 1661.590 3018.560 1661.910 3018.620 ;
        RECT 1730.130 3018.560 1730.450 3018.620 ;
      LAYER via ;
        RECT 1661.620 3018.560 1661.880 3018.820 ;
        RECT 1730.160 3018.560 1730.420 3018.820 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3104.610 1662.740 3517.600 ;
        RECT 1662.140 3104.470 1662.740 3104.610 ;
        RECT 1662.140 3057.010 1662.280 3104.470 ;
        RECT 1661.680 3056.870 1662.280 3057.010 ;
        RECT 1661.680 3018.850 1661.820 3056.870 ;
        RECT 1661.620 3018.530 1661.880 3018.850 ;
        RECT 1730.160 3018.530 1730.420 3018.850 ;
        RECT 1730.220 3010.000 1730.360 3018.530 ;
        RECT 1730.220 3009.340 1730.570 3010.000 ;
        RECT 1730.290 3006.000 1730.570 3009.340 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3018.760 1338.530 3018.820 ;
        RECT 1527.270 3018.760 1527.590 3018.820 ;
        RECT 1338.210 3018.620 1527.590 3018.760 ;
        RECT 1338.210 3018.560 1338.530 3018.620 ;
        RECT 1527.270 3018.560 1527.590 3018.620 ;
      LAYER via ;
        RECT 1338.240 3018.560 1338.500 3018.820 ;
        RECT 1527.300 3018.560 1527.560 3018.820 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3018.850 1338.440 3517.600 ;
        RECT 1338.240 3018.530 1338.500 3018.850 ;
        RECT 1527.300 3018.530 1527.560 3018.850 ;
        RECT 1527.360 3010.000 1527.500 3018.530 ;
        RECT 1527.360 3009.340 1527.710 3010.000 ;
        RECT 1527.430 3006.000 1527.710 3009.340 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 441.560 2523.490 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2523.170 441.420 2901.150 441.560 ;
        RECT 2523.170 441.360 2523.490 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2523.200 441.360 2523.460 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2523.190 807.995 2523.470 808.365 ;
        RECT 2523.260 441.650 2523.400 807.995 ;
        RECT 2523.200 441.330 2523.460 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2523.190 808.040 2523.470 808.320 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2506.000 808.330 2510.000 808.480 ;
        RECT 2523.165 808.330 2523.495 808.345 ;
        RECT 2506.000 808.030 2523.495 808.330 ;
        RECT 2506.000 807.880 2510.000 808.030 ;
        RECT 2523.165 808.015 2523.495 808.030 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3019.440 1014.230 3019.500 ;
        RECT 1323.950 3019.440 1324.270 3019.500 ;
        RECT 1013.910 3019.300 1324.270 3019.440 ;
        RECT 1013.910 3019.240 1014.230 3019.300 ;
        RECT 1323.950 3019.240 1324.270 3019.300 ;
      LAYER via ;
        RECT 1013.940 3019.240 1014.200 3019.500 ;
        RECT 1323.980 3019.240 1324.240 3019.500 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3019.530 1014.140 3517.600 ;
        RECT 1013.940 3019.210 1014.200 3019.530 ;
        RECT 1323.980 3019.210 1324.240 3019.530 ;
        RECT 1324.040 3010.000 1324.180 3019.210 ;
        RECT 1324.040 3009.340 1324.390 3010.000 ;
        RECT 1324.110 3006.000 1324.390 3009.340 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3270.700 689.010 3270.760 ;
        RECT 689.610 3270.700 689.930 3270.760 ;
        RECT 688.690 3270.560 689.930 3270.700 ;
        RECT 688.690 3270.500 689.010 3270.560 ;
        RECT 689.610 3270.500 689.930 3270.560 ;
        RECT 688.690 3174.140 689.010 3174.200 ;
        RECT 689.610 3174.140 689.930 3174.200 ;
        RECT 688.690 3174.000 689.930 3174.140 ;
        RECT 688.690 3173.940 689.010 3174.000 ;
        RECT 689.610 3173.940 689.930 3174.000 ;
        RECT 688.690 3077.580 689.010 3077.640 ;
        RECT 689.610 3077.580 689.930 3077.640 ;
        RECT 688.690 3077.440 689.930 3077.580 ;
        RECT 688.690 3077.380 689.010 3077.440 ;
        RECT 689.610 3077.380 689.930 3077.440 ;
        RECT 688.690 3020.800 689.010 3020.860 ;
        RECT 1120.630 3020.800 1120.950 3020.860 ;
        RECT 688.690 3020.660 1120.950 3020.800 ;
        RECT 688.690 3020.600 689.010 3020.660 ;
        RECT 1120.630 3020.600 1120.950 3020.660 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3270.500 688.980 3270.760 ;
        RECT 689.640 3270.500 689.900 3270.760 ;
        RECT 688.720 3173.940 688.980 3174.200 ;
        RECT 689.640 3173.940 689.900 3174.200 ;
        RECT 688.720 3077.380 688.980 3077.640 ;
        RECT 689.640 3077.380 689.900 3077.640 ;
        RECT 688.720 3020.600 688.980 3020.860 ;
        RECT 1120.660 3020.600 1120.920 3020.860 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3270.790 688.920 3318.670 ;
        RECT 688.720 3270.470 688.980 3270.790 ;
        RECT 689.640 3270.470 689.900 3270.790 ;
        RECT 689.700 3222.250 689.840 3270.470 ;
        RECT 688.780 3222.110 689.840 3222.250 ;
        RECT 688.780 3174.230 688.920 3222.110 ;
        RECT 688.720 3173.910 688.980 3174.230 ;
        RECT 689.640 3173.910 689.900 3174.230 ;
        RECT 689.700 3125.690 689.840 3173.910 ;
        RECT 688.780 3125.550 689.840 3125.690 ;
        RECT 688.780 3077.670 688.920 3125.550 ;
        RECT 688.720 3077.350 688.980 3077.670 ;
        RECT 689.640 3077.350 689.900 3077.670 ;
        RECT 689.700 3029.130 689.840 3077.350 ;
        RECT 688.780 3028.990 689.840 3029.130 ;
        RECT 688.780 3020.890 688.920 3028.990 ;
        RECT 688.720 3020.570 688.980 3020.890 ;
        RECT 1120.660 3020.570 1120.920 3020.890 ;
        RECT 1120.720 3010.000 1120.860 3020.570 ;
        RECT 1120.720 3009.340 1121.070 3010.000 ;
        RECT 1120.790 3006.000 1121.070 3009.340 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
        RECT 364.925 3236.205 365.095 3284.315 ;
        RECT 364.005 3139.645 364.175 3187.755 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
        RECT 364.925 3284.145 365.095 3284.315 ;
        RECT 364.005 3187.585 364.175 3187.755 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 364.390 3298.240 364.710 3298.300 ;
        RECT 365.310 3298.240 365.630 3298.300 ;
        RECT 364.390 3298.100 365.630 3298.240 ;
        RECT 364.390 3298.040 364.710 3298.100 ;
        RECT 365.310 3298.040 365.630 3298.100 ;
        RECT 364.865 3284.300 365.155 3284.345 ;
        RECT 365.310 3284.300 365.630 3284.360 ;
        RECT 364.865 3284.160 365.630 3284.300 ;
        RECT 364.865 3284.115 365.155 3284.160 ;
        RECT 365.310 3284.100 365.630 3284.160 ;
        RECT 364.850 3236.360 365.170 3236.420 ;
        RECT 364.655 3236.220 365.170 3236.360 ;
        RECT 364.850 3236.160 365.170 3236.220 ;
        RECT 364.850 3202.020 365.170 3202.080 ;
        RECT 364.020 3201.880 365.170 3202.020 ;
        RECT 364.020 3201.400 364.160 3201.880 ;
        RECT 364.850 3201.820 365.170 3201.880 ;
        RECT 363.930 3201.140 364.250 3201.400 ;
        RECT 363.930 3187.740 364.250 3187.800 ;
        RECT 363.735 3187.600 364.250 3187.740 ;
        RECT 363.930 3187.540 364.250 3187.600 ;
        RECT 363.945 3139.800 364.235 3139.845 ;
        RECT 365.310 3139.800 365.630 3139.860 ;
        RECT 363.945 3139.660 365.630 3139.800 ;
        RECT 363.945 3139.615 364.235 3139.660 ;
        RECT 365.310 3139.600 365.630 3139.660 ;
        RECT 365.310 3019.780 365.630 3019.840 ;
        RECT 917.310 3019.780 917.630 3019.840 ;
        RECT 365.310 3019.640 917.630 3019.780 ;
        RECT 365.310 3019.580 365.630 3019.640 ;
        RECT 917.310 3019.580 917.630 3019.640 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 364.420 3298.040 364.680 3298.300 ;
        RECT 365.340 3298.040 365.600 3298.300 ;
        RECT 365.340 3284.100 365.600 3284.360 ;
        RECT 364.880 3236.160 365.140 3236.420 ;
        RECT 364.880 3201.820 365.140 3202.080 ;
        RECT 363.960 3201.140 364.220 3201.400 ;
        RECT 363.960 3187.540 364.220 3187.800 ;
        RECT 365.340 3139.600 365.600 3139.860 ;
        RECT 365.340 3019.580 365.600 3019.840 ;
        RECT 917.340 3019.580 917.600 3019.840 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.330 364.620 3298.410 ;
        RECT 364.020 3298.270 364.680 3298.330 ;
        RECT 364.420 3298.010 364.680 3298.270 ;
        RECT 365.340 3298.010 365.600 3298.330 ;
        RECT 365.400 3284.390 365.540 3298.010 ;
        RECT 365.340 3284.070 365.600 3284.390 ;
        RECT 364.880 3236.130 365.140 3236.450 ;
        RECT 364.940 3202.110 365.080 3236.130 ;
        RECT 364.880 3201.790 365.140 3202.110 ;
        RECT 363.960 3201.110 364.220 3201.430 ;
        RECT 364.020 3187.830 364.160 3201.110 ;
        RECT 363.960 3187.510 364.220 3187.830 ;
        RECT 365.340 3139.570 365.600 3139.890 ;
        RECT 365.400 3019.870 365.540 3139.570 ;
        RECT 365.340 3019.550 365.600 3019.870 ;
        RECT 917.340 3019.550 917.600 3019.870 ;
        RECT 917.400 3010.000 917.540 3019.550 ;
        RECT 917.400 3009.340 917.750 3010.000 ;
        RECT 917.470 3006.000 917.750 3009.340 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 3018.760 40.410 3018.820 ;
        RECT 714.450 3018.760 714.770 3018.820 ;
        RECT 40.090 3018.620 714.770 3018.760 ;
        RECT 40.090 3018.560 40.410 3018.620 ;
        RECT 714.450 3018.560 714.770 3018.620 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 3018.560 40.380 3018.820 ;
        RECT 714.480 3018.560 714.740 3018.820 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 3018.850 40.320 3028.990 ;
        RECT 40.120 3018.530 40.380 3018.850 ;
        RECT 714.480 3018.530 714.740 3018.850 ;
        RECT 714.540 3010.000 714.680 3018.530 ;
        RECT 714.540 3009.340 714.890 3010.000 ;
        RECT 714.610 3006.000 714.890 3009.340 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 72.290 3263.900 72.610 3263.960 ;
        RECT 15.250 3263.760 72.610 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 72.290 3263.700 72.610 3263.760 ;
        RECT 72.290 2870.180 72.610 2870.240 ;
        RECT 393.370 2870.180 393.690 2870.240 ;
        RECT 72.290 2870.040 393.690 2870.180 ;
        RECT 72.290 2869.980 72.610 2870.040 ;
        RECT 393.370 2869.980 393.690 2870.040 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 72.320 3263.700 72.580 3263.960 ;
        RECT 72.320 2869.980 72.580 2870.240 ;
        RECT 393.400 2869.980 393.660 2870.240 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 72.320 3263.670 72.580 3263.990 ;
        RECT 72.380 2870.270 72.520 3263.670 ;
        RECT 72.320 2869.950 72.580 2870.270 ;
        RECT 393.400 2869.950 393.660 2870.270 ;
        RECT 393.460 2864.005 393.600 2869.950 ;
        RECT 393.390 2863.635 393.670 2864.005 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 393.390 2863.680 393.670 2863.960 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 393.365 2863.970 393.695 2863.985 ;
        RECT 410.000 2863.970 414.000 2864.120 ;
        RECT 393.365 2863.670 414.000 2863.970 ;
        RECT 393.365 2863.655 393.695 2863.670 ;
        RECT 410.000 2863.520 414.000 2863.670 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 45.150 2974.220 45.470 2974.280 ;
        RECT 16.630 2974.080 45.470 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 45.150 2974.020 45.470 2974.080 ;
        RECT 45.150 2839.240 45.470 2839.300 ;
        RECT 396.590 2839.240 396.910 2839.300 ;
        RECT 45.150 2839.100 396.910 2839.240 ;
        RECT 45.150 2839.040 45.470 2839.100 ;
        RECT 396.590 2839.040 396.910 2839.100 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 45.180 2974.020 45.440 2974.280 ;
        RECT 45.180 2839.040 45.440 2839.300 ;
        RECT 396.620 2839.040 396.880 2839.300 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 45.180 2973.990 45.440 2974.310 ;
        RECT 45.240 2839.330 45.380 2973.990 ;
        RECT 45.180 2839.010 45.440 2839.330 ;
        RECT 396.620 2839.010 396.880 2839.330 ;
        RECT 396.680 2689.925 396.820 2839.010 ;
        RECT 396.610 2689.555 396.890 2689.925 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
        RECT 396.610 2689.600 396.890 2689.880 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
        RECT 396.585 2689.890 396.915 2689.905 ;
        RECT 410.000 2689.890 414.000 2690.040 ;
        RECT 396.585 2689.590 414.000 2689.890 ;
        RECT 396.585 2689.575 396.915 2689.590 ;
        RECT 410.000 2689.440 414.000 2689.590 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2518.280 17.870 2518.340 ;
        RECT 393.370 2518.280 393.690 2518.340 ;
        RECT 17.550 2518.140 393.690 2518.280 ;
        RECT 17.550 2518.080 17.870 2518.140 ;
        RECT 393.370 2518.080 393.690 2518.140 ;
      LAYER via ;
        RECT 17.580 2518.080 17.840 2518.340 ;
        RECT 393.400 2518.080 393.660 2518.340 ;
      LAYER met2 ;
        RECT 17.570 2692.955 17.850 2693.325 ;
        RECT 17.640 2518.370 17.780 2692.955 ;
        RECT 17.580 2518.050 17.840 2518.370 ;
        RECT 393.400 2518.050 393.660 2518.370 ;
        RECT 393.460 2515.165 393.600 2518.050 ;
        RECT 393.390 2514.795 393.670 2515.165 ;
      LAYER via2 ;
        RECT 17.570 2693.000 17.850 2693.280 ;
        RECT 393.390 2514.840 393.670 2515.120 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.545 2693.290 17.875 2693.305 ;
        RECT -4.800 2692.990 17.875 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.545 2692.975 17.875 2692.990 ;
        RECT 393.365 2515.130 393.695 2515.145 ;
        RECT 410.000 2515.130 414.000 2515.280 ;
        RECT 393.365 2514.830 414.000 2515.130 ;
        RECT 393.365 2514.815 393.695 2514.830 ;
        RECT 410.000 2514.680 414.000 2514.830 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2345.900 17.410 2345.960 ;
        RECT 393.370 2345.900 393.690 2345.960 ;
        RECT 17.090 2345.760 393.690 2345.900 ;
        RECT 17.090 2345.700 17.410 2345.760 ;
        RECT 393.370 2345.700 393.690 2345.760 ;
      LAYER via ;
        RECT 17.120 2345.700 17.380 2345.960 ;
        RECT 393.400 2345.700 393.660 2345.960 ;
      LAYER met2 ;
        RECT 17.110 2405.315 17.390 2405.685 ;
        RECT 17.180 2345.990 17.320 2405.315 ;
        RECT 17.120 2345.670 17.380 2345.990 ;
        RECT 393.400 2345.670 393.660 2345.990 ;
        RECT 393.460 2341.085 393.600 2345.670 ;
        RECT 393.390 2340.715 393.670 2341.085 ;
      LAYER via2 ;
        RECT 17.110 2405.360 17.390 2405.640 ;
        RECT 393.390 2340.760 393.670 2341.040 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 17.085 2405.650 17.415 2405.665 ;
        RECT -4.800 2405.350 17.415 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 17.085 2405.335 17.415 2405.350 ;
        RECT 393.365 2341.050 393.695 2341.065 ;
        RECT 410.000 2341.050 414.000 2341.200 ;
        RECT 393.365 2340.750 414.000 2341.050 ;
        RECT 393.365 2340.735 393.695 2340.750 ;
        RECT 410.000 2340.600 414.000 2340.750 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 396.590 2125.240 396.910 2125.300 ;
        RECT 16.170 2125.100 396.910 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 396.590 2125.040 396.910 2125.100 ;
      LAYER via ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 396.620 2125.040 396.880 2125.300 ;
      LAYER met2 ;
        RECT 396.610 2165.955 396.890 2166.325 ;
        RECT 396.680 2125.330 396.820 2165.955 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 396.620 2125.010 396.880 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 396.610 2166.000 396.890 2166.280 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT 396.585 2166.290 396.915 2166.305 ;
        RECT 410.000 2166.290 414.000 2166.440 ;
        RECT 396.585 2165.990 414.000 2166.290 ;
        RECT 396.585 2165.975 396.915 2165.990 ;
        RECT 410.000 2165.840 414.000 2165.990 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 396.590 1835.220 396.910 1835.280 ;
        RECT 15.710 1835.080 396.910 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 396.590 1835.020 396.910 1835.080 ;
      LAYER via ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 396.620 1835.020 396.880 1835.280 ;
      LAYER met2 ;
        RECT 396.610 1991.875 396.890 1992.245 ;
        RECT 396.680 1835.310 396.820 1991.875 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 396.620 1834.990 396.880 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 396.610 1991.920 396.890 1992.200 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 396.585 1992.210 396.915 1992.225 ;
        RECT 410.000 1992.210 414.000 1992.360 ;
        RECT 396.585 1991.910 414.000 1992.210 ;
        RECT 396.585 1991.895 396.915 1991.910 ;
        RECT 410.000 1991.760 414.000 1991.910 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 676.160 2522.110 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2521.790 676.020 2901.150 676.160 ;
        RECT 2521.790 675.960 2522.110 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2521.820 675.960 2522.080 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2521.810 971.195 2522.090 971.565 ;
        RECT 2521.880 676.250 2522.020 971.195 ;
        RECT 2521.820 675.930 2522.080 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2521.810 971.240 2522.090 971.520 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2506.000 971.530 2510.000 971.680 ;
        RECT 2521.785 971.530 2522.115 971.545 ;
        RECT 2506.000 971.230 2522.115 971.530 ;
        RECT 2506.000 971.080 2510.000 971.230 ;
        RECT 2521.785 971.215 2522.115 971.230 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 396.590 1545.540 396.910 1545.600 ;
        RECT 16.630 1545.400 396.910 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 396.590 1545.340 396.910 1545.400 ;
      LAYER via ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 396.620 1545.340 396.880 1545.600 ;
      LAYER met2 ;
        RECT 396.610 1817.115 396.890 1817.485 ;
        RECT 396.680 1545.630 396.820 1817.115 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 396.620 1545.310 396.880 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 396.610 1817.160 396.890 1817.440 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 396.585 1817.450 396.915 1817.465 ;
        RECT 410.000 1817.450 414.000 1817.600 ;
        RECT 396.585 1817.150 414.000 1817.450 ;
        RECT 396.585 1817.135 396.915 1817.150 ;
        RECT 410.000 1817.000 414.000 1817.150 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 397.050 1331.680 397.370 1331.740 ;
        RECT 15.710 1331.540 397.370 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 397.050 1331.480 397.370 1331.540 ;
      LAYER via ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 397.080 1331.480 397.340 1331.740 ;
      LAYER met2 ;
        RECT 397.070 1643.035 397.350 1643.405 ;
        RECT 397.140 1331.770 397.280 1643.035 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 397.080 1331.450 397.340 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 397.070 1643.080 397.350 1643.360 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
        RECT 397.045 1643.370 397.375 1643.385 ;
        RECT 410.000 1643.370 414.000 1643.520 ;
        RECT 397.045 1643.070 414.000 1643.370 ;
        RECT 397.045 1643.055 397.375 1643.070 ;
        RECT 410.000 1642.920 414.000 1643.070 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 15.705 1328.215 16.035 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 397.970 1117.820 398.290 1117.880 ;
        RECT 15.710 1117.680 398.290 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 397.970 1117.620 398.290 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 398.000 1117.620 398.260 1117.880 ;
      LAYER met2 ;
        RECT 397.990 1468.275 398.270 1468.645 ;
        RECT 398.060 1117.910 398.200 1468.275 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 398.000 1117.590 398.260 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 397.990 1468.320 398.270 1468.600 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 397.965 1468.610 398.295 1468.625 ;
        RECT 410.000 1468.610 414.000 1468.760 ;
        RECT 397.965 1468.310 414.000 1468.610 ;
        RECT 397.965 1468.295 398.295 1468.310 ;
        RECT 410.000 1468.160 414.000 1468.310 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 397.050 903.960 397.370 904.020 ;
        RECT 16.170 903.820 397.370 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 397.050 903.760 397.370 903.820 ;
      LAYER via ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 397.080 903.760 397.340 904.020 ;
      LAYER met2 ;
        RECT 397.070 1294.195 397.350 1294.565 ;
        RECT 397.140 904.050 397.280 1294.195 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 397.080 903.730 397.340 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 397.070 1294.240 397.350 1294.520 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 397.045 1294.530 397.375 1294.545 ;
        RECT 410.000 1294.530 414.000 1294.680 ;
        RECT 397.045 1294.230 414.000 1294.530 ;
        RECT 397.045 1294.215 397.375 1294.230 ;
        RECT 410.000 1294.080 414.000 1294.230 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 1118.160 72.610 1118.220 ;
        RECT 393.370 1118.160 393.690 1118.220 ;
        RECT 72.290 1118.020 393.690 1118.160 ;
        RECT 72.290 1117.960 72.610 1118.020 ;
        RECT 393.370 1117.960 393.690 1118.020 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 72.290 682.960 72.610 683.020 ;
        RECT 16.170 682.820 72.610 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 72.290 682.760 72.610 682.820 ;
      LAYER via ;
        RECT 72.320 1117.960 72.580 1118.220 ;
        RECT 393.400 1117.960 393.660 1118.220 ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 72.320 682.760 72.580 683.020 ;
      LAYER met2 ;
        RECT 393.390 1119.435 393.670 1119.805 ;
        RECT 393.460 1118.250 393.600 1119.435 ;
        RECT 72.320 1117.930 72.580 1118.250 ;
        RECT 393.400 1117.930 393.660 1118.250 ;
        RECT 72.380 683.050 72.520 1117.930 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 72.320 682.730 72.580 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 393.390 1119.480 393.670 1119.760 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 393.365 1119.770 393.695 1119.785 ;
        RECT 410.000 1119.770 414.000 1119.920 ;
        RECT 393.365 1119.470 414.000 1119.770 ;
        RECT 393.365 1119.455 393.695 1119.470 ;
        RECT 410.000 1119.320 414.000 1119.470 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 945.440 100.210 945.500 ;
        RECT 393.370 945.440 393.690 945.500 ;
        RECT 99.890 945.300 393.690 945.440 ;
        RECT 99.890 945.240 100.210 945.300 ;
        RECT 393.370 945.240 393.690 945.300 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 99.890 469.100 100.210 469.160 ;
        RECT 17.090 468.960 100.210 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 99.890 468.900 100.210 468.960 ;
      LAYER via ;
        RECT 99.920 945.240 100.180 945.500 ;
        RECT 393.400 945.240 393.660 945.500 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 99.920 468.900 100.180 469.160 ;
      LAYER met2 ;
        RECT 99.920 945.210 100.180 945.530 ;
        RECT 393.390 945.355 393.670 945.725 ;
        RECT 393.400 945.210 393.660 945.355 ;
        RECT 99.980 469.190 100.120 945.210 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 99.920 468.870 100.180 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 393.390 945.400 393.670 945.680 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 393.365 945.690 393.695 945.705 ;
        RECT 410.000 945.690 414.000 945.840 ;
        RECT 393.365 945.390 414.000 945.690 ;
        RECT 393.365 945.375 393.695 945.390 ;
        RECT 410.000 945.240 414.000 945.390 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 397.510 255.240 397.830 255.300 ;
        RECT 17.090 255.100 397.830 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 397.510 255.040 397.830 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 397.540 255.040 397.800 255.300 ;
      LAYER met2 ;
        RECT 397.530 770.595 397.810 770.965 ;
        RECT 397.600 255.330 397.740 770.595 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 397.540 255.010 397.800 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 397.530 770.640 397.810 770.920 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 397.505 770.930 397.835 770.945 ;
        RECT 410.000 770.930 414.000 771.080 ;
        RECT 397.505 770.630 414.000 770.930 ;
        RECT 397.505 770.615 397.835 770.630 ;
        RECT 410.000 770.480 414.000 770.630 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 41.380 20.630 41.440 ;
        RECT 396.590 41.380 396.910 41.440 ;
        RECT 20.310 41.240 396.910 41.380 ;
        RECT 20.310 41.180 20.630 41.240 ;
        RECT 396.590 41.180 396.910 41.240 ;
      LAYER via ;
        RECT 20.340 41.180 20.600 41.440 ;
        RECT 396.620 41.180 396.880 41.440 ;
      LAYER met2 ;
        RECT 396.610 596.515 396.890 596.885 ;
        RECT 396.680 41.470 396.820 596.515 ;
        RECT 20.340 41.150 20.600 41.470 ;
        RECT 396.620 41.150 396.880 41.470 ;
        RECT 20.400 35.885 20.540 41.150 ;
        RECT 20.330 35.515 20.610 35.885 ;
      LAYER via2 ;
        RECT 396.610 596.560 396.890 596.840 ;
        RECT 20.330 35.560 20.610 35.840 ;
      LAYER met3 ;
        RECT 396.585 596.850 396.915 596.865 ;
        RECT 410.000 596.850 414.000 597.000 ;
        RECT 396.585 596.550 414.000 596.850 ;
        RECT 396.585 596.535 396.915 596.550 ;
        RECT 410.000 596.400 414.000 596.550 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 20.305 35.850 20.635 35.865 ;
        RECT -4.800 35.550 20.635 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 20.305 35.535 20.635 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2523.170 910.760 2523.490 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2523.170 910.620 2901.150 910.760 ;
        RECT 2523.170 910.560 2523.490 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2523.200 910.560 2523.460 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2523.190 1134.395 2523.470 1134.765 ;
        RECT 2523.260 910.850 2523.400 1134.395 ;
        RECT 2523.200 910.530 2523.460 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2523.190 1134.440 2523.470 1134.720 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2506.000 1134.730 2510.000 1134.880 ;
        RECT 2523.165 1134.730 2523.495 1134.745 ;
        RECT 2506.000 1134.430 2523.495 1134.730 ;
        RECT 2506.000 1134.280 2510.000 1134.430 ;
        RECT 2523.165 1134.415 2523.495 1134.430 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 1145.360 2523.030 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2522.710 1145.220 2901.150 1145.360 ;
        RECT 2522.710 1145.160 2523.030 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2522.740 1145.160 2523.000 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2522.730 1296.915 2523.010 1297.285 ;
        RECT 2522.800 1145.450 2522.940 1296.915 ;
        RECT 2522.740 1145.130 2523.000 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2522.730 1296.960 2523.010 1297.240 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2506.000 1297.250 2510.000 1297.400 ;
        RECT 2522.705 1297.250 2523.035 1297.265 ;
        RECT 2506.000 1296.950 2523.035 1297.250 ;
        RECT 2506.000 1296.800 2510.000 1296.950 ;
        RECT 2522.705 1296.935 2523.035 1296.950 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 1379.960 2522.110 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2521.790 1379.820 2901.150 1379.960 ;
        RECT 2521.790 1379.760 2522.110 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2521.820 1379.760 2522.080 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2521.810 1460.115 2522.090 1460.485 ;
        RECT 2521.880 1380.050 2522.020 1460.115 ;
        RECT 2521.820 1379.730 2522.080 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2521.810 1460.160 2522.090 1460.440 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2506.000 1460.450 2510.000 1460.600 ;
        RECT 2521.785 1460.450 2522.115 1460.465 ;
        RECT 2506.000 1460.150 2522.115 1460.450 ;
        RECT 2506.000 1460.000 2510.000 1460.150 ;
        RECT 2521.785 1460.135 2522.115 1460.150 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1614.560 2525.330 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2525.010 1614.420 2901.150 1614.560 ;
        RECT 2525.010 1614.360 2525.330 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2525.040 1614.360 2525.300 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2525.030 1623.315 2525.310 1623.685 ;
        RECT 2525.100 1614.650 2525.240 1623.315 ;
        RECT 2525.040 1614.330 2525.300 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2525.030 1623.360 2525.310 1623.640 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2506.000 1623.650 2510.000 1623.800 ;
        RECT 2525.005 1623.650 2525.335 1623.665 ;
        RECT 2506.000 1623.350 2525.335 1623.650 ;
        RECT 2506.000 1623.200 2510.000 1623.350 ;
        RECT 2525.005 1623.335 2525.335 1623.350 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1786.940 2525.330 1787.000 ;
        RECT 2901.290 1786.940 2901.610 1787.000 ;
        RECT 2525.010 1786.800 2901.610 1786.940 ;
        RECT 2525.010 1786.740 2525.330 1786.800 ;
        RECT 2901.290 1786.740 2901.610 1786.800 ;
      LAYER via ;
        RECT 2525.040 1786.740 2525.300 1787.000 ;
        RECT 2901.320 1786.740 2901.580 1787.000 ;
      LAYER met2 ;
        RECT 2901.310 1847.715 2901.590 1848.085 ;
        RECT 2901.380 1787.030 2901.520 1847.715 ;
        RECT 2525.040 1786.885 2525.300 1787.030 ;
        RECT 2525.030 1786.515 2525.310 1786.885 ;
        RECT 2901.320 1786.710 2901.580 1787.030 ;
      LAYER via2 ;
        RECT 2901.310 1847.760 2901.590 1848.040 ;
        RECT 2525.030 1786.560 2525.310 1786.840 ;
      LAYER met3 ;
        RECT 2901.285 1848.050 2901.615 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.285 1847.750 2924.800 1848.050 ;
        RECT 2901.285 1847.735 2901.615 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2506.000 1786.850 2510.000 1787.000 ;
        RECT 2525.005 1786.850 2525.335 1786.865 ;
        RECT 2506.000 1786.550 2525.335 1786.850 ;
        RECT 2506.000 1786.400 2510.000 1786.550 ;
        RECT 2525.005 1786.535 2525.335 1786.550 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1952.520 2525.330 1952.580 ;
        RECT 2902.210 1952.520 2902.530 1952.580 ;
        RECT 2525.010 1952.380 2902.530 1952.520 ;
        RECT 2525.010 1952.320 2525.330 1952.380 ;
        RECT 2902.210 1952.320 2902.530 1952.380 ;
      LAYER via ;
        RECT 2525.040 1952.320 2525.300 1952.580 ;
        RECT 2902.240 1952.320 2902.500 1952.580 ;
      LAYER met2 ;
        RECT 2902.230 2082.315 2902.510 2082.685 ;
        RECT 2902.300 1952.610 2902.440 2082.315 ;
        RECT 2525.040 1952.290 2525.300 1952.610 ;
        RECT 2902.240 1952.290 2902.500 1952.610 ;
        RECT 2525.100 1949.405 2525.240 1952.290 ;
        RECT 2525.030 1949.035 2525.310 1949.405 ;
      LAYER via2 ;
        RECT 2902.230 2082.360 2902.510 2082.640 ;
        RECT 2525.030 1949.080 2525.310 1949.360 ;
      LAYER met3 ;
        RECT 2902.205 2082.650 2902.535 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2902.205 2082.350 2924.800 2082.650 ;
        RECT 2902.205 2082.335 2902.535 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2506.000 1949.370 2510.000 1949.520 ;
        RECT 2525.005 1949.370 2525.335 1949.385 ;
        RECT 2506.000 1949.070 2525.335 1949.370 ;
        RECT 2506.000 1948.920 2510.000 1949.070 ;
        RECT 2525.005 1949.055 2525.335 1949.070 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2528.690 2311.900 2529.010 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2528.690 2311.760 2901.150 2311.900 ;
        RECT 2528.690 2311.700 2529.010 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 2518.570 2117.420 2518.890 2117.480 ;
        RECT 2528.690 2117.420 2529.010 2117.480 ;
        RECT 2518.570 2117.280 2529.010 2117.420 ;
        RECT 2518.570 2117.220 2518.890 2117.280 ;
        RECT 2528.690 2117.220 2529.010 2117.280 ;
      LAYER via ;
        RECT 2528.720 2311.700 2528.980 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 2518.600 2117.220 2518.860 2117.480 ;
        RECT 2528.720 2117.220 2528.980 2117.480 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2528.720 2311.670 2528.980 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2528.780 2117.510 2528.920 2311.670 ;
        RECT 2518.600 2117.190 2518.860 2117.510 ;
        RECT 2528.720 2117.190 2528.980 2117.510 ;
        RECT 2518.660 2112.605 2518.800 2117.190 ;
        RECT 2518.590 2112.235 2518.870 2112.605 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2518.590 2112.280 2518.870 2112.560 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2506.000 2112.570 2510.000 2112.720 ;
        RECT 2518.565 2112.570 2518.895 2112.585 ;
        RECT 2506.000 2112.270 2518.895 2112.570 ;
        RECT 2506.000 2112.120 2510.000 2112.270 ;
        RECT 2518.565 2112.255 2518.895 2112.270 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 151.540 2522.110 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2521.790 151.400 2901.150 151.540 ;
        RECT 2521.790 151.340 2522.110 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2521.820 151.340 2522.080 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2521.810 590.395 2522.090 590.765 ;
        RECT 2521.880 151.630 2522.020 590.395 ;
        RECT 2521.820 151.310 2522.080 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2521.810 590.440 2522.090 590.720 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2506.000 590.730 2510.000 590.880 ;
        RECT 2521.785 590.730 2522.115 590.745 ;
        RECT 2506.000 590.430 2522.115 590.730 ;
        RECT 2506.000 590.280 2510.000 590.430 ;
        RECT 2521.785 590.415 2522.115 590.430 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2221.800 2525.330 2221.860 ;
        RECT 2901.290 2221.800 2901.610 2221.860 ;
        RECT 2525.010 2221.660 2901.610 2221.800 ;
        RECT 2525.010 2221.600 2525.330 2221.660 ;
        RECT 2901.290 2221.600 2901.610 2221.660 ;
      LAYER via ;
        RECT 2525.040 2221.600 2525.300 2221.860 ;
        RECT 2901.320 2221.600 2901.580 2221.860 ;
      LAYER met2 ;
        RECT 2901.310 2493.035 2901.590 2493.405 ;
        RECT 2901.380 2221.890 2901.520 2493.035 ;
        RECT 2525.040 2221.570 2525.300 2221.890 ;
        RECT 2901.320 2221.570 2901.580 2221.890 ;
        RECT 2525.100 2221.405 2525.240 2221.570 ;
        RECT 2525.030 2221.035 2525.310 2221.405 ;
      LAYER via2 ;
        RECT 2901.310 2493.080 2901.590 2493.360 ;
        RECT 2525.030 2221.080 2525.310 2221.360 ;
      LAYER met3 ;
        RECT 2901.285 2493.370 2901.615 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2901.285 2493.070 2924.800 2493.370 ;
        RECT 2901.285 2493.055 2901.615 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2506.000 2221.370 2510.000 2221.520 ;
        RECT 2525.005 2221.370 2525.335 2221.385 ;
        RECT 2506.000 2221.070 2525.335 2221.370 ;
        RECT 2506.000 2220.920 2510.000 2221.070 ;
        RECT 2525.005 2221.055 2525.335 2221.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2528.690 2725.680 2529.010 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2528.690 2725.540 2901.150 2725.680 ;
        RECT 2528.690 2725.480 2529.010 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 2518.570 2386.360 2518.890 2386.420 ;
        RECT 2528.690 2386.360 2529.010 2386.420 ;
        RECT 2518.570 2386.220 2529.010 2386.360 ;
        RECT 2518.570 2386.160 2518.890 2386.220 ;
        RECT 2528.690 2386.160 2529.010 2386.220 ;
      LAYER via ;
        RECT 2528.720 2725.480 2528.980 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 2518.600 2386.160 2518.860 2386.420 ;
        RECT 2528.720 2386.160 2528.980 2386.420 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2528.720 2725.450 2528.980 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2528.780 2386.450 2528.920 2725.450 ;
        RECT 2518.600 2386.130 2518.860 2386.450 ;
        RECT 2528.720 2386.130 2528.980 2386.450 ;
        RECT 2518.660 2384.605 2518.800 2386.130 ;
        RECT 2518.590 2384.235 2518.870 2384.605 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2518.590 2384.280 2518.870 2384.560 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2506.000 2384.570 2510.000 2384.720 ;
        RECT 2518.565 2384.570 2518.895 2384.585 ;
        RECT 2506.000 2384.270 2518.895 2384.570 ;
        RECT 2506.000 2384.120 2510.000 2384.270 ;
        RECT 2518.565 2384.255 2518.895 2384.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2604.590 2960.280 2604.910 2960.340 ;
        RECT 2899.450 2960.280 2899.770 2960.340 ;
        RECT 2604.590 2960.140 2899.770 2960.280 ;
        RECT 2604.590 2960.080 2604.910 2960.140 ;
        RECT 2899.450 2960.080 2899.770 2960.140 ;
        RECT 2525.010 2552.960 2525.330 2553.020 ;
        RECT 2604.590 2552.960 2604.910 2553.020 ;
        RECT 2525.010 2552.820 2604.910 2552.960 ;
        RECT 2525.010 2552.760 2525.330 2552.820 ;
        RECT 2604.590 2552.760 2604.910 2552.820 ;
      LAYER via ;
        RECT 2604.620 2960.080 2604.880 2960.340 ;
        RECT 2899.480 2960.080 2899.740 2960.340 ;
        RECT 2525.040 2552.760 2525.300 2553.020 ;
        RECT 2604.620 2552.760 2604.880 2553.020 ;
      LAYER met2 ;
        RECT 2899.470 2962.235 2899.750 2962.605 ;
        RECT 2899.540 2960.370 2899.680 2962.235 ;
        RECT 2604.620 2960.050 2604.880 2960.370 ;
        RECT 2899.480 2960.050 2899.740 2960.370 ;
        RECT 2604.680 2553.050 2604.820 2960.050 ;
        RECT 2525.040 2552.730 2525.300 2553.050 ;
        RECT 2604.620 2552.730 2604.880 2553.050 ;
        RECT 2525.100 2547.125 2525.240 2552.730 ;
        RECT 2525.030 2546.755 2525.310 2547.125 ;
      LAYER via2 ;
        RECT 2899.470 2962.280 2899.750 2962.560 ;
        RECT 2525.030 2546.800 2525.310 2547.080 ;
      LAYER met3 ;
        RECT 2899.445 2962.570 2899.775 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2899.445 2962.270 2924.800 2962.570 ;
        RECT 2899.445 2962.255 2899.775 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2506.000 2547.090 2510.000 2547.240 ;
        RECT 2525.005 2547.090 2525.335 2547.105 ;
        RECT 2506.000 2546.790 2525.335 2547.090 ;
        RECT 2506.000 2546.640 2510.000 2546.790 ;
        RECT 2525.005 2546.775 2525.335 2546.790 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2711.740 2525.330 2711.800 ;
        RECT 2901.750 2711.740 2902.070 2711.800 ;
        RECT 2525.010 2711.600 2902.070 2711.740 ;
        RECT 2525.010 2711.540 2525.330 2711.600 ;
        RECT 2901.750 2711.540 2902.070 2711.600 ;
      LAYER via ;
        RECT 2525.040 2711.540 2525.300 2711.800 ;
        RECT 2901.780 2711.540 2902.040 2711.800 ;
      LAYER met2 ;
        RECT 2901.770 3196.835 2902.050 3197.205 ;
        RECT 2901.840 2711.830 2901.980 3196.835 ;
        RECT 2525.040 2711.510 2525.300 2711.830 ;
        RECT 2901.780 2711.510 2902.040 2711.830 ;
        RECT 2525.100 2710.325 2525.240 2711.510 ;
        RECT 2525.030 2709.955 2525.310 2710.325 ;
      LAYER via2 ;
        RECT 2901.770 3196.880 2902.050 3197.160 ;
        RECT 2525.030 2710.000 2525.310 2710.280 ;
      LAYER met3 ;
        RECT 2901.745 3197.170 2902.075 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.745 3196.870 2924.800 3197.170 ;
        RECT 2901.745 3196.855 2902.075 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2506.000 2710.290 2510.000 2710.440 ;
        RECT 2525.005 2710.290 2525.335 2710.305 ;
        RECT 2506.000 2709.990 2525.335 2710.290 ;
        RECT 2506.000 2709.840 2510.000 2709.990 ;
        RECT 2525.005 2709.975 2525.335 2709.990 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2877.320 2525.330 2877.380 ;
        RECT 2901.290 2877.320 2901.610 2877.380 ;
        RECT 2525.010 2877.180 2901.610 2877.320 ;
        RECT 2525.010 2877.120 2525.330 2877.180 ;
        RECT 2901.290 2877.120 2901.610 2877.180 ;
      LAYER via ;
        RECT 2525.040 2877.120 2525.300 2877.380 ;
        RECT 2901.320 2877.120 2901.580 2877.380 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 2901.380 2877.410 2901.520 3431.435 ;
        RECT 2525.040 2877.090 2525.300 2877.410 ;
        RECT 2901.320 2877.090 2901.580 2877.410 ;
        RECT 2525.100 2873.525 2525.240 2877.090 ;
        RECT 2525.030 2873.155 2525.310 2873.525 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
        RECT 2525.030 2873.200 2525.310 2873.480 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2506.000 2873.490 2510.000 2873.640 ;
        RECT 2525.005 2873.490 2525.335 2873.505 ;
        RECT 2506.000 2873.190 2525.335 2873.490 ;
        RECT 2506.000 2873.040 2510.000 2873.190 ;
        RECT 2525.005 2873.175 2525.335 2873.190 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3415.555 ;
      LAYER mcon ;
        RECT 2713.685 3415.385 2713.855 3415.555 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2712.690 3470.620 2713.010 3470.680 ;
        RECT 2713.610 3470.620 2713.930 3470.680 ;
        RECT 2712.690 3470.480 2713.930 3470.620 ;
        RECT 2712.690 3470.420 2713.010 3470.480 ;
        RECT 2713.610 3470.420 2713.930 3470.480 ;
        RECT 2712.690 3463.820 2713.010 3463.880 ;
        RECT 2713.610 3463.820 2713.930 3463.880 ;
        RECT 2712.690 3463.680 2713.930 3463.820 ;
        RECT 2712.690 3463.620 2713.010 3463.680 ;
        RECT 2713.610 3463.620 2713.930 3463.680 ;
        RECT 2711.770 3415.540 2712.090 3415.600 ;
        RECT 2713.625 3415.540 2713.915 3415.585 ;
        RECT 2711.770 3415.400 2713.915 3415.540 ;
        RECT 2711.770 3415.340 2712.090 3415.400 ;
        RECT 2713.625 3415.355 2713.915 3415.400 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2407.710 3019.100 2408.030 3019.160 ;
        RECT 2712.230 3019.100 2712.550 3019.160 ;
        RECT 2407.710 3018.960 2712.550 3019.100 ;
        RECT 2407.710 3018.900 2408.030 3018.960 ;
        RECT 2712.230 3018.900 2712.550 3018.960 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2712.720 3470.420 2712.980 3470.680 ;
        RECT 2713.640 3470.420 2713.900 3470.680 ;
        RECT 2712.720 3463.620 2712.980 3463.880 ;
        RECT 2713.640 3463.620 2713.900 3463.880 ;
        RECT 2711.800 3415.340 2712.060 3415.600 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2407.740 3018.900 2408.000 3019.160 ;
        RECT 2712.260 3018.900 2712.520 3019.160 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3470.710 2713.840 3491.130 ;
        RECT 2712.720 3470.390 2712.980 3470.710 ;
        RECT 2713.640 3470.390 2713.900 3470.710 ;
        RECT 2712.780 3463.910 2712.920 3470.390 ;
        RECT 2712.720 3463.590 2712.980 3463.910 ;
        RECT 2713.640 3463.590 2713.900 3463.910 ;
        RECT 2713.700 3416.165 2713.840 3463.590 ;
        RECT 2711.790 3415.795 2712.070 3416.165 ;
        RECT 2713.630 3415.795 2713.910 3416.165 ;
        RECT 2711.860 3415.630 2712.000 3415.795 ;
        RECT 2711.800 3415.310 2712.060 3415.630 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3019.190 2712.460 3056.610 ;
        RECT 2407.740 3018.870 2408.000 3019.190 ;
        RECT 2712.260 3018.870 2712.520 3019.190 ;
        RECT 2407.800 3010.000 2407.940 3018.870 ;
        RECT 2407.800 3009.340 2408.150 3010.000 ;
        RECT 2407.870 3006.000 2408.150 3009.340 ;
      LAYER via2 ;
        RECT 2711.790 3415.840 2712.070 3416.120 ;
        RECT 2713.630 3415.840 2713.910 3416.120 ;
      LAYER met3 ;
        RECT 2711.765 3416.130 2712.095 3416.145 ;
        RECT 2713.605 3416.130 2713.935 3416.145 ;
        RECT 2711.765 3415.830 2713.935 3416.130 ;
        RECT 2711.765 3415.815 2712.095 3415.830 ;
        RECT 2713.605 3415.815 2713.935 3415.830 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.470 3464.160 2387.790 3464.220 ;
        RECT 2392.990 3464.160 2393.310 3464.220 ;
        RECT 2387.470 3464.020 2393.310 3464.160 ;
        RECT 2387.470 3463.960 2387.790 3464.020 ;
        RECT 2392.990 3463.960 2393.310 3464.020 ;
        RECT 2387.470 3367.600 2387.790 3367.660 ;
        RECT 2388.390 3367.600 2388.710 3367.660 ;
        RECT 2387.470 3367.460 2388.710 3367.600 ;
        RECT 2387.470 3367.400 2387.790 3367.460 ;
        RECT 2388.390 3367.400 2388.710 3367.460 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 2387.470 3077.580 2387.790 3077.640 ;
        RECT 2388.390 3077.580 2388.710 3077.640 ;
        RECT 2387.470 3077.440 2388.710 3077.580 ;
        RECT 2387.470 3077.380 2387.790 3077.440 ;
        RECT 2388.390 3077.380 2388.710 3077.440 ;
        RECT 2204.390 3019.100 2204.710 3019.160 ;
        RECT 2388.390 3019.100 2388.710 3019.160 ;
        RECT 2204.390 3018.960 2388.710 3019.100 ;
        RECT 2204.390 3018.900 2204.710 3018.960 ;
        RECT 2388.390 3018.900 2388.710 3018.960 ;
      LAYER via ;
        RECT 2387.500 3463.960 2387.760 3464.220 ;
        RECT 2393.020 3463.960 2393.280 3464.220 ;
        RECT 2387.500 3367.400 2387.760 3367.660 ;
        RECT 2388.420 3367.400 2388.680 3367.660 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 2387.500 3077.380 2387.760 3077.640 ;
        RECT 2388.420 3077.380 2388.680 3077.640 ;
        RECT 2204.420 3018.900 2204.680 3019.160 ;
        RECT 2388.420 3018.900 2388.680 3019.160 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3464.250 2393.220 3517.230 ;
        RECT 2387.500 3463.930 2387.760 3464.250 ;
        RECT 2393.020 3463.930 2393.280 3464.250 ;
        RECT 2387.560 3415.370 2387.700 3463.930 ;
        RECT 2387.560 3415.230 2388.620 3415.370 ;
        RECT 2388.480 3367.690 2388.620 3415.230 ;
        RECT 2387.500 3367.370 2387.760 3367.690 ;
        RECT 2388.420 3367.370 2388.680 3367.690 ;
        RECT 2387.560 3318.810 2387.700 3367.370 ;
        RECT 2387.560 3318.670 2388.620 3318.810 ;
        RECT 2388.480 3270.790 2388.620 3318.670 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 3019.190 2388.620 3028.990 ;
        RECT 2204.420 3018.870 2204.680 3019.190 ;
        RECT 2388.420 3018.870 2388.680 3019.190 ;
        RECT 2204.480 3010.000 2204.620 3018.870 ;
        RECT 2204.480 3009.340 2204.830 3010.000 ;
        RECT 2204.550 3006.000 2204.830 3009.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2063.245 3416.065 2063.415 3463.835 ;
        RECT 2065.085 3332.765 2065.255 3415.555 ;
      LAYER mcon ;
        RECT 2063.245 3463.665 2063.415 3463.835 ;
        RECT 2065.085 3415.385 2065.255 3415.555 ;
      LAYER met1 ;
        RECT 2065.010 3491.360 2065.330 3491.420 ;
        RECT 2068.690 3491.360 2069.010 3491.420 ;
        RECT 2065.010 3491.220 2069.010 3491.360 ;
        RECT 2065.010 3491.160 2065.330 3491.220 ;
        RECT 2068.690 3491.160 2069.010 3491.220 ;
        RECT 2064.090 3470.620 2064.410 3470.680 ;
        RECT 2065.010 3470.620 2065.330 3470.680 ;
        RECT 2064.090 3470.480 2065.330 3470.620 ;
        RECT 2064.090 3470.420 2064.410 3470.480 ;
        RECT 2065.010 3470.420 2065.330 3470.480 ;
        RECT 2063.185 3463.820 2063.475 3463.865 ;
        RECT 2064.090 3463.820 2064.410 3463.880 ;
        RECT 2063.185 3463.680 2064.410 3463.820 ;
        RECT 2063.185 3463.635 2063.475 3463.680 ;
        RECT 2064.090 3463.620 2064.410 3463.680 ;
        RECT 2063.170 3416.220 2063.490 3416.280 ;
        RECT 2063.170 3416.080 2063.685 3416.220 ;
        RECT 2063.170 3416.020 2063.490 3416.080 ;
        RECT 2063.170 3415.540 2063.490 3415.600 ;
        RECT 2065.025 3415.540 2065.315 3415.585 ;
        RECT 2063.170 3415.400 2065.315 3415.540 ;
        RECT 2063.170 3415.340 2063.490 3415.400 ;
        RECT 2065.025 3415.355 2065.315 3415.400 ;
        RECT 2065.025 3332.920 2065.315 3332.965 ;
        RECT 2065.470 3332.920 2065.790 3332.980 ;
        RECT 2065.025 3332.780 2065.790 3332.920 ;
        RECT 2065.025 3332.735 2065.315 3332.780 ;
        RECT 2065.470 3332.720 2065.790 3332.780 ;
        RECT 2064.090 3236.360 2064.410 3236.420 ;
        RECT 2064.550 3236.360 2064.870 3236.420 ;
        RECT 2064.090 3236.220 2064.870 3236.360 ;
        RECT 2064.090 3236.160 2064.410 3236.220 ;
        RECT 2064.550 3236.160 2064.870 3236.220 ;
        RECT 2064.090 3202.020 2064.410 3202.080 ;
        RECT 2064.550 3202.020 2064.870 3202.080 ;
        RECT 2064.090 3201.880 2064.870 3202.020 ;
        RECT 2064.090 3201.820 2064.410 3201.880 ;
        RECT 2064.550 3201.820 2064.870 3201.880 ;
        RECT 2063.630 3153.400 2063.950 3153.460 ;
        RECT 2064.550 3153.400 2064.870 3153.460 ;
        RECT 2063.630 3153.260 2064.870 3153.400 ;
        RECT 2063.630 3153.200 2063.950 3153.260 ;
        RECT 2064.550 3153.200 2064.870 3153.260 ;
        RECT 2063.630 3056.840 2063.950 3056.900 ;
        RECT 2064.550 3056.840 2064.870 3056.900 ;
        RECT 2063.630 3056.700 2064.870 3056.840 ;
        RECT 2063.630 3056.640 2063.950 3056.700 ;
        RECT 2064.550 3056.640 2064.870 3056.700 ;
        RECT 2001.070 3018.760 2001.390 3018.820 ;
        RECT 2063.630 3018.760 2063.950 3018.820 ;
        RECT 2001.070 3018.620 2063.950 3018.760 ;
        RECT 2001.070 3018.560 2001.390 3018.620 ;
        RECT 2063.630 3018.560 2063.950 3018.620 ;
      LAYER via ;
        RECT 2065.040 3491.160 2065.300 3491.420 ;
        RECT 2068.720 3491.160 2068.980 3491.420 ;
        RECT 2064.120 3470.420 2064.380 3470.680 ;
        RECT 2065.040 3470.420 2065.300 3470.680 ;
        RECT 2064.120 3463.620 2064.380 3463.880 ;
        RECT 2063.200 3416.020 2063.460 3416.280 ;
        RECT 2063.200 3415.340 2063.460 3415.600 ;
        RECT 2065.500 3332.720 2065.760 3332.980 ;
        RECT 2064.120 3236.160 2064.380 3236.420 ;
        RECT 2064.580 3236.160 2064.840 3236.420 ;
        RECT 2064.120 3201.820 2064.380 3202.080 ;
        RECT 2064.580 3201.820 2064.840 3202.080 ;
        RECT 2063.660 3153.200 2063.920 3153.460 ;
        RECT 2064.580 3153.200 2064.840 3153.460 ;
        RECT 2063.660 3056.640 2063.920 3056.900 ;
        RECT 2064.580 3056.640 2064.840 3056.900 ;
        RECT 2001.100 3018.560 2001.360 3018.820 ;
        RECT 2063.660 3018.560 2063.920 3018.820 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3470.710 2065.240 3491.130 ;
        RECT 2064.120 3470.390 2064.380 3470.710 ;
        RECT 2065.040 3470.390 2065.300 3470.710 ;
        RECT 2064.180 3463.910 2064.320 3470.390 ;
        RECT 2064.120 3463.590 2064.380 3463.910 ;
        RECT 2063.200 3415.990 2063.460 3416.310 ;
        RECT 2063.260 3415.630 2063.400 3415.990 ;
        RECT 2063.200 3415.310 2063.460 3415.630 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3018.850 2063.860 3056.610 ;
        RECT 2001.100 3018.530 2001.360 3018.850 ;
        RECT 2063.660 3018.530 2063.920 3018.850 ;
        RECT 2001.160 3010.000 2001.300 3018.530 ;
        RECT 2001.160 3009.340 2001.510 3010.000 ;
        RECT 2001.230 3006.000 2001.510 3009.340 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1743.545 3429.325 1743.715 3477.435 ;
        RECT 1743.545 3332.765 1743.715 3380.875 ;
        RECT 1744.925 3236.205 1745.095 3284.315 ;
        RECT 1744.005 3139.645 1744.175 3187.755 ;
      LAYER mcon ;
        RECT 1743.545 3477.265 1743.715 3477.435 ;
        RECT 1743.545 3380.705 1743.715 3380.875 ;
        RECT 1744.925 3284.145 1745.095 3284.315 ;
        RECT 1744.005 3187.585 1744.175 3187.755 ;
      LAYER met1 ;
        RECT 1743.470 3477.420 1743.790 3477.480 ;
        RECT 1743.275 3477.280 1743.790 3477.420 ;
        RECT 1743.470 3477.220 1743.790 3477.280 ;
        RECT 1743.485 3429.480 1743.775 3429.525 ;
        RECT 1743.930 3429.480 1744.250 3429.540 ;
        RECT 1743.485 3429.340 1744.250 3429.480 ;
        RECT 1743.485 3429.295 1743.775 3429.340 ;
        RECT 1743.930 3429.280 1744.250 3429.340 ;
        RECT 1743.470 3380.860 1743.790 3380.920 ;
        RECT 1743.275 3380.720 1743.790 3380.860 ;
        RECT 1743.470 3380.660 1743.790 3380.720 ;
        RECT 1743.485 3332.920 1743.775 3332.965 ;
        RECT 1743.930 3332.920 1744.250 3332.980 ;
        RECT 1743.485 3332.780 1744.250 3332.920 ;
        RECT 1743.485 3332.735 1743.775 3332.780 ;
        RECT 1743.930 3332.720 1744.250 3332.780 ;
        RECT 1744.390 3298.240 1744.710 3298.300 ;
        RECT 1745.310 3298.240 1745.630 3298.300 ;
        RECT 1744.390 3298.100 1745.630 3298.240 ;
        RECT 1744.390 3298.040 1744.710 3298.100 ;
        RECT 1745.310 3298.040 1745.630 3298.100 ;
        RECT 1744.865 3284.300 1745.155 3284.345 ;
        RECT 1745.310 3284.300 1745.630 3284.360 ;
        RECT 1744.865 3284.160 1745.630 3284.300 ;
        RECT 1744.865 3284.115 1745.155 3284.160 ;
        RECT 1745.310 3284.100 1745.630 3284.160 ;
        RECT 1744.850 3236.360 1745.170 3236.420 ;
        RECT 1744.655 3236.220 1745.170 3236.360 ;
        RECT 1744.850 3236.160 1745.170 3236.220 ;
        RECT 1744.850 3202.020 1745.170 3202.080 ;
        RECT 1744.020 3201.880 1745.170 3202.020 ;
        RECT 1744.020 3201.400 1744.160 3201.880 ;
        RECT 1744.850 3201.820 1745.170 3201.880 ;
        RECT 1743.930 3201.140 1744.250 3201.400 ;
        RECT 1743.930 3187.740 1744.250 3187.800 ;
        RECT 1743.735 3187.600 1744.250 3187.740 ;
        RECT 1743.930 3187.540 1744.250 3187.600 ;
        RECT 1743.945 3139.800 1744.235 3139.845 ;
        RECT 1745.310 3139.800 1745.630 3139.860 ;
        RECT 1743.945 3139.660 1745.630 3139.800 ;
        RECT 1743.945 3139.615 1744.235 3139.660 ;
        RECT 1745.310 3139.600 1745.630 3139.660 ;
        RECT 1745.310 3018.760 1745.630 3018.820 ;
        RECT 1798.210 3018.760 1798.530 3018.820 ;
        RECT 1745.310 3018.620 1798.530 3018.760 ;
        RECT 1745.310 3018.560 1745.630 3018.620 ;
        RECT 1798.210 3018.560 1798.530 3018.620 ;
      LAYER via ;
        RECT 1743.500 3477.220 1743.760 3477.480 ;
        RECT 1743.960 3429.280 1744.220 3429.540 ;
        RECT 1743.500 3380.660 1743.760 3380.920 ;
        RECT 1743.960 3332.720 1744.220 3332.980 ;
        RECT 1744.420 3298.040 1744.680 3298.300 ;
        RECT 1745.340 3298.040 1745.600 3298.300 ;
        RECT 1745.340 3284.100 1745.600 3284.360 ;
        RECT 1744.880 3236.160 1745.140 3236.420 ;
        RECT 1744.880 3201.820 1745.140 3202.080 ;
        RECT 1743.960 3201.140 1744.220 3201.400 ;
        RECT 1743.960 3187.540 1744.220 3187.800 ;
        RECT 1745.340 3139.600 1745.600 3139.860 ;
        RECT 1745.340 3018.560 1745.600 3018.820 ;
        RECT 1798.240 3018.560 1798.500 3018.820 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3517.370 1744.160 3517.600 ;
        RECT 1743.560 3517.230 1744.160 3517.370 ;
        RECT 1743.560 3477.510 1743.700 3517.230 ;
        RECT 1743.500 3477.190 1743.760 3477.510 ;
        RECT 1743.960 3429.250 1744.220 3429.570 ;
        RECT 1744.020 3394.970 1744.160 3429.250 ;
        RECT 1743.560 3394.830 1744.160 3394.970 ;
        RECT 1743.560 3380.950 1743.700 3394.830 ;
        RECT 1743.500 3380.630 1743.760 3380.950 ;
        RECT 1743.960 3332.690 1744.220 3333.010 ;
        RECT 1744.020 3298.410 1744.160 3332.690 ;
        RECT 1744.020 3298.330 1744.620 3298.410 ;
        RECT 1744.020 3298.270 1744.680 3298.330 ;
        RECT 1744.420 3298.010 1744.680 3298.270 ;
        RECT 1745.340 3298.010 1745.600 3298.330 ;
        RECT 1745.400 3284.390 1745.540 3298.010 ;
        RECT 1745.340 3284.070 1745.600 3284.390 ;
        RECT 1744.880 3236.130 1745.140 3236.450 ;
        RECT 1744.940 3202.110 1745.080 3236.130 ;
        RECT 1744.880 3201.790 1745.140 3202.110 ;
        RECT 1743.960 3201.110 1744.220 3201.430 ;
        RECT 1744.020 3187.830 1744.160 3201.110 ;
        RECT 1743.960 3187.510 1744.220 3187.830 ;
        RECT 1745.340 3139.570 1745.600 3139.890 ;
        RECT 1745.400 3018.850 1745.540 3139.570 ;
        RECT 1745.340 3018.530 1745.600 3018.850 ;
        RECT 1798.240 3018.530 1798.500 3018.850 ;
        RECT 1798.300 3010.000 1798.440 3018.530 ;
        RECT 1798.300 3009.340 1798.650 3010.000 ;
        RECT 1798.370 3006.000 1798.650 3009.340 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3270.700 1420.410 3270.760 ;
        RECT 1421.010 3270.700 1421.330 3270.760 ;
        RECT 1420.090 3270.560 1421.330 3270.700 ;
        RECT 1420.090 3270.500 1420.410 3270.560 ;
        RECT 1421.010 3270.500 1421.330 3270.560 ;
        RECT 1420.090 3174.140 1420.410 3174.200 ;
        RECT 1421.010 3174.140 1421.330 3174.200 ;
        RECT 1420.090 3174.000 1421.330 3174.140 ;
        RECT 1420.090 3173.940 1420.410 3174.000 ;
        RECT 1421.010 3173.940 1421.330 3174.000 ;
        RECT 1420.090 3077.580 1420.410 3077.640 ;
        RECT 1421.010 3077.580 1421.330 3077.640 ;
        RECT 1420.090 3077.440 1421.330 3077.580 ;
        RECT 1420.090 3077.380 1420.410 3077.440 ;
        RECT 1421.010 3077.380 1421.330 3077.440 ;
        RECT 1420.090 3019.100 1420.410 3019.160 ;
        RECT 1594.890 3019.100 1595.210 3019.160 ;
        RECT 1420.090 3018.960 1595.210 3019.100 ;
        RECT 1420.090 3018.900 1420.410 3018.960 ;
        RECT 1594.890 3018.900 1595.210 3018.960 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3270.500 1420.380 3270.760 ;
        RECT 1421.040 3270.500 1421.300 3270.760 ;
        RECT 1420.120 3173.940 1420.380 3174.200 ;
        RECT 1421.040 3173.940 1421.300 3174.200 ;
        RECT 1420.120 3077.380 1420.380 3077.640 ;
        RECT 1421.040 3077.380 1421.300 3077.640 ;
        RECT 1420.120 3018.900 1420.380 3019.160 ;
        RECT 1594.920 3018.900 1595.180 3019.160 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3222.250 1421.240 3270.470 ;
        RECT 1420.180 3222.110 1421.240 3222.250 ;
        RECT 1420.180 3174.230 1420.320 3222.110 ;
        RECT 1420.120 3173.910 1420.380 3174.230 ;
        RECT 1421.040 3173.910 1421.300 3174.230 ;
        RECT 1421.100 3125.690 1421.240 3173.910 ;
        RECT 1420.180 3125.550 1421.240 3125.690 ;
        RECT 1420.180 3077.670 1420.320 3125.550 ;
        RECT 1420.120 3077.350 1420.380 3077.670 ;
        RECT 1421.040 3077.350 1421.300 3077.670 ;
        RECT 1421.100 3029.130 1421.240 3077.350 ;
        RECT 1420.180 3028.990 1421.240 3029.130 ;
        RECT 1420.180 3019.190 1420.320 3028.990 ;
        RECT 1420.120 3018.870 1420.380 3019.190 ;
        RECT 1594.920 3018.870 1595.180 3019.190 ;
        RECT 1594.980 3010.000 1595.120 3018.870 ;
        RECT 1594.980 3009.340 1595.330 3010.000 ;
        RECT 1595.050 3006.000 1595.330 3009.340 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 386.140 2523.030 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2522.710 386.000 2901.150 386.140 ;
        RECT 2522.710 385.940 2523.030 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2522.740 385.940 2523.000 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2522.730 753.595 2523.010 753.965 ;
        RECT 2522.800 386.230 2522.940 753.595 ;
        RECT 2522.740 385.910 2523.000 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2522.730 753.640 2523.010 753.920 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2506.000 753.930 2510.000 754.080 ;
        RECT 2522.705 753.930 2523.035 753.945 ;
        RECT 2506.000 753.630 2523.035 753.930 ;
        RECT 2506.000 753.480 2510.000 753.630 ;
        RECT 2522.705 753.615 2523.035 753.630 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1095.405 3139.645 1095.575 3187.755 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1095.405 3187.585 1095.575 3187.755 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.135 3187.600 1095.650 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.345 3139.800 1095.635 3139.845 ;
        RECT 1096.710 3139.800 1097.030 3139.860 ;
        RECT 1095.345 3139.660 1097.030 3139.800 ;
        RECT 1095.345 3139.615 1095.635 3139.660 ;
        RECT 1096.710 3139.600 1097.030 3139.660 ;
        RECT 1096.710 3019.780 1097.030 3019.840 ;
        RECT 1391.570 3019.780 1391.890 3019.840 ;
        RECT 1096.710 3019.640 1391.890 3019.780 ;
        RECT 1096.710 3019.580 1097.030 3019.640 ;
        RECT 1391.570 3019.580 1391.890 3019.640 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1096.740 3139.600 1097.000 3139.860 ;
        RECT 1096.740 3019.580 1097.000 3019.840 ;
        RECT 1391.600 3019.580 1391.860 3019.840 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1096.740 3139.570 1097.000 3139.890 ;
        RECT 1096.800 3019.870 1096.940 3139.570 ;
        RECT 1096.740 3019.550 1097.000 3019.870 ;
        RECT 1391.600 3019.550 1391.860 3019.870 ;
        RECT 1391.660 3010.000 1391.800 3019.550 ;
        RECT 1391.660 3009.340 1392.010 3010.000 ;
        RECT 1391.730 3006.000 1392.010 3009.340 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 3018.760 771.810 3018.820 ;
        RECT 1188.250 3018.760 1188.570 3018.820 ;
        RECT 771.490 3018.620 1188.570 3018.760 ;
        RECT 771.490 3018.560 771.810 3018.620 ;
        RECT 1188.250 3018.560 1188.570 3018.620 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 3018.560 771.780 3018.820 ;
        RECT 1188.280 3018.560 1188.540 3018.820 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 3018.850 771.720 3028.990 ;
        RECT 771.520 3018.530 771.780 3018.850 ;
        RECT 1188.280 3018.530 1188.540 3018.850 ;
        RECT 1188.340 3010.000 1188.480 3018.530 ;
        RECT 1188.340 3009.340 1188.690 3010.000 ;
        RECT 1188.410 3006.000 1188.690 3009.340 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 3020.120 448.430 3020.180 ;
        RECT 985.390 3020.120 985.710 3020.180 ;
        RECT 448.110 3019.980 985.710 3020.120 ;
        RECT 448.110 3019.920 448.430 3019.980 ;
        RECT 985.390 3019.920 985.710 3019.980 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 3019.920 448.400 3020.180 ;
        RECT 985.420 3019.920 985.680 3020.180 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 3020.210 448.340 3498.270 ;
        RECT 448.140 3019.890 448.400 3020.210 ;
        RECT 985.420 3019.890 985.680 3020.210 ;
        RECT 985.480 3010.000 985.620 3019.890 ;
        RECT 985.480 3009.340 985.830 3010.000 ;
        RECT 985.550 3006.000 985.830 3009.340 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 3019.100 124.130 3019.160 ;
        RECT 782.070 3019.100 782.390 3019.160 ;
        RECT 123.810 3018.960 782.390 3019.100 ;
        RECT 123.810 3018.900 124.130 3018.960 ;
        RECT 782.070 3018.900 782.390 3018.960 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 3018.900 124.100 3019.160 ;
        RECT 782.100 3018.900 782.360 3019.160 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 3019.190 124.040 3498.270 ;
        RECT 123.840 3018.870 124.100 3019.190 ;
        RECT 782.100 3018.870 782.360 3019.190 ;
        RECT 782.160 3010.000 782.300 3018.870 ;
        RECT 782.160 3009.340 782.510 3010.000 ;
        RECT 782.230 3006.000 782.510 3009.340 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2925.600 17.410 2925.660 ;
        RECT 393.370 2925.600 393.690 2925.660 ;
        RECT 17.090 2925.460 393.690 2925.600 ;
        RECT 17.090 2925.400 17.410 2925.460 ;
        RECT 393.370 2925.400 393.690 2925.460 ;
      LAYER via ;
        RECT 17.120 2925.400 17.380 2925.660 ;
        RECT 393.400 2925.400 393.660 2925.660 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 2925.690 17.320 3339.635 ;
        RECT 17.120 2925.370 17.380 2925.690 ;
        RECT 393.400 2925.370 393.660 2925.690 ;
        RECT 393.460 2922.485 393.600 2925.370 ;
        RECT 393.390 2922.115 393.670 2922.485 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 393.390 2922.160 393.670 2922.440 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 393.365 2922.450 393.695 2922.465 ;
        RECT 410.000 2922.450 414.000 2922.600 ;
        RECT 393.365 2922.150 414.000 2922.450 ;
        RECT 393.365 2922.135 393.695 2922.150 ;
        RECT 410.000 2922.000 414.000 2922.150 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2752.880 17.870 2752.940 ;
        RECT 393.370 2752.880 393.690 2752.940 ;
        RECT 17.550 2752.740 393.690 2752.880 ;
        RECT 17.550 2752.680 17.870 2752.740 ;
        RECT 393.370 2752.680 393.690 2752.740 ;
      LAYER via ;
        RECT 17.580 2752.680 17.840 2752.940 ;
        RECT 393.400 2752.680 393.660 2752.940 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 2752.970 17.780 3051.995 ;
        RECT 17.580 2752.650 17.840 2752.970 ;
        RECT 393.400 2752.650 393.660 2752.970 ;
        RECT 393.460 2747.725 393.600 2752.650 ;
        RECT 393.390 2747.355 393.670 2747.725 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 393.390 2747.400 393.670 2747.680 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 393.365 2747.690 393.695 2747.705 ;
        RECT 410.000 2747.690 414.000 2747.840 ;
        RECT 393.365 2747.390 414.000 2747.690 ;
        RECT 393.365 2747.375 393.695 2747.390 ;
        RECT 410.000 2747.240 414.000 2747.390 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2573.700 17.410 2573.760 ;
        RECT 393.370 2573.700 393.690 2573.760 ;
        RECT 17.090 2573.560 393.690 2573.700 ;
        RECT 17.090 2573.500 17.410 2573.560 ;
        RECT 393.370 2573.500 393.690 2573.560 ;
      LAYER via ;
        RECT 17.120 2573.500 17.380 2573.760 ;
        RECT 393.400 2573.500 393.660 2573.760 ;
      LAYER met2 ;
        RECT 17.110 2765.035 17.390 2765.405 ;
        RECT 17.180 2573.790 17.320 2765.035 ;
        RECT 17.120 2573.470 17.380 2573.790 ;
        RECT 393.400 2573.645 393.660 2573.790 ;
        RECT 393.390 2573.275 393.670 2573.645 ;
      LAYER via2 ;
        RECT 17.110 2765.080 17.390 2765.360 ;
        RECT 393.390 2573.320 393.670 2573.600 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.085 2765.370 17.415 2765.385 ;
        RECT -4.800 2765.070 17.415 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.085 2765.055 17.415 2765.070 ;
        RECT 393.365 2573.610 393.695 2573.625 ;
        RECT 410.000 2573.610 414.000 2573.760 ;
        RECT 393.365 2573.310 414.000 2573.610 ;
        RECT 393.365 2573.295 393.695 2573.310 ;
        RECT 410.000 2573.160 414.000 2573.310 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2400.980 17.870 2401.040 ;
        RECT 393.370 2400.980 393.690 2401.040 ;
        RECT 17.550 2400.840 393.690 2400.980 ;
        RECT 17.550 2400.780 17.870 2400.840 ;
        RECT 393.370 2400.780 393.690 2400.840 ;
      LAYER via ;
        RECT 17.580 2400.780 17.840 2401.040 ;
        RECT 393.400 2400.780 393.660 2401.040 ;
      LAYER met2 ;
        RECT 17.570 2477.395 17.850 2477.765 ;
        RECT 17.640 2401.070 17.780 2477.395 ;
        RECT 17.580 2400.750 17.840 2401.070 ;
        RECT 393.400 2400.750 393.660 2401.070 ;
        RECT 393.460 2398.885 393.600 2400.750 ;
        RECT 393.390 2398.515 393.670 2398.885 ;
      LAYER via2 ;
        RECT 17.570 2477.440 17.850 2477.720 ;
        RECT 393.390 2398.560 393.670 2398.840 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.545 2477.730 17.875 2477.745 ;
        RECT -4.800 2477.430 17.875 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.545 2477.415 17.875 2477.430 ;
        RECT 393.365 2398.850 393.695 2398.865 ;
        RECT 410.000 2398.850 414.000 2399.000 ;
        RECT 393.365 2398.550 414.000 2398.850 ;
        RECT 393.365 2398.535 393.695 2398.550 ;
        RECT 410.000 2398.400 414.000 2398.550 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2194.260 16.030 2194.320 ;
        RECT 396.590 2194.260 396.910 2194.320 ;
        RECT 15.710 2194.120 396.910 2194.260 ;
        RECT 15.710 2194.060 16.030 2194.120 ;
        RECT 396.590 2194.060 396.910 2194.120 ;
      LAYER via ;
        RECT 15.740 2194.060 16.000 2194.320 ;
        RECT 396.620 2194.060 396.880 2194.320 ;
      LAYER met2 ;
        RECT 396.610 2224.435 396.890 2224.805 ;
        RECT 396.680 2194.350 396.820 2224.435 ;
        RECT 15.740 2194.030 16.000 2194.350 ;
        RECT 396.620 2194.030 396.880 2194.350 ;
        RECT 15.800 2190.125 15.940 2194.030 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 396.610 2224.480 396.890 2224.760 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT 396.585 2224.770 396.915 2224.785 ;
        RECT 410.000 2224.770 414.000 2224.920 ;
        RECT 396.585 2224.470 414.000 2224.770 ;
        RECT 396.585 2224.455 396.915 2224.470 ;
        RECT 410.000 2224.320 414.000 2224.470 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 397.510 1904.240 397.830 1904.300 ;
        RECT 16.170 1904.100 397.830 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 397.510 1904.040 397.830 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 397.540 1904.040 397.800 1904.300 ;
      LAYER met2 ;
        RECT 397.530 2049.675 397.810 2050.045 ;
        RECT 397.600 1904.330 397.740 2049.675 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 397.540 1904.010 397.800 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 397.530 2049.720 397.810 2050.000 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 397.505 2050.010 397.835 2050.025 ;
        RECT 410.000 2050.010 414.000 2050.160 ;
        RECT 397.505 2049.710 414.000 2050.010 ;
        RECT 397.505 2049.695 397.835 2049.710 ;
        RECT 410.000 2049.560 414.000 2049.710 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2524.090 620.740 2524.410 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2524.090 620.600 2901.150 620.740 ;
        RECT 2524.090 620.540 2524.410 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2524.120 620.540 2524.380 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2524.110 916.795 2524.390 917.165 ;
        RECT 2524.180 620.830 2524.320 916.795 ;
        RECT 2524.120 620.510 2524.380 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2524.110 916.840 2524.390 917.120 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2506.000 917.130 2510.000 917.280 ;
        RECT 2524.085 917.130 2524.415 917.145 ;
        RECT 2506.000 916.830 2524.415 917.130 ;
        RECT 2506.000 916.680 2510.000 916.830 ;
        RECT 2524.085 916.815 2524.415 916.830 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 398.430 1621.360 398.750 1621.420 ;
        RECT 16.170 1621.220 398.750 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 398.430 1621.160 398.750 1621.220 ;
      LAYER via ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 398.460 1621.160 398.720 1621.420 ;
      LAYER met2 ;
        RECT 398.450 1875.595 398.730 1875.965 ;
        RECT 398.520 1621.450 398.660 1875.595 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 398.460 1621.130 398.720 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 398.450 1875.640 398.730 1875.920 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 398.425 1875.930 398.755 1875.945 ;
        RECT 410.000 1875.930 414.000 1876.080 ;
        RECT 398.425 1875.630 414.000 1875.930 ;
        RECT 398.425 1875.615 398.755 1875.630 ;
        RECT 410.000 1875.480 414.000 1875.630 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 397.510 1400.700 397.830 1400.760 ;
        RECT 17.090 1400.560 397.830 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 397.510 1400.500 397.830 1400.560 ;
      LAYER via ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 397.540 1400.500 397.800 1400.760 ;
      LAYER met2 ;
        RECT 397.530 1700.835 397.810 1701.205 ;
        RECT 397.600 1400.790 397.740 1700.835 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 397.540 1400.470 397.800 1400.790 ;
      LAYER via2 ;
        RECT 397.530 1700.880 397.810 1701.160 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 397.505 1701.170 397.835 1701.185 ;
        RECT 410.000 1701.170 414.000 1701.320 ;
        RECT 397.505 1700.870 414.000 1701.170 ;
        RECT 397.505 1700.855 397.835 1700.870 ;
        RECT 410.000 1700.720 414.000 1700.870 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 396.590 1186.840 396.910 1186.900 ;
        RECT 17.090 1186.700 396.910 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 396.590 1186.640 396.910 1186.700 ;
      LAYER via ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 396.620 1186.640 396.880 1186.900 ;
      LAYER met2 ;
        RECT 396.610 1526.755 396.890 1527.125 ;
        RECT 396.680 1186.930 396.820 1526.755 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 396.620 1186.610 396.880 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 396.610 1526.800 396.890 1527.080 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 396.585 1527.090 396.915 1527.105 ;
        RECT 410.000 1527.090 414.000 1527.240 ;
        RECT 396.585 1526.790 414.000 1527.090 ;
        RECT 396.585 1526.775 396.915 1526.790 ;
        RECT 410.000 1526.640 414.000 1526.790 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 397.510 972.640 397.830 972.700 ;
        RECT 15.710 972.500 397.830 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 397.510 972.440 397.830 972.500 ;
      LAYER via ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 397.540 972.440 397.800 972.700 ;
      LAYER met2 ;
        RECT 397.530 1351.995 397.810 1352.365 ;
        RECT 397.600 972.730 397.740 1351.995 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 397.540 972.410 397.800 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 397.530 1352.040 397.810 1352.320 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 397.505 1352.330 397.835 1352.345 ;
        RECT 410.000 1352.330 414.000 1352.480 ;
        RECT 397.505 1352.030 414.000 1352.330 ;
        RECT 397.505 1352.015 397.835 1352.030 ;
        RECT 410.000 1351.880 414.000 1352.030 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 396.590 758.780 396.910 758.840 ;
        RECT 15.710 758.640 396.910 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 396.590 758.580 396.910 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 396.620 758.580 396.880 758.840 ;
      LAYER met2 ;
        RECT 396.610 1177.915 396.890 1178.285 ;
        RECT 396.680 758.870 396.820 1177.915 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 396.620 758.550 396.880 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 396.610 1177.960 396.890 1178.240 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 396.585 1178.250 396.915 1178.265 ;
        RECT 410.000 1178.250 414.000 1178.400 ;
        RECT 396.585 1177.950 414.000 1178.250 ;
        RECT 396.585 1177.935 396.915 1177.950 ;
        RECT 410.000 1177.800 414.000 1177.950 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 398.430 544.920 398.750 544.980 ;
        RECT 16.170 544.780 398.750 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 398.430 544.720 398.750 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 398.460 544.720 398.720 544.980 ;
      LAYER met2 ;
        RECT 398.450 1003.155 398.730 1003.525 ;
        RECT 398.520 545.010 398.660 1003.155 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 398.460 544.690 398.720 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 398.450 1003.200 398.730 1003.480 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 398.425 1003.490 398.755 1003.505 ;
        RECT 410.000 1003.490 414.000 1003.640 ;
        RECT 398.425 1003.190 414.000 1003.490 ;
        RECT 398.425 1003.175 398.755 1003.190 ;
        RECT 410.000 1003.040 414.000 1003.190 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 397.970 324.260 398.290 324.320 ;
        RECT 16.630 324.120 398.290 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 397.970 324.060 398.290 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 398.000 324.060 398.260 324.320 ;
      LAYER met2 ;
        RECT 397.990 829.075 398.270 829.445 ;
        RECT 398.060 324.350 398.200 829.075 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 398.000 324.030 398.260 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 397.990 829.120 398.270 829.400 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 397.965 829.410 398.295 829.425 ;
        RECT 410.000 829.410 414.000 829.560 ;
        RECT 397.965 829.110 414.000 829.410 ;
        RECT 397.965 829.095 398.295 829.110 ;
        RECT 410.000 828.960 414.000 829.110 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 397.050 110.400 397.370 110.460 ;
        RECT 15.710 110.260 397.370 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 397.050 110.200 397.370 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 397.080 110.200 397.340 110.460 ;
      LAYER met2 ;
        RECT 397.070 654.315 397.350 654.685 ;
        RECT 397.140 110.490 397.280 654.315 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 397.080 110.170 397.340 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 397.070 654.360 397.350 654.640 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 397.045 654.650 397.375 654.665 ;
        RECT 410.000 654.650 414.000 654.800 ;
        RECT 397.045 654.350 414.000 654.650 ;
        RECT 397.045 654.335 397.375 654.350 ;
        RECT 410.000 654.200 414.000 654.350 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 855.340 2523.030 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2522.710 855.200 2901.150 855.340 ;
        RECT 2522.710 855.140 2523.030 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2522.740 855.140 2523.000 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2522.730 1079.995 2523.010 1080.365 ;
        RECT 2522.800 855.430 2522.940 1079.995 ;
        RECT 2522.740 855.110 2523.000 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2522.730 1080.040 2523.010 1080.320 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2506.000 1080.330 2510.000 1080.480 ;
        RECT 2522.705 1080.330 2523.035 1080.345 ;
        RECT 2506.000 1080.030 2523.035 1080.330 ;
        RECT 2506.000 1079.880 2510.000 1080.030 ;
        RECT 2522.705 1080.015 2523.035 1080.030 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 1089.940 2522.570 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2522.250 1089.800 2901.150 1089.940 ;
        RECT 2522.250 1089.740 2522.570 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2522.280 1089.740 2522.540 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2522.270 1242.515 2522.550 1242.885 ;
        RECT 2522.340 1090.030 2522.480 1242.515 ;
        RECT 2522.280 1089.710 2522.540 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2522.270 1242.560 2522.550 1242.840 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2506.000 1242.850 2510.000 1243.000 ;
        RECT 2522.245 1242.850 2522.575 1242.865 ;
        RECT 2506.000 1242.550 2522.575 1242.850 ;
        RECT 2506.000 1242.400 2510.000 1242.550 ;
        RECT 2522.245 1242.535 2522.575 1242.550 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 1324.540 2522.570 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2522.250 1324.400 2901.150 1324.540 ;
        RECT 2522.250 1324.340 2522.570 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2522.280 1324.340 2522.540 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2522.270 1405.715 2522.550 1406.085 ;
        RECT 2522.340 1324.630 2522.480 1405.715 ;
        RECT 2522.280 1324.310 2522.540 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2522.270 1405.760 2522.550 1406.040 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2506.000 1406.050 2510.000 1406.200 ;
        RECT 2522.245 1406.050 2522.575 1406.065 ;
        RECT 2506.000 1405.750 2522.575 1406.050 ;
        RECT 2506.000 1405.600 2510.000 1405.750 ;
        RECT 2522.245 1405.735 2522.575 1405.750 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1559.140 2520.730 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2520.410 1559.000 2901.150 1559.140 ;
        RECT 2520.410 1558.940 2520.730 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2520.440 1558.940 2520.700 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2520.430 1568.915 2520.710 1569.285 ;
        RECT 2520.500 1559.230 2520.640 1568.915 ;
        RECT 2520.440 1558.910 2520.700 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2520.430 1568.960 2520.710 1569.240 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2506.000 1569.250 2510.000 1569.400 ;
        RECT 2520.405 1569.250 2520.735 1569.265 ;
        RECT 2506.000 1568.950 2520.735 1569.250 ;
        RECT 2506.000 1568.800 2510.000 1568.950 ;
        RECT 2520.405 1568.935 2520.735 1568.950 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1738.660 2525.330 1738.720 ;
        RECT 2901.750 1738.660 2902.070 1738.720 ;
        RECT 2525.010 1738.520 2902.070 1738.660 ;
        RECT 2525.010 1738.460 2525.330 1738.520 ;
        RECT 2901.750 1738.460 2902.070 1738.520 ;
      LAYER via ;
        RECT 2525.040 1738.460 2525.300 1738.720 ;
        RECT 2901.780 1738.460 2902.040 1738.720 ;
      LAYER met2 ;
        RECT 2901.770 1789.235 2902.050 1789.605 ;
        RECT 2901.840 1738.750 2901.980 1789.235 ;
        RECT 2525.040 1738.430 2525.300 1738.750 ;
        RECT 2901.780 1738.430 2902.040 1738.750 ;
        RECT 2525.100 1732.485 2525.240 1738.430 ;
        RECT 2525.030 1732.115 2525.310 1732.485 ;
      LAYER via2 ;
        RECT 2901.770 1789.280 2902.050 1789.560 ;
        RECT 2525.030 1732.160 2525.310 1732.440 ;
      LAYER met3 ;
        RECT 2901.745 1789.570 2902.075 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.745 1789.270 2924.800 1789.570 ;
        RECT 2901.745 1789.255 2902.075 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2506.000 1732.450 2510.000 1732.600 ;
        RECT 2525.005 1732.450 2525.335 1732.465 ;
        RECT 2506.000 1732.150 2525.335 1732.450 ;
        RECT 2506.000 1732.000 2510.000 1732.150 ;
        RECT 2525.005 1732.135 2525.335 1732.150 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1897.440 2519.810 1897.500 ;
        RECT 2901.290 1897.440 2901.610 1897.500 ;
        RECT 2519.490 1897.300 2901.610 1897.440 ;
        RECT 2519.490 1897.240 2519.810 1897.300 ;
        RECT 2901.290 1897.240 2901.610 1897.300 ;
      LAYER via ;
        RECT 2519.520 1897.240 2519.780 1897.500 ;
        RECT 2901.320 1897.240 2901.580 1897.500 ;
      LAYER met2 ;
        RECT 2901.310 2023.835 2901.590 2024.205 ;
        RECT 2901.380 1897.530 2901.520 2023.835 ;
        RECT 2519.520 1897.210 2519.780 1897.530 ;
        RECT 2901.320 1897.210 2901.580 1897.530 ;
        RECT 2519.580 1895.005 2519.720 1897.210 ;
        RECT 2519.510 1894.635 2519.790 1895.005 ;
      LAYER via2 ;
        RECT 2901.310 2023.880 2901.590 2024.160 ;
        RECT 2519.510 1894.680 2519.790 1894.960 ;
      LAYER met3 ;
        RECT 2901.285 2024.170 2901.615 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.285 2023.870 2924.800 2024.170 ;
        RECT 2901.285 2023.855 2901.615 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2506.000 1894.970 2510.000 1895.120 ;
        RECT 2519.485 1894.970 2519.815 1894.985 ;
        RECT 2506.000 1894.670 2519.815 1894.970 ;
        RECT 2506.000 1894.520 2510.000 1894.670 ;
        RECT 2519.485 1894.655 2519.815 1894.670 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 2063.020 2525.330 2063.080 ;
        RECT 2901.750 2063.020 2902.070 2063.080 ;
        RECT 2525.010 2062.880 2902.070 2063.020 ;
        RECT 2525.010 2062.820 2525.330 2062.880 ;
        RECT 2901.750 2062.820 2902.070 2062.880 ;
      LAYER via ;
        RECT 2525.040 2062.820 2525.300 2063.080 ;
        RECT 2901.780 2062.820 2902.040 2063.080 ;
      LAYER met2 ;
        RECT 2901.770 2258.435 2902.050 2258.805 ;
        RECT 2901.840 2063.110 2901.980 2258.435 ;
        RECT 2525.040 2062.790 2525.300 2063.110 ;
        RECT 2901.780 2062.790 2902.040 2063.110 ;
        RECT 2525.100 2058.205 2525.240 2062.790 ;
        RECT 2525.030 2057.835 2525.310 2058.205 ;
      LAYER via2 ;
        RECT 2901.770 2258.480 2902.050 2258.760 ;
        RECT 2525.030 2057.880 2525.310 2058.160 ;
      LAYER met3 ;
        RECT 2901.745 2258.770 2902.075 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2901.745 2258.470 2924.800 2258.770 ;
        RECT 2901.745 2258.455 2902.075 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2506.000 2058.170 2510.000 2058.320 ;
        RECT 2525.005 2058.170 2525.335 2058.185 ;
        RECT 2506.000 2057.870 2525.335 2058.170 ;
        RECT 2506.000 2057.720 2510.000 2057.870 ;
        RECT 2525.005 2057.855 2525.335 2057.870 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 24.040 633.350 24.100 ;
        RECT 862.570 24.040 862.890 24.100 ;
        RECT 633.030 23.900 862.890 24.040 ;
        RECT 633.030 23.840 633.350 23.900 ;
        RECT 862.570 23.840 862.890 23.900 ;
      LAYER via ;
        RECT 633.060 23.840 633.320 24.100 ;
        RECT 862.600 23.840 862.860 24.100 ;
      LAYER met2 ;
        RECT 864.110 510.410 864.390 514.000 ;
        RECT 862.660 510.270 864.390 510.410 ;
        RECT 862.660 24.130 862.800 510.270 ;
        RECT 864.110 510.000 864.390 510.270 ;
        RECT 633.060 23.810 633.320 24.130 ;
        RECT 862.600 23.810 862.860 24.130 ;
        RECT 633.120 2.400 633.260 23.810 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2144.205 338.045 2144.375 403.835 ;
        RECT 2144.205 241.485 2144.375 259.335 ;
        RECT 2145.125 138.465 2145.295 159.375 ;
        RECT 2144.665 23.885 2144.835 48.195 ;
      LAYER mcon ;
        RECT 2144.205 403.665 2144.375 403.835 ;
        RECT 2144.205 259.165 2144.375 259.335 ;
        RECT 2145.125 159.205 2145.295 159.375 ;
        RECT 2144.665 48.025 2144.835 48.195 ;
      LAYER met1 ;
        RECT 2144.130 476.240 2144.450 476.300 ;
        RECT 2145.050 476.240 2145.370 476.300 ;
        RECT 2144.130 476.100 2145.370 476.240 ;
        RECT 2144.130 476.040 2144.450 476.100 ;
        RECT 2145.050 476.040 2145.370 476.100 ;
        RECT 2144.130 427.960 2144.450 428.020 ;
        RECT 2144.590 427.960 2144.910 428.020 ;
        RECT 2144.130 427.820 2144.910 427.960 ;
        RECT 2144.130 427.760 2144.450 427.820 ;
        RECT 2144.590 427.760 2144.910 427.820 ;
        RECT 2143.210 403.820 2143.530 403.880 ;
        RECT 2144.145 403.820 2144.435 403.865 ;
        RECT 2143.210 403.680 2144.435 403.820 ;
        RECT 2143.210 403.620 2143.530 403.680 ;
        RECT 2144.145 403.635 2144.435 403.680 ;
        RECT 2144.145 338.200 2144.435 338.245 ;
        RECT 2144.590 338.200 2144.910 338.260 ;
        RECT 2144.145 338.060 2144.910 338.200 ;
        RECT 2144.145 338.015 2144.435 338.060 ;
        RECT 2144.590 338.000 2144.910 338.060 ;
        RECT 2144.145 259.320 2144.435 259.365 ;
        RECT 2145.050 259.320 2145.370 259.380 ;
        RECT 2144.145 259.180 2145.370 259.320 ;
        RECT 2144.145 259.135 2144.435 259.180 ;
        RECT 2145.050 259.120 2145.370 259.180 ;
        RECT 2144.130 241.640 2144.450 241.700 ;
        RECT 2143.935 241.500 2144.450 241.640 ;
        RECT 2144.130 241.440 2144.450 241.500 ;
        RECT 2145.050 159.360 2145.370 159.420 ;
        RECT 2144.855 159.220 2145.370 159.360 ;
        RECT 2145.050 159.160 2145.370 159.220 ;
        RECT 2145.050 138.620 2145.370 138.680 ;
        RECT 2144.855 138.480 2145.370 138.620 ;
        RECT 2145.050 138.420 2145.370 138.480 ;
        RECT 2143.670 137.940 2143.990 138.000 ;
        RECT 2145.050 137.940 2145.370 138.000 ;
        RECT 2143.670 137.800 2145.370 137.940 ;
        RECT 2143.670 137.740 2143.990 137.800 ;
        RECT 2145.050 137.740 2145.370 137.800 ;
        RECT 2144.590 48.180 2144.910 48.240 ;
        RECT 2144.395 48.040 2144.910 48.180 ;
        RECT 2144.590 47.980 2144.910 48.040 ;
        RECT 2144.605 24.040 2144.895 24.085 ;
        RECT 2417.370 24.040 2417.690 24.100 ;
        RECT 2144.605 23.900 2417.690 24.040 ;
        RECT 2144.605 23.855 2144.895 23.900 ;
        RECT 2417.370 23.840 2417.690 23.900 ;
      LAYER via ;
        RECT 2144.160 476.040 2144.420 476.300 ;
        RECT 2145.080 476.040 2145.340 476.300 ;
        RECT 2144.160 427.760 2144.420 428.020 ;
        RECT 2144.620 427.760 2144.880 428.020 ;
        RECT 2143.240 403.620 2143.500 403.880 ;
        RECT 2144.620 338.000 2144.880 338.260 ;
        RECT 2145.080 259.120 2145.340 259.380 ;
        RECT 2144.160 241.440 2144.420 241.700 ;
        RECT 2145.080 159.160 2145.340 159.420 ;
        RECT 2145.080 138.420 2145.340 138.680 ;
        RECT 2143.700 137.740 2143.960 138.000 ;
        RECT 2145.080 137.740 2145.340 138.000 ;
        RECT 2144.620 47.980 2144.880 48.240 ;
        RECT 2417.400 23.840 2417.660 24.100 ;
      LAYER met2 ;
        RECT 2144.750 510.410 2145.030 514.000 ;
        RECT 2144.220 510.270 2145.030 510.410 ;
        RECT 2144.220 476.330 2144.360 510.270 ;
        RECT 2144.750 510.000 2145.030 510.270 ;
        RECT 2144.160 476.010 2144.420 476.330 ;
        RECT 2145.080 476.010 2145.340 476.330 ;
        RECT 2145.140 475.730 2145.280 476.010 ;
        RECT 2144.220 475.590 2145.280 475.730 ;
        RECT 2144.220 428.050 2144.360 475.590 ;
        RECT 2144.160 427.730 2144.420 428.050 ;
        RECT 2144.620 427.730 2144.880 428.050 ;
        RECT 2144.680 427.565 2144.820 427.730 ;
        RECT 2143.230 427.195 2143.510 427.565 ;
        RECT 2144.610 427.195 2144.890 427.565 ;
        RECT 2143.300 403.910 2143.440 427.195 ;
        RECT 2143.240 403.590 2143.500 403.910 ;
        RECT 2144.620 337.970 2144.880 338.290 ;
        RECT 2144.680 303.690 2144.820 337.970 ;
        RECT 2144.680 303.550 2145.280 303.690 ;
        RECT 2145.140 259.410 2145.280 303.550 ;
        RECT 2145.080 259.090 2145.340 259.410 ;
        RECT 2144.160 241.410 2144.420 241.730 ;
        RECT 2144.220 207.130 2144.360 241.410 ;
        RECT 2144.220 206.990 2145.280 207.130 ;
        RECT 2145.140 159.450 2145.280 206.990 ;
        RECT 2145.080 159.130 2145.340 159.450 ;
        RECT 2145.080 138.390 2145.340 138.710 ;
        RECT 2145.140 138.030 2145.280 138.390 ;
        RECT 2143.700 137.710 2143.960 138.030 ;
        RECT 2145.080 137.710 2145.340 138.030 ;
        RECT 2143.760 71.810 2143.900 137.710 ;
        RECT 2143.760 71.670 2144.820 71.810 ;
        RECT 2144.680 48.270 2144.820 71.670 ;
        RECT 2144.620 47.950 2144.880 48.270 ;
        RECT 2417.400 23.810 2417.660 24.130 ;
        RECT 2417.460 2.400 2417.600 23.810 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 2143.230 427.240 2143.510 427.520 ;
        RECT 2144.610 427.240 2144.890 427.520 ;
      LAYER met3 ;
        RECT 2143.205 427.530 2143.535 427.545 ;
        RECT 2144.585 427.530 2144.915 427.545 ;
        RECT 2143.205 427.230 2144.915 427.530 ;
        RECT 2143.205 427.215 2143.535 427.230 ;
        RECT 2144.585 427.215 2144.915 427.230 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2157.010 500.040 2157.330 500.100 ;
        RECT 2418.290 500.040 2418.610 500.100 ;
        RECT 2157.010 499.900 2418.610 500.040 ;
        RECT 2157.010 499.840 2157.330 499.900 ;
        RECT 2418.290 499.840 2418.610 499.900 ;
        RECT 2418.290 20.980 2418.610 21.040 ;
        RECT 2434.850 20.980 2435.170 21.040 ;
        RECT 2418.290 20.840 2435.170 20.980 ;
        RECT 2418.290 20.780 2418.610 20.840 ;
        RECT 2434.850 20.780 2435.170 20.840 ;
      LAYER via ;
        RECT 2157.040 499.840 2157.300 500.100 ;
        RECT 2418.320 499.840 2418.580 500.100 ;
        RECT 2418.320 20.780 2418.580 21.040 ;
        RECT 2434.880 20.780 2435.140 21.040 ;
      LAYER met2 ;
        RECT 2157.170 510.340 2157.450 514.000 ;
        RECT 2157.100 510.000 2157.450 510.340 ;
        RECT 2157.100 500.130 2157.240 510.000 ;
        RECT 2157.040 499.810 2157.300 500.130 ;
        RECT 2418.320 499.810 2418.580 500.130 ;
        RECT 2418.380 21.070 2418.520 499.810 ;
        RECT 2418.320 20.750 2418.580 21.070 ;
        RECT 2434.880 20.750 2435.140 21.070 ;
        RECT 2434.940 2.400 2435.080 20.750 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.110 30.840 2173.430 30.900 ;
        RECT 2452.790 30.840 2453.110 30.900 ;
        RECT 2173.110 30.700 2453.110 30.840 ;
        RECT 2173.110 30.640 2173.430 30.700 ;
        RECT 2452.790 30.640 2453.110 30.700 ;
      LAYER via ;
        RECT 2173.140 30.640 2173.400 30.900 ;
        RECT 2452.820 30.640 2453.080 30.900 ;
      LAYER met2 ;
        RECT 2170.050 510.410 2170.330 514.000 ;
        RECT 2170.050 510.270 2173.340 510.410 ;
        RECT 2170.050 510.000 2170.330 510.270 ;
        RECT 2173.200 30.930 2173.340 510.270 ;
        RECT 2173.140 30.610 2173.400 30.930 ;
        RECT 2452.820 30.610 2453.080 30.930 ;
        RECT 2452.880 2.400 2453.020 30.610 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2182.770 496.980 2183.090 497.040 ;
        RECT 2190.590 496.980 2190.910 497.040 ;
        RECT 2182.770 496.840 2190.910 496.980 ;
        RECT 2182.770 496.780 2183.090 496.840 ;
        RECT 2190.590 496.780 2190.910 496.840 ;
        RECT 2190.590 37.980 2190.910 38.040 ;
        RECT 2470.730 37.980 2471.050 38.040 ;
        RECT 2190.590 37.840 2471.050 37.980 ;
        RECT 2190.590 37.780 2190.910 37.840 ;
        RECT 2470.730 37.780 2471.050 37.840 ;
      LAYER via ;
        RECT 2182.800 496.780 2183.060 497.040 ;
        RECT 2190.620 496.780 2190.880 497.040 ;
        RECT 2190.620 37.780 2190.880 38.040 ;
        RECT 2470.760 37.780 2471.020 38.040 ;
      LAYER met2 ;
        RECT 2182.930 510.340 2183.210 514.000 ;
        RECT 2182.860 510.000 2183.210 510.340 ;
        RECT 2182.860 497.070 2183.000 510.000 ;
        RECT 2182.800 496.750 2183.060 497.070 ;
        RECT 2190.620 496.750 2190.880 497.070 ;
        RECT 2190.680 38.070 2190.820 496.750 ;
        RECT 2190.620 37.750 2190.880 38.070 ;
        RECT 2470.760 37.750 2471.020 38.070 ;
        RECT 2470.820 2.400 2470.960 37.750 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2195.650 503.440 2195.970 503.500 ;
        RECT 2200.710 503.440 2201.030 503.500 ;
        RECT 2195.650 503.300 2201.030 503.440 ;
        RECT 2195.650 503.240 2195.970 503.300 ;
        RECT 2200.710 503.240 2201.030 503.300 ;
        RECT 2200.710 44.780 2201.030 44.840 ;
        RECT 2488.670 44.780 2488.990 44.840 ;
        RECT 2200.710 44.640 2488.990 44.780 ;
        RECT 2200.710 44.580 2201.030 44.640 ;
        RECT 2488.670 44.580 2488.990 44.640 ;
      LAYER via ;
        RECT 2195.680 503.240 2195.940 503.500 ;
        RECT 2200.740 503.240 2201.000 503.500 ;
        RECT 2200.740 44.580 2201.000 44.840 ;
        RECT 2488.700 44.580 2488.960 44.840 ;
      LAYER met2 ;
        RECT 2195.810 510.340 2196.090 514.000 ;
        RECT 2195.740 510.000 2196.090 510.340 ;
        RECT 2195.740 503.530 2195.880 510.000 ;
        RECT 2195.680 503.210 2195.940 503.530 ;
        RECT 2200.740 503.210 2201.000 503.530 ;
        RECT 2200.800 44.870 2200.940 503.210 ;
        RECT 2200.740 44.550 2201.000 44.870 ;
        RECT 2488.700 44.550 2488.960 44.870 ;
        RECT 2488.760 2.400 2488.900 44.550 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2208.530 493.240 2208.850 493.300 ;
        RECT 2504.770 493.240 2505.090 493.300 ;
        RECT 2208.530 493.100 2505.090 493.240 ;
        RECT 2208.530 493.040 2208.850 493.100 ;
        RECT 2504.770 493.040 2505.090 493.100 ;
      LAYER via ;
        RECT 2208.560 493.040 2208.820 493.300 ;
        RECT 2504.800 493.040 2505.060 493.300 ;
      LAYER met2 ;
        RECT 2208.690 510.340 2208.970 514.000 ;
        RECT 2208.620 510.000 2208.970 510.340 ;
        RECT 2208.620 493.330 2208.760 510.000 ;
        RECT 2208.560 493.010 2208.820 493.330 ;
        RECT 2504.800 493.010 2505.060 493.330 ;
        RECT 2504.860 3.130 2505.000 493.010 ;
        RECT 2504.860 2.990 2506.380 3.130 ;
        RECT 2506.240 2.400 2506.380 2.990 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2221.410 503.440 2221.730 503.500 ;
        RECT 2225.090 503.440 2225.410 503.500 ;
        RECT 2221.410 503.300 2225.410 503.440 ;
        RECT 2221.410 503.240 2221.730 503.300 ;
        RECT 2225.090 503.240 2225.410 503.300 ;
        RECT 2225.090 148.140 2225.410 148.200 ;
        RECT 2518.570 148.140 2518.890 148.200 ;
        RECT 2225.090 148.000 2518.890 148.140 ;
        RECT 2225.090 147.940 2225.410 148.000 ;
        RECT 2518.570 147.940 2518.890 148.000 ;
      LAYER via ;
        RECT 2221.440 503.240 2221.700 503.500 ;
        RECT 2225.120 503.240 2225.380 503.500 ;
        RECT 2225.120 147.940 2225.380 148.200 ;
        RECT 2518.600 147.940 2518.860 148.200 ;
      LAYER met2 ;
        RECT 2221.570 510.340 2221.850 514.000 ;
        RECT 2221.500 510.000 2221.850 510.340 ;
        RECT 2221.500 503.530 2221.640 510.000 ;
        RECT 2221.440 503.210 2221.700 503.530 ;
        RECT 2225.120 503.210 2225.380 503.530 ;
        RECT 2225.180 148.230 2225.320 503.210 ;
        RECT 2225.120 147.910 2225.380 148.230 ;
        RECT 2518.600 147.910 2518.860 148.230 ;
        RECT 2518.660 16.730 2518.800 147.910 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2235.210 51.580 2235.530 51.640 ;
        RECT 2539.270 51.580 2539.590 51.640 ;
        RECT 2235.210 51.440 2539.590 51.580 ;
        RECT 2235.210 51.380 2235.530 51.440 ;
        RECT 2539.270 51.380 2539.590 51.440 ;
      LAYER via ;
        RECT 2235.240 51.380 2235.500 51.640 ;
        RECT 2539.300 51.380 2539.560 51.640 ;
      LAYER met2 ;
        RECT 2233.990 510.410 2234.270 514.000 ;
        RECT 2233.990 510.270 2235.440 510.410 ;
        RECT 2233.990 510.000 2234.270 510.270 ;
        RECT 2235.300 51.670 2235.440 510.270 ;
        RECT 2235.240 51.350 2235.500 51.670 ;
        RECT 2539.300 51.350 2539.560 51.670 ;
        RECT 2539.360 16.730 2539.500 51.350 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.400 2542.260 16.590 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2249.010 58.720 2249.330 58.780 ;
        RECT 2560.430 58.720 2560.750 58.780 ;
        RECT 2249.010 58.580 2560.750 58.720 ;
        RECT 2249.010 58.520 2249.330 58.580 ;
        RECT 2560.430 58.520 2560.750 58.580 ;
      LAYER via ;
        RECT 2249.040 58.520 2249.300 58.780 ;
        RECT 2560.460 58.520 2560.720 58.780 ;
      LAYER met2 ;
        RECT 2246.870 510.410 2247.150 514.000 ;
        RECT 2246.870 510.270 2249.240 510.410 ;
        RECT 2246.870 510.000 2247.150 510.270 ;
        RECT 2249.100 58.810 2249.240 510.270 ;
        RECT 2249.040 58.490 2249.300 58.810 ;
        RECT 2560.460 58.490 2560.720 58.810 ;
        RECT 2560.520 7.210 2560.660 58.490 ;
        RECT 2560.060 7.070 2560.660 7.210 ;
        RECT 2560.060 2.400 2560.200 7.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2262.810 65.520 2263.130 65.580 ;
        RECT 2573.770 65.520 2574.090 65.580 ;
        RECT 2262.810 65.380 2574.090 65.520 ;
        RECT 2262.810 65.320 2263.130 65.380 ;
        RECT 2573.770 65.320 2574.090 65.380 ;
      LAYER via ;
        RECT 2262.840 65.320 2263.100 65.580 ;
        RECT 2573.800 65.320 2574.060 65.580 ;
      LAYER met2 ;
        RECT 2259.750 510.410 2260.030 514.000 ;
        RECT 2259.750 510.270 2263.040 510.410 ;
        RECT 2259.750 510.000 2260.030 510.270 ;
        RECT 2262.900 65.610 2263.040 510.270 ;
        RECT 2262.840 65.290 2263.100 65.610 ;
        RECT 2573.800 65.290 2574.060 65.610 ;
        RECT 2573.860 17.410 2574.000 65.290 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.770 472.840 987.090 472.900 ;
        RECT 989.990 472.840 990.310 472.900 ;
        RECT 986.770 472.700 990.310 472.840 ;
        RECT 986.770 472.640 987.090 472.700 ;
        RECT 989.990 472.640 990.310 472.700 ;
        RECT 811.510 30.840 811.830 30.900 ;
        RECT 986.770 30.840 987.090 30.900 ;
        RECT 811.510 30.700 987.090 30.840 ;
        RECT 811.510 30.640 811.830 30.700 ;
        RECT 986.770 30.640 987.090 30.700 ;
      LAYER via ;
        RECT 986.800 472.640 987.060 472.900 ;
        RECT 990.020 472.640 990.280 472.900 ;
        RECT 811.540 30.640 811.800 30.900 ;
        RECT 986.800 30.640 987.060 30.900 ;
      LAYER met2 ;
        RECT 991.990 510.410 992.270 514.000 ;
        RECT 990.080 510.270 992.270 510.410 ;
        RECT 990.080 472.930 990.220 510.270 ;
        RECT 991.990 510.000 992.270 510.270 ;
        RECT 986.800 472.610 987.060 472.930 ;
        RECT 990.020 472.610 990.280 472.930 ;
        RECT 986.860 30.930 987.000 472.610 ;
        RECT 811.540 30.610 811.800 30.930 ;
        RECT 986.800 30.610 987.060 30.930 ;
        RECT 811.600 2.400 811.740 30.610 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2272.470 486.440 2272.790 486.500 ;
        RECT 2594.470 486.440 2594.790 486.500 ;
        RECT 2272.470 486.300 2594.790 486.440 ;
        RECT 2272.470 486.240 2272.790 486.300 ;
        RECT 2594.470 486.240 2594.790 486.300 ;
      LAYER via ;
        RECT 2272.500 486.240 2272.760 486.500 ;
        RECT 2594.500 486.240 2594.760 486.500 ;
      LAYER met2 ;
        RECT 2272.630 510.340 2272.910 514.000 ;
        RECT 2272.560 510.000 2272.910 510.340 ;
        RECT 2272.560 486.530 2272.700 510.000 ;
        RECT 2272.500 486.210 2272.760 486.530 ;
        RECT 2594.500 486.210 2594.760 486.530 ;
        RECT 2594.560 17.410 2594.700 486.210 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2285.350 479.640 2285.670 479.700 ;
        RECT 2608.270 479.640 2608.590 479.700 ;
        RECT 2285.350 479.500 2608.590 479.640 ;
        RECT 2285.350 479.440 2285.670 479.500 ;
        RECT 2608.270 479.440 2608.590 479.500 ;
      LAYER via ;
        RECT 2285.380 479.440 2285.640 479.700 ;
        RECT 2608.300 479.440 2608.560 479.700 ;
      LAYER met2 ;
        RECT 2285.510 510.340 2285.790 514.000 ;
        RECT 2285.440 510.000 2285.790 510.340 ;
        RECT 2285.440 479.730 2285.580 510.000 ;
        RECT 2285.380 479.410 2285.640 479.730 ;
        RECT 2608.300 479.410 2608.560 479.730 ;
        RECT 2608.360 17.410 2608.500 479.410 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2298.230 496.980 2298.550 497.040 ;
        RECT 2304.210 496.980 2304.530 497.040 ;
        RECT 2298.230 496.840 2304.530 496.980 ;
        RECT 2298.230 496.780 2298.550 496.840 ;
        RECT 2304.210 496.780 2304.530 496.840 ;
        RECT 2304.210 72.320 2304.530 72.380 ;
        RECT 2628.970 72.320 2629.290 72.380 ;
        RECT 2304.210 72.180 2629.290 72.320 ;
        RECT 2304.210 72.120 2304.530 72.180 ;
        RECT 2628.970 72.120 2629.290 72.180 ;
      LAYER via ;
        RECT 2298.260 496.780 2298.520 497.040 ;
        RECT 2304.240 496.780 2304.500 497.040 ;
        RECT 2304.240 72.120 2304.500 72.380 ;
        RECT 2629.000 72.120 2629.260 72.380 ;
      LAYER met2 ;
        RECT 2298.390 510.340 2298.670 514.000 ;
        RECT 2298.320 510.000 2298.670 510.340 ;
        RECT 2298.320 497.070 2298.460 510.000 ;
        RECT 2298.260 496.750 2298.520 497.070 ;
        RECT 2304.240 496.750 2304.500 497.070 ;
        RECT 2304.300 72.410 2304.440 496.750 ;
        RECT 2304.240 72.090 2304.500 72.410 ;
        RECT 2629.000 72.090 2629.260 72.410 ;
        RECT 2629.060 17.410 2629.200 72.090 ;
        RECT 2629.060 17.270 2631.500 17.410 ;
        RECT 2631.360 2.400 2631.500 17.270 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2312.030 472.500 2312.350 472.560 ;
        RECT 2642.770 472.500 2643.090 472.560 ;
        RECT 2312.030 472.360 2643.090 472.500 ;
        RECT 2312.030 472.300 2312.350 472.360 ;
        RECT 2642.770 472.300 2643.090 472.360 ;
        RECT 2642.770 16.900 2643.090 16.960 ;
        RECT 2649.210 16.900 2649.530 16.960 ;
        RECT 2642.770 16.760 2649.530 16.900 ;
        RECT 2642.770 16.700 2643.090 16.760 ;
        RECT 2649.210 16.700 2649.530 16.760 ;
      LAYER via ;
        RECT 2312.060 472.300 2312.320 472.560 ;
        RECT 2642.800 472.300 2643.060 472.560 ;
        RECT 2642.800 16.700 2643.060 16.960 ;
        RECT 2649.240 16.700 2649.500 16.960 ;
      LAYER met2 ;
        RECT 2310.810 510.340 2311.090 514.000 ;
        RECT 2310.740 510.000 2311.090 510.340 ;
        RECT 2310.740 497.490 2310.880 510.000 ;
        RECT 2310.740 497.350 2312.260 497.490 ;
        RECT 2312.120 472.590 2312.260 497.350 ;
        RECT 2312.060 472.270 2312.320 472.590 ;
        RECT 2642.800 472.270 2643.060 472.590 ;
        RECT 2642.860 16.990 2643.000 472.270 ;
        RECT 2642.800 16.670 2643.060 16.990 ;
        RECT 2649.240 16.670 2649.500 16.990 ;
        RECT 2649.300 2.400 2649.440 16.670 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2324.910 79.460 2325.230 79.520 ;
        RECT 2663.470 79.460 2663.790 79.520 ;
        RECT 2324.910 79.320 2663.790 79.460 ;
        RECT 2324.910 79.260 2325.230 79.320 ;
        RECT 2663.470 79.260 2663.790 79.320 ;
      LAYER via ;
        RECT 2324.940 79.260 2325.200 79.520 ;
        RECT 2663.500 79.260 2663.760 79.520 ;
      LAYER met2 ;
        RECT 2323.690 510.410 2323.970 514.000 ;
        RECT 2323.690 510.270 2325.140 510.410 ;
        RECT 2323.690 510.000 2323.970 510.270 ;
        RECT 2325.000 79.550 2325.140 510.270 ;
        RECT 2324.940 79.230 2325.200 79.550 ;
        RECT 2663.500 79.230 2663.760 79.550 ;
        RECT 2663.560 17.410 2663.700 79.230 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2338.250 465.700 2338.570 465.760 ;
        RECT 2684.170 465.700 2684.490 465.760 ;
        RECT 2338.250 465.560 2684.490 465.700 ;
        RECT 2338.250 465.500 2338.570 465.560 ;
        RECT 2684.170 465.500 2684.490 465.560 ;
      LAYER via ;
        RECT 2338.280 465.500 2338.540 465.760 ;
        RECT 2684.200 465.500 2684.460 465.760 ;
      LAYER met2 ;
        RECT 2336.570 510.410 2336.850 514.000 ;
        RECT 2336.570 510.270 2338.480 510.410 ;
        RECT 2336.570 510.000 2336.850 510.270 ;
        RECT 2338.340 465.790 2338.480 510.270 ;
        RECT 2338.280 465.470 2338.540 465.790 ;
        RECT 2684.200 465.470 2684.460 465.790 ;
        RECT 2684.260 17.410 2684.400 465.470 ;
        RECT 2684.260 17.270 2684.860 17.410 ;
        RECT 2684.720 2.400 2684.860 17.270 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2352.510 120.600 2352.830 120.660 ;
        RECT 2697.970 120.600 2698.290 120.660 ;
        RECT 2352.510 120.460 2698.290 120.600 ;
        RECT 2352.510 120.400 2352.830 120.460 ;
        RECT 2697.970 120.400 2698.290 120.460 ;
      LAYER via ;
        RECT 2352.540 120.400 2352.800 120.660 ;
        RECT 2698.000 120.400 2698.260 120.660 ;
      LAYER met2 ;
        RECT 2349.450 510.410 2349.730 514.000 ;
        RECT 2349.450 510.270 2352.740 510.410 ;
        RECT 2349.450 510.000 2349.730 510.270 ;
        RECT 2352.600 120.690 2352.740 510.270 ;
        RECT 2352.540 120.370 2352.800 120.690 ;
        RECT 2698.000 120.370 2698.260 120.690 ;
        RECT 2698.060 16.730 2698.200 120.370 ;
        RECT 2698.060 16.590 2702.800 16.730 ;
        RECT 2702.660 2.400 2702.800 16.590 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2362.170 500.380 2362.490 500.440 ;
        RECT 2535.590 500.380 2535.910 500.440 ;
        RECT 2362.170 500.240 2535.910 500.380 ;
        RECT 2362.170 500.180 2362.490 500.240 ;
        RECT 2535.590 500.180 2535.910 500.240 ;
        RECT 2535.590 24.040 2535.910 24.100 ;
        RECT 2720.510 24.040 2720.830 24.100 ;
        RECT 2535.590 23.900 2720.830 24.040 ;
        RECT 2535.590 23.840 2535.910 23.900 ;
        RECT 2720.510 23.840 2720.830 23.900 ;
      LAYER via ;
        RECT 2362.200 500.180 2362.460 500.440 ;
        RECT 2535.620 500.180 2535.880 500.440 ;
        RECT 2535.620 23.840 2535.880 24.100 ;
        RECT 2720.540 23.840 2720.800 24.100 ;
      LAYER met2 ;
        RECT 2362.330 510.340 2362.610 514.000 ;
        RECT 2362.260 510.000 2362.610 510.340 ;
        RECT 2362.260 500.470 2362.400 510.000 ;
        RECT 2362.200 500.150 2362.460 500.470 ;
        RECT 2535.620 500.150 2535.880 500.470 ;
        RECT 2535.680 24.130 2535.820 500.150 ;
        RECT 2535.620 23.810 2535.880 24.130 ;
        RECT 2720.540 23.810 2720.800 24.130 ;
        RECT 2720.600 2.400 2720.740 23.810 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2375.050 503.440 2375.370 503.500 ;
        RECT 2379.650 503.440 2379.970 503.500 ;
        RECT 2375.050 503.300 2379.970 503.440 ;
        RECT 2375.050 503.240 2375.370 503.300 ;
        RECT 2379.650 503.240 2379.970 503.300 ;
        RECT 2379.650 458.900 2379.970 458.960 ;
        RECT 2732.930 458.900 2733.250 458.960 ;
        RECT 2379.650 458.760 2733.250 458.900 ;
        RECT 2379.650 458.700 2379.970 458.760 ;
        RECT 2732.930 458.700 2733.250 458.760 ;
      LAYER via ;
        RECT 2375.080 503.240 2375.340 503.500 ;
        RECT 2379.680 503.240 2379.940 503.500 ;
        RECT 2379.680 458.700 2379.940 458.960 ;
        RECT 2732.960 458.700 2733.220 458.960 ;
      LAYER met2 ;
        RECT 2375.210 510.340 2375.490 514.000 ;
        RECT 2375.140 510.000 2375.490 510.340 ;
        RECT 2375.140 503.530 2375.280 510.000 ;
        RECT 2375.080 503.210 2375.340 503.530 ;
        RECT 2379.680 503.210 2379.940 503.530 ;
        RECT 2379.740 458.990 2379.880 503.210 ;
        RECT 2379.680 458.670 2379.940 458.990 ;
        RECT 2732.960 458.670 2733.220 458.990 ;
        RECT 2733.020 16.730 2733.160 458.670 ;
        RECT 2733.020 16.590 2738.680 16.730 ;
        RECT 2738.540 2.400 2738.680 16.590 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.470 496.980 2387.790 497.040 ;
        RECT 2393.910 496.980 2394.230 497.040 ;
        RECT 2387.470 496.840 2394.230 496.980 ;
        RECT 2387.470 496.780 2387.790 496.840 ;
        RECT 2393.910 496.780 2394.230 496.840 ;
        RECT 2393.910 93.060 2394.230 93.120 ;
        RECT 2753.170 93.060 2753.490 93.120 ;
        RECT 2393.910 92.920 2753.490 93.060 ;
        RECT 2393.910 92.860 2394.230 92.920 ;
        RECT 2753.170 92.860 2753.490 92.920 ;
      LAYER via ;
        RECT 2387.500 496.780 2387.760 497.040 ;
        RECT 2393.940 496.780 2394.200 497.040 ;
        RECT 2393.940 92.860 2394.200 93.120 ;
        RECT 2753.200 92.860 2753.460 93.120 ;
      LAYER met2 ;
        RECT 2387.630 510.340 2387.910 514.000 ;
        RECT 2387.560 510.000 2387.910 510.340 ;
        RECT 2387.560 497.070 2387.700 510.000 ;
        RECT 2387.500 496.750 2387.760 497.070 ;
        RECT 2393.940 496.750 2394.200 497.070 ;
        RECT 2394.000 93.150 2394.140 496.750 ;
        RECT 2393.940 92.830 2394.200 93.150 ;
        RECT 2753.200 92.830 2753.460 93.150 ;
        RECT 2753.260 17.410 2753.400 92.830 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 838.190 500.380 838.510 500.440 ;
        RECT 1004.710 500.380 1005.030 500.440 ;
        RECT 838.190 500.240 1005.030 500.380 ;
        RECT 838.190 500.180 838.510 500.240 ;
        RECT 1004.710 500.180 1005.030 500.240 ;
        RECT 829.450 24.380 829.770 24.440 ;
        RECT 838.190 24.380 838.510 24.440 ;
        RECT 829.450 24.240 838.510 24.380 ;
        RECT 829.450 24.180 829.770 24.240 ;
        RECT 838.190 24.180 838.510 24.240 ;
      LAYER via ;
        RECT 838.220 500.180 838.480 500.440 ;
        RECT 1004.740 500.180 1005.000 500.440 ;
        RECT 829.480 24.180 829.740 24.440 ;
        RECT 838.220 24.180 838.480 24.440 ;
      LAYER met2 ;
        RECT 1004.870 510.340 1005.150 514.000 ;
        RECT 1004.800 510.000 1005.150 510.340 ;
        RECT 1004.800 500.470 1004.940 510.000 ;
        RECT 838.220 500.150 838.480 500.470 ;
        RECT 1004.740 500.150 1005.000 500.470 ;
        RECT 838.280 24.470 838.420 500.150 ;
        RECT 829.480 24.150 829.740 24.470 ;
        RECT 838.220 24.150 838.480 24.470 ;
        RECT 829.540 2.400 829.680 24.150 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.350 451.760 2400.670 451.820 ;
        RECT 2773.870 451.760 2774.190 451.820 ;
        RECT 2400.350 451.620 2774.190 451.760 ;
        RECT 2400.350 451.560 2400.670 451.620 ;
        RECT 2773.870 451.560 2774.190 451.620 ;
      LAYER via ;
        RECT 2400.380 451.560 2400.640 451.820 ;
        RECT 2773.900 451.560 2774.160 451.820 ;
      LAYER met2 ;
        RECT 2400.510 510.340 2400.790 514.000 ;
        RECT 2400.440 510.000 2400.790 510.340 ;
        RECT 2400.440 451.850 2400.580 510.000 ;
        RECT 2400.380 451.530 2400.640 451.850 ;
        RECT 2773.900 451.530 2774.160 451.850 ;
        RECT 2773.960 2.400 2774.100 451.530 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2414.150 444.960 2414.470 445.020 ;
        RECT 2787.670 444.960 2787.990 445.020 ;
        RECT 2414.150 444.820 2787.990 444.960 ;
        RECT 2414.150 444.760 2414.470 444.820 ;
        RECT 2787.670 444.760 2787.990 444.820 ;
      LAYER via ;
        RECT 2414.180 444.760 2414.440 445.020 ;
        RECT 2787.700 444.760 2787.960 445.020 ;
      LAYER met2 ;
        RECT 2413.390 510.410 2413.670 514.000 ;
        RECT 2413.390 510.270 2414.380 510.410 ;
        RECT 2413.390 510.000 2413.670 510.270 ;
        RECT 2414.240 445.050 2414.380 510.270 ;
        RECT 2414.180 444.730 2414.440 445.050 ;
        RECT 2787.700 444.730 2787.960 445.050 ;
        RECT 2787.760 17.410 2787.900 444.730 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2426.110 500.720 2426.430 500.780 ;
        RECT 2514.890 500.720 2515.210 500.780 ;
        RECT 2426.110 500.580 2515.210 500.720 ;
        RECT 2426.110 500.520 2426.430 500.580 ;
        RECT 2514.890 500.520 2515.210 500.580 ;
        RECT 2514.890 30.840 2515.210 30.900 ;
        RECT 2809.750 30.840 2810.070 30.900 ;
        RECT 2514.890 30.700 2810.070 30.840 ;
        RECT 2514.890 30.640 2515.210 30.700 ;
        RECT 2809.750 30.640 2810.070 30.700 ;
      LAYER via ;
        RECT 2426.140 500.520 2426.400 500.780 ;
        RECT 2514.920 500.520 2515.180 500.780 ;
        RECT 2514.920 30.640 2515.180 30.900 ;
        RECT 2809.780 30.640 2810.040 30.900 ;
      LAYER met2 ;
        RECT 2426.270 510.340 2426.550 514.000 ;
        RECT 2426.200 510.000 2426.550 510.340 ;
        RECT 2426.200 500.810 2426.340 510.000 ;
        RECT 2426.140 500.490 2426.400 500.810 ;
        RECT 2514.920 500.490 2515.180 500.810 ;
        RECT 2514.980 30.930 2515.120 500.490 ;
        RECT 2514.920 30.610 2515.180 30.930 ;
        RECT 2809.780 30.610 2810.040 30.930 ;
        RECT 2809.840 2.400 2809.980 30.610 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2442.210 134.540 2442.530 134.600 ;
        RECT 2822.170 134.540 2822.490 134.600 ;
        RECT 2442.210 134.400 2822.490 134.540 ;
        RECT 2442.210 134.340 2442.530 134.400 ;
        RECT 2822.170 134.340 2822.490 134.400 ;
      LAYER via ;
        RECT 2442.240 134.340 2442.500 134.600 ;
        RECT 2822.200 134.340 2822.460 134.600 ;
      LAYER met2 ;
        RECT 2439.150 510.410 2439.430 514.000 ;
        RECT 2439.150 510.270 2442.440 510.410 ;
        RECT 2439.150 510.000 2439.430 510.270 ;
        RECT 2442.300 134.630 2442.440 510.270 ;
        RECT 2442.240 134.310 2442.500 134.630 ;
        RECT 2822.200 134.310 2822.460 134.630 ;
        RECT 2822.260 17.410 2822.400 134.310 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2451.870 496.980 2452.190 497.040 ;
        RECT 2459.690 496.980 2460.010 497.040 ;
        RECT 2451.870 496.840 2460.010 496.980 ;
        RECT 2451.870 496.780 2452.190 496.840 ;
        RECT 2459.690 496.780 2460.010 496.840 ;
        RECT 2459.690 431.360 2460.010 431.420 ;
        RECT 2842.870 431.360 2843.190 431.420 ;
        RECT 2459.690 431.220 2843.190 431.360 ;
        RECT 2459.690 431.160 2460.010 431.220 ;
        RECT 2842.870 431.160 2843.190 431.220 ;
      LAYER via ;
        RECT 2451.900 496.780 2452.160 497.040 ;
        RECT 2459.720 496.780 2459.980 497.040 ;
        RECT 2459.720 431.160 2459.980 431.420 ;
        RECT 2842.900 431.160 2843.160 431.420 ;
      LAYER met2 ;
        RECT 2452.030 510.340 2452.310 514.000 ;
        RECT 2451.960 510.000 2452.310 510.340 ;
        RECT 2451.960 497.070 2452.100 510.000 ;
        RECT 2451.900 496.750 2452.160 497.070 ;
        RECT 2459.720 496.750 2459.980 497.070 ;
        RECT 2459.780 431.450 2459.920 496.750 ;
        RECT 2459.720 431.130 2459.980 431.450 ;
        RECT 2842.900 431.130 2843.160 431.450 ;
        RECT 2842.960 17.410 2843.100 431.130 ;
        RECT 2842.960 17.270 2845.400 17.410 ;
        RECT 2845.260 2.400 2845.400 17.270 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2464.290 496.980 2464.610 497.040 ;
        RECT 2469.350 496.980 2469.670 497.040 ;
        RECT 2464.290 496.840 2469.670 496.980 ;
        RECT 2464.290 496.780 2464.610 496.840 ;
        RECT 2469.350 496.780 2469.670 496.840 ;
        RECT 2469.350 424.220 2469.670 424.280 ;
        RECT 2857.130 424.220 2857.450 424.280 ;
        RECT 2469.350 424.080 2857.450 424.220 ;
        RECT 2469.350 424.020 2469.670 424.080 ;
        RECT 2857.130 424.020 2857.450 424.080 ;
        RECT 2857.130 17.920 2857.450 17.980 ;
        RECT 2863.110 17.920 2863.430 17.980 ;
        RECT 2857.130 17.780 2863.430 17.920 ;
        RECT 2857.130 17.720 2857.450 17.780 ;
        RECT 2863.110 17.720 2863.430 17.780 ;
      LAYER via ;
        RECT 2464.320 496.780 2464.580 497.040 ;
        RECT 2469.380 496.780 2469.640 497.040 ;
        RECT 2469.380 424.020 2469.640 424.280 ;
        RECT 2857.160 424.020 2857.420 424.280 ;
        RECT 2857.160 17.720 2857.420 17.980 ;
        RECT 2863.140 17.720 2863.400 17.980 ;
      LAYER met2 ;
        RECT 2464.450 510.340 2464.730 514.000 ;
        RECT 2464.380 510.000 2464.730 510.340 ;
        RECT 2464.380 497.070 2464.520 510.000 ;
        RECT 2464.320 496.750 2464.580 497.070 ;
        RECT 2469.380 496.750 2469.640 497.070 ;
        RECT 2469.440 424.310 2469.580 496.750 ;
        RECT 2469.380 423.990 2469.640 424.310 ;
        RECT 2857.160 423.990 2857.420 424.310 ;
        RECT 2857.220 18.010 2857.360 423.990 ;
        RECT 2857.160 17.690 2857.420 18.010 ;
        RECT 2863.140 17.690 2863.400 18.010 ;
        RECT 2863.200 2.400 2863.340 17.690 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2477.170 496.980 2477.490 497.040 ;
        RECT 2483.150 496.980 2483.470 497.040 ;
        RECT 2477.170 496.840 2483.470 496.980 ;
        RECT 2477.170 496.780 2477.490 496.840 ;
        RECT 2483.150 496.780 2483.470 496.840 ;
        RECT 2483.150 417.420 2483.470 417.480 ;
        RECT 2873.690 417.420 2874.010 417.480 ;
        RECT 2483.150 417.280 2874.010 417.420 ;
        RECT 2483.150 417.220 2483.470 417.280 ;
        RECT 2873.690 417.220 2874.010 417.280 ;
        RECT 2873.690 16.560 2874.010 16.620 ;
        RECT 2881.050 16.560 2881.370 16.620 ;
        RECT 2873.690 16.420 2881.370 16.560 ;
        RECT 2873.690 16.360 2874.010 16.420 ;
        RECT 2881.050 16.360 2881.370 16.420 ;
      LAYER via ;
        RECT 2477.200 496.780 2477.460 497.040 ;
        RECT 2483.180 496.780 2483.440 497.040 ;
        RECT 2483.180 417.220 2483.440 417.480 ;
        RECT 2873.720 417.220 2873.980 417.480 ;
        RECT 2873.720 16.360 2873.980 16.620 ;
        RECT 2881.080 16.360 2881.340 16.620 ;
      LAYER met2 ;
        RECT 2477.330 510.340 2477.610 514.000 ;
        RECT 2477.260 510.000 2477.610 510.340 ;
        RECT 2477.260 497.070 2477.400 510.000 ;
        RECT 2477.200 496.750 2477.460 497.070 ;
        RECT 2483.180 496.750 2483.440 497.070 ;
        RECT 2483.240 417.510 2483.380 496.750 ;
        RECT 2483.180 417.190 2483.440 417.510 ;
        RECT 2873.720 417.190 2873.980 417.510 ;
        RECT 2873.780 16.650 2873.920 417.190 ;
        RECT 2873.720 16.330 2873.980 16.650 ;
        RECT 2881.080 16.330 2881.340 16.650 ;
        RECT 2881.140 2.400 2881.280 16.330 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.050 500.040 2490.370 500.100 ;
        RECT 2728.790 500.040 2729.110 500.100 ;
        RECT 2490.050 499.900 2729.110 500.040 ;
        RECT 2490.050 499.840 2490.370 499.900 ;
        RECT 2728.790 499.840 2729.110 499.900 ;
        RECT 2728.790 24.040 2729.110 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 2728.790 23.900 2899.310 24.040 ;
        RECT 2728.790 23.840 2729.110 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 2490.080 499.840 2490.340 500.100 ;
        RECT 2728.820 499.840 2729.080 500.100 ;
        RECT 2728.820 23.840 2729.080 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 2490.210 510.340 2490.490 514.000 ;
        RECT 2490.140 510.000 2490.490 510.340 ;
        RECT 2490.140 500.130 2490.280 510.000 ;
        RECT 2490.080 499.810 2490.340 500.130 ;
        RECT 2728.820 499.810 2729.080 500.130 ;
        RECT 2728.880 24.130 2729.020 499.810 ;
        RECT 2728.820 23.810 2729.080 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 38.320 847.250 38.380 ;
        RECT 1014.370 38.320 1014.690 38.380 ;
        RECT 846.930 38.180 1014.690 38.320 ;
        RECT 846.930 38.120 847.250 38.180 ;
        RECT 1014.370 38.120 1014.690 38.180 ;
      LAYER via ;
        RECT 846.960 38.120 847.220 38.380 ;
        RECT 1014.400 38.120 1014.660 38.380 ;
      LAYER met2 ;
        RECT 1017.750 510.410 1018.030 514.000 ;
        RECT 1014.460 510.270 1018.030 510.410 ;
        RECT 1014.460 38.410 1014.600 510.270 ;
        RECT 1017.750 510.000 1018.030 510.270 ;
        RECT 846.960 38.090 847.220 38.410 ;
        RECT 1014.400 38.090 1014.660 38.410 ;
        RECT 847.020 2.400 847.160 38.090 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1017.590 496.980 1017.910 497.040 ;
        RECT 1030.470 496.980 1030.790 497.040 ;
        RECT 1017.590 496.840 1030.790 496.980 ;
        RECT 1017.590 496.780 1017.910 496.840 ;
        RECT 1030.470 496.780 1030.790 496.840 ;
        RECT 864.870 24.040 865.190 24.100 ;
        RECT 1017.590 24.040 1017.910 24.100 ;
        RECT 864.870 23.900 1017.910 24.040 ;
        RECT 864.870 23.840 865.190 23.900 ;
        RECT 1017.590 23.840 1017.910 23.900 ;
      LAYER via ;
        RECT 1017.620 496.780 1017.880 497.040 ;
        RECT 1030.500 496.780 1030.760 497.040 ;
        RECT 864.900 23.840 865.160 24.100 ;
        RECT 1017.620 23.840 1017.880 24.100 ;
      LAYER met2 ;
        RECT 1030.630 510.340 1030.910 514.000 ;
        RECT 1030.560 510.000 1030.910 510.340 ;
        RECT 1030.560 497.070 1030.700 510.000 ;
        RECT 1017.620 496.750 1017.880 497.070 ;
        RECT 1030.500 496.750 1030.760 497.070 ;
        RECT 1017.680 24.130 1017.820 496.750 ;
        RECT 864.900 23.810 865.160 24.130 ;
        RECT 1017.620 23.810 1017.880 24.130 ;
        RECT 864.960 2.400 865.100 23.810 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 44.780 883.130 44.840 ;
        RECT 1041.970 44.780 1042.290 44.840 ;
        RECT 882.810 44.640 1042.290 44.780 ;
        RECT 882.810 44.580 883.130 44.640 ;
        RECT 1041.970 44.580 1042.290 44.640 ;
      LAYER via ;
        RECT 882.840 44.580 883.100 44.840 ;
        RECT 1042.000 44.580 1042.260 44.840 ;
      LAYER met2 ;
        RECT 1043.510 510.410 1043.790 514.000 ;
        RECT 1042.060 510.270 1043.790 510.410 ;
        RECT 1042.060 44.870 1042.200 510.270 ;
        RECT 1043.510 510.000 1043.790 510.270 ;
        RECT 882.840 44.550 883.100 44.870 ;
        RECT 1042.000 44.550 1042.260 44.870 ;
        RECT 882.900 2.400 883.040 44.550 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 51.580 901.070 51.640 ;
        RECT 1055.770 51.580 1056.090 51.640 ;
        RECT 900.750 51.440 1056.090 51.580 ;
        RECT 900.750 51.380 901.070 51.440 ;
        RECT 1055.770 51.380 1056.090 51.440 ;
      LAYER via ;
        RECT 900.780 51.380 901.040 51.640 ;
        RECT 1055.800 51.380 1056.060 51.640 ;
      LAYER met2 ;
        RECT 1056.390 510.410 1056.670 514.000 ;
        RECT 1055.860 510.270 1056.670 510.410 ;
        RECT 1055.860 51.670 1056.000 510.270 ;
        RECT 1056.390 510.000 1056.670 510.270 ;
        RECT 900.780 51.350 901.040 51.670 ;
        RECT 1055.800 51.350 1056.060 51.670 ;
        RECT 900.840 2.400 900.980 51.350 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1063.665 338.045 1063.835 352.495 ;
        RECT 1063.665 269.025 1063.835 331.075 ;
        RECT 1064.125 144.245 1064.295 220.575 ;
        RECT 1064.585 96.305 1064.755 131.155 ;
      LAYER mcon ;
        RECT 1063.665 352.325 1063.835 352.495 ;
        RECT 1063.665 330.905 1063.835 331.075 ;
        RECT 1064.125 220.405 1064.295 220.575 ;
        RECT 1064.585 130.985 1064.755 131.155 ;
      LAYER met1 ;
        RECT 1063.590 410.620 1063.910 410.680 ;
        RECT 1065.430 410.620 1065.750 410.680 ;
        RECT 1063.590 410.480 1065.750 410.620 ;
        RECT 1063.590 410.420 1063.910 410.480 ;
        RECT 1065.430 410.420 1065.750 410.480 ;
        RECT 1063.590 352.480 1063.910 352.540 ;
        RECT 1063.395 352.340 1063.910 352.480 ;
        RECT 1063.590 352.280 1063.910 352.340 ;
        RECT 1063.590 338.200 1063.910 338.260 ;
        RECT 1063.395 338.060 1063.910 338.200 ;
        RECT 1063.590 338.000 1063.910 338.060 ;
        RECT 1063.590 331.060 1063.910 331.120 ;
        RECT 1063.395 330.920 1063.910 331.060 ;
        RECT 1063.590 330.860 1063.910 330.920 ;
        RECT 1063.605 269.180 1063.895 269.225 ;
        RECT 1064.050 269.180 1064.370 269.240 ;
        RECT 1063.605 269.040 1064.370 269.180 ;
        RECT 1063.605 268.995 1063.895 269.040 ;
        RECT 1064.050 268.980 1064.370 269.040 ;
        RECT 1064.050 220.560 1064.370 220.620 ;
        RECT 1063.855 220.420 1064.370 220.560 ;
        RECT 1064.050 220.360 1064.370 220.420 ;
        RECT 1064.050 144.400 1064.370 144.460 ;
        RECT 1063.855 144.260 1064.370 144.400 ;
        RECT 1064.050 144.200 1064.370 144.260 ;
        RECT 1064.050 131.140 1064.370 131.200 ;
        RECT 1064.525 131.140 1064.815 131.185 ;
        RECT 1064.050 131.000 1064.815 131.140 ;
        RECT 1064.050 130.940 1064.370 131.000 ;
        RECT 1064.525 130.955 1064.815 131.000 ;
        RECT 1064.510 96.460 1064.830 96.520 ;
        RECT 1064.315 96.320 1064.830 96.460 ;
        RECT 1064.510 96.260 1064.830 96.320 ;
        RECT 918.690 58.720 919.010 58.780 ;
        RECT 1064.510 58.720 1064.830 58.780 ;
        RECT 918.690 58.580 1064.830 58.720 ;
        RECT 918.690 58.520 919.010 58.580 ;
        RECT 1064.510 58.520 1064.830 58.580 ;
      LAYER via ;
        RECT 1063.620 410.420 1063.880 410.680 ;
        RECT 1065.460 410.420 1065.720 410.680 ;
        RECT 1063.620 352.280 1063.880 352.540 ;
        RECT 1063.620 338.000 1063.880 338.260 ;
        RECT 1063.620 330.860 1063.880 331.120 ;
        RECT 1064.080 268.980 1064.340 269.240 ;
        RECT 1064.080 220.360 1064.340 220.620 ;
        RECT 1064.080 144.200 1064.340 144.460 ;
        RECT 1064.080 130.940 1064.340 131.200 ;
        RECT 1064.540 96.260 1064.800 96.520 ;
        RECT 918.720 58.520 918.980 58.780 ;
        RECT 1064.540 58.520 1064.800 58.780 ;
      LAYER met2 ;
        RECT 1068.810 510.340 1069.090 514.000 ;
        RECT 1068.740 510.000 1069.090 510.340 ;
        RECT 1068.740 483.325 1068.880 510.000 ;
        RECT 1065.450 482.955 1065.730 483.325 ;
        RECT 1068.670 482.955 1068.950 483.325 ;
        RECT 1065.520 410.710 1065.660 482.955 ;
        RECT 1063.620 410.390 1063.880 410.710 ;
        RECT 1065.460 410.390 1065.720 410.710 ;
        RECT 1063.680 352.570 1063.820 410.390 ;
        RECT 1063.620 352.250 1063.880 352.570 ;
        RECT 1063.620 337.970 1063.880 338.290 ;
        RECT 1063.680 331.150 1063.820 337.970 ;
        RECT 1063.620 330.830 1063.880 331.150 ;
        RECT 1064.080 268.950 1064.340 269.270 ;
        RECT 1064.140 220.650 1064.280 268.950 ;
        RECT 1064.080 220.330 1064.340 220.650 ;
        RECT 1064.080 144.170 1064.340 144.490 ;
        RECT 1064.140 131.230 1064.280 144.170 ;
        RECT 1064.080 130.910 1064.340 131.230 ;
        RECT 1064.540 96.230 1064.800 96.550 ;
        RECT 1064.600 58.810 1064.740 96.230 ;
        RECT 918.720 58.490 918.980 58.810 ;
        RECT 1064.540 58.490 1064.800 58.810 ;
        RECT 918.780 2.400 918.920 58.490 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 1065.450 483.000 1065.730 483.280 ;
        RECT 1068.670 483.000 1068.950 483.280 ;
      LAYER met3 ;
        RECT 1065.425 483.290 1065.755 483.305 ;
        RECT 1068.645 483.290 1068.975 483.305 ;
        RECT 1065.425 482.990 1068.975 483.290 ;
        RECT 1065.425 482.975 1065.755 482.990 ;
        RECT 1068.645 482.975 1068.975 482.990 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1077.005 379.525 1077.175 427.635 ;
      LAYER mcon ;
        RECT 1077.005 427.465 1077.175 427.635 ;
      LAYER met1 ;
        RECT 1077.850 476.240 1078.170 476.300 ;
        RECT 1081.530 476.240 1081.850 476.300 ;
        RECT 1077.850 476.100 1081.850 476.240 ;
        RECT 1077.850 476.040 1078.170 476.100 ;
        RECT 1081.530 476.040 1081.850 476.100 ;
        RECT 1076.945 427.620 1077.235 427.665 ;
        RECT 1077.390 427.620 1077.710 427.680 ;
        RECT 1076.945 427.480 1077.710 427.620 ;
        RECT 1076.945 427.435 1077.235 427.480 ;
        RECT 1077.390 427.420 1077.710 427.480 ;
        RECT 1076.930 379.680 1077.250 379.740 ;
        RECT 1076.735 379.540 1077.250 379.680 ;
        RECT 1076.930 379.480 1077.250 379.540 ;
        RECT 1076.930 314.060 1077.250 314.120 ;
        RECT 1077.850 314.060 1078.170 314.120 ;
        RECT 1076.930 313.920 1078.170 314.060 ;
        RECT 1076.930 313.860 1077.250 313.920 ;
        RECT 1077.850 313.860 1078.170 313.920 ;
        RECT 1077.390 241.640 1077.710 241.700 ;
        RECT 1077.850 241.640 1078.170 241.700 ;
        RECT 1077.390 241.500 1078.170 241.640 ;
        RECT 1077.390 241.440 1077.710 241.500 ;
        RECT 1077.850 241.440 1078.170 241.500 ;
        RECT 938.010 65.520 938.330 65.580 ;
        RECT 1077.390 65.520 1077.710 65.580 ;
        RECT 938.010 65.380 1077.710 65.520 ;
        RECT 938.010 65.320 938.330 65.380 ;
        RECT 1077.390 65.320 1077.710 65.380 ;
      LAYER via ;
        RECT 1077.880 476.040 1078.140 476.300 ;
        RECT 1081.560 476.040 1081.820 476.300 ;
        RECT 1077.420 427.420 1077.680 427.680 ;
        RECT 1076.960 379.480 1077.220 379.740 ;
        RECT 1076.960 313.860 1077.220 314.120 ;
        RECT 1077.880 313.860 1078.140 314.120 ;
        RECT 1077.420 241.440 1077.680 241.700 ;
        RECT 1077.880 241.440 1078.140 241.700 ;
        RECT 938.040 65.320 938.300 65.580 ;
        RECT 1077.420 65.320 1077.680 65.580 ;
      LAYER met2 ;
        RECT 1081.690 510.340 1081.970 514.000 ;
        RECT 1081.620 510.000 1081.970 510.340 ;
        RECT 1081.620 476.330 1081.760 510.000 ;
        RECT 1077.880 476.010 1078.140 476.330 ;
        RECT 1081.560 476.010 1081.820 476.330 ;
        RECT 1077.940 434.930 1078.080 476.010 ;
        RECT 1077.480 434.790 1078.080 434.930 ;
        RECT 1077.480 427.710 1077.620 434.790 ;
        RECT 1077.420 427.390 1077.680 427.710 ;
        RECT 1076.960 379.450 1077.220 379.770 ;
        RECT 1077.020 314.150 1077.160 379.450 ;
        RECT 1076.960 313.830 1077.220 314.150 ;
        RECT 1077.880 313.830 1078.140 314.150 ;
        RECT 1077.940 241.730 1078.080 313.830 ;
        RECT 1077.420 241.410 1077.680 241.730 ;
        RECT 1077.880 241.410 1078.140 241.730 ;
        RECT 1077.480 207.810 1077.620 241.410 ;
        RECT 1077.480 207.670 1078.080 207.810 ;
        RECT 1077.940 206.960 1078.080 207.670 ;
        RECT 1077.480 206.820 1078.080 206.960 ;
        RECT 1077.480 65.610 1077.620 206.820 ;
        RECT 938.040 65.290 938.300 65.610 ;
        RECT 1077.420 65.290 1077.680 65.610 ;
        RECT 938.100 17.410 938.240 65.290 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1090.805 379.525 1090.975 427.635 ;
      LAYER mcon ;
        RECT 1090.805 427.465 1090.975 427.635 ;
      LAYER met1 ;
        RECT 1091.650 484.400 1091.970 484.460 ;
        RECT 1094.410 484.400 1094.730 484.460 ;
        RECT 1091.650 484.260 1094.730 484.400 ;
        RECT 1091.650 484.200 1091.970 484.260 ;
        RECT 1094.410 484.200 1094.730 484.260 ;
        RECT 1091.650 435.780 1091.970 435.840 ;
        RECT 1091.280 435.640 1091.970 435.780 ;
        RECT 1091.280 435.160 1091.420 435.640 ;
        RECT 1091.650 435.580 1091.970 435.640 ;
        RECT 1091.190 434.900 1091.510 435.160 ;
        RECT 1090.745 427.620 1091.035 427.665 ;
        RECT 1091.190 427.620 1091.510 427.680 ;
        RECT 1090.745 427.480 1091.510 427.620 ;
        RECT 1090.745 427.435 1091.035 427.480 ;
        RECT 1091.190 427.420 1091.510 427.480 ;
        RECT 1090.730 379.680 1091.050 379.740 ;
        RECT 1090.535 379.540 1091.050 379.680 ;
        RECT 1090.730 379.480 1091.050 379.540 ;
        RECT 1090.730 314.060 1091.050 314.120 ;
        RECT 1091.650 314.060 1091.970 314.120 ;
        RECT 1090.730 313.920 1091.970 314.060 ;
        RECT 1090.730 313.860 1091.050 313.920 ;
        RECT 1091.650 313.860 1091.970 313.920 ;
        RECT 1091.190 241.640 1091.510 241.700 ;
        RECT 1091.650 241.640 1091.970 241.700 ;
        RECT 1091.190 241.500 1091.970 241.640 ;
        RECT 1091.190 241.440 1091.510 241.500 ;
        RECT 1091.650 241.440 1091.970 241.500 ;
        RECT 958.710 72.320 959.030 72.380 ;
        RECT 1091.190 72.320 1091.510 72.380 ;
        RECT 958.710 72.180 1091.510 72.320 ;
        RECT 958.710 72.120 959.030 72.180 ;
        RECT 1091.190 72.120 1091.510 72.180 ;
        RECT 954.110 16.900 954.430 16.960 ;
        RECT 958.710 16.900 959.030 16.960 ;
        RECT 954.110 16.760 959.030 16.900 ;
        RECT 954.110 16.700 954.430 16.760 ;
        RECT 958.710 16.700 959.030 16.760 ;
      LAYER via ;
        RECT 1091.680 484.200 1091.940 484.460 ;
        RECT 1094.440 484.200 1094.700 484.460 ;
        RECT 1091.680 435.580 1091.940 435.840 ;
        RECT 1091.220 434.900 1091.480 435.160 ;
        RECT 1091.220 427.420 1091.480 427.680 ;
        RECT 1090.760 379.480 1091.020 379.740 ;
        RECT 1090.760 313.860 1091.020 314.120 ;
        RECT 1091.680 313.860 1091.940 314.120 ;
        RECT 1091.220 241.440 1091.480 241.700 ;
        RECT 1091.680 241.440 1091.940 241.700 ;
        RECT 958.740 72.120 959.000 72.380 ;
        RECT 1091.220 72.120 1091.480 72.380 ;
        RECT 954.140 16.700 954.400 16.960 ;
        RECT 958.740 16.700 959.000 16.960 ;
      LAYER met2 ;
        RECT 1094.570 510.340 1094.850 514.000 ;
        RECT 1094.500 510.000 1094.850 510.340 ;
        RECT 1094.500 484.490 1094.640 510.000 ;
        RECT 1091.680 484.170 1091.940 484.490 ;
        RECT 1094.440 484.170 1094.700 484.490 ;
        RECT 1091.740 435.870 1091.880 484.170 ;
        RECT 1091.680 435.550 1091.940 435.870 ;
        RECT 1091.220 434.870 1091.480 435.190 ;
        RECT 1091.280 427.710 1091.420 434.870 ;
        RECT 1091.220 427.390 1091.480 427.710 ;
        RECT 1090.760 379.450 1091.020 379.770 ;
        RECT 1090.820 314.150 1090.960 379.450 ;
        RECT 1090.760 313.830 1091.020 314.150 ;
        RECT 1091.680 313.830 1091.940 314.150 ;
        RECT 1091.740 241.730 1091.880 313.830 ;
        RECT 1091.220 241.410 1091.480 241.730 ;
        RECT 1091.680 241.410 1091.940 241.730 ;
        RECT 1091.280 72.410 1091.420 241.410 ;
        RECT 958.740 72.090 959.000 72.410 ;
        RECT 1091.220 72.090 1091.480 72.410 ;
        RECT 958.800 16.990 958.940 72.090 ;
        RECT 954.140 16.670 954.400 16.990 ;
        RECT 958.740 16.670 959.000 16.990 ;
        RECT 954.200 2.400 954.340 16.670 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 31.180 972.370 31.240 ;
        RECT 1104.070 31.180 1104.390 31.240 ;
        RECT 972.050 31.040 1104.390 31.180 ;
        RECT 972.050 30.980 972.370 31.040 ;
        RECT 1104.070 30.980 1104.390 31.040 ;
      LAYER via ;
        RECT 972.080 30.980 972.340 31.240 ;
        RECT 1104.100 30.980 1104.360 31.240 ;
      LAYER met2 ;
        RECT 1107.450 510.410 1107.730 514.000 ;
        RECT 1104.160 510.270 1107.730 510.410 ;
        RECT 1104.160 31.270 1104.300 510.270 ;
        RECT 1107.450 510.000 1107.730 510.270 ;
        RECT 972.080 30.950 972.340 31.270 ;
        RECT 1104.100 30.950 1104.360 31.270 ;
        RECT 972.140 2.400 972.280 30.950 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 45.120 651.290 45.180 ;
        RECT 876.370 45.120 876.690 45.180 ;
        RECT 650.970 44.980 876.690 45.120 ;
        RECT 650.970 44.920 651.290 44.980 ;
        RECT 876.370 44.920 876.690 44.980 ;
      LAYER via ;
        RECT 651.000 44.920 651.260 45.180 ;
        RECT 876.400 44.920 876.660 45.180 ;
      LAYER met2 ;
        RECT 876.990 510.410 877.270 514.000 ;
        RECT 876.460 510.270 877.270 510.410 ;
        RECT 876.460 45.210 876.600 510.270 ;
        RECT 876.990 510.000 877.270 510.270 ;
        RECT 651.000 44.890 651.260 45.210 ;
        RECT 876.400 44.890 876.660 45.210 ;
        RECT 651.060 2.400 651.200 44.890 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1038.290 500.040 1038.610 500.100 ;
        RECT 1120.170 500.040 1120.490 500.100 ;
        RECT 1038.290 499.900 1120.490 500.040 ;
        RECT 1038.290 499.840 1038.610 499.900 ;
        RECT 1120.170 499.840 1120.490 499.900 ;
        RECT 993.210 79.460 993.530 79.520 ;
        RECT 1038.290 79.460 1038.610 79.520 ;
        RECT 993.210 79.320 1038.610 79.460 ;
        RECT 993.210 79.260 993.530 79.320 ;
        RECT 1038.290 79.260 1038.610 79.320 ;
        RECT 989.990 16.900 990.310 16.960 ;
        RECT 993.210 16.900 993.530 16.960 ;
        RECT 989.990 16.760 993.530 16.900 ;
        RECT 989.990 16.700 990.310 16.760 ;
        RECT 993.210 16.700 993.530 16.760 ;
      LAYER via ;
        RECT 1038.320 499.840 1038.580 500.100 ;
        RECT 1120.200 499.840 1120.460 500.100 ;
        RECT 993.240 79.260 993.500 79.520 ;
        RECT 1038.320 79.260 1038.580 79.520 ;
        RECT 990.020 16.700 990.280 16.960 ;
        RECT 993.240 16.700 993.500 16.960 ;
      LAYER met2 ;
        RECT 1120.330 510.340 1120.610 514.000 ;
        RECT 1120.260 510.000 1120.610 510.340 ;
        RECT 1120.260 500.130 1120.400 510.000 ;
        RECT 1038.320 499.810 1038.580 500.130 ;
        RECT 1120.200 499.810 1120.460 500.130 ;
        RECT 1038.380 79.550 1038.520 499.810 ;
        RECT 993.240 79.230 993.500 79.550 ;
        RECT 1038.320 79.230 1038.580 79.550 ;
        RECT 993.300 16.990 993.440 79.230 ;
        RECT 990.020 16.670 990.280 16.990 ;
        RECT 993.240 16.670 993.500 16.990 ;
        RECT 990.080 2.400 990.220 16.670 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 24.380 1007.790 24.440 ;
        RECT 1131.670 24.380 1131.990 24.440 ;
        RECT 1007.470 24.240 1131.990 24.380 ;
        RECT 1007.470 24.180 1007.790 24.240 ;
        RECT 1131.670 24.180 1131.990 24.240 ;
      LAYER via ;
        RECT 1007.500 24.180 1007.760 24.440 ;
        RECT 1131.700 24.180 1131.960 24.440 ;
      LAYER met2 ;
        RECT 1133.210 510.410 1133.490 514.000 ;
        RECT 1131.760 510.270 1133.490 510.410 ;
        RECT 1131.760 24.470 1131.900 510.270 ;
        RECT 1133.210 510.000 1133.490 510.270 ;
        RECT 1007.500 24.150 1007.760 24.470 ;
        RECT 1131.700 24.150 1131.960 24.470 ;
        RECT 1007.560 2.400 1007.700 24.150 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.410 37.980 1025.730 38.040 ;
        RECT 1145.470 37.980 1145.790 38.040 ;
        RECT 1025.410 37.840 1145.790 37.980 ;
        RECT 1025.410 37.780 1025.730 37.840 ;
        RECT 1145.470 37.780 1145.790 37.840 ;
      LAYER via ;
        RECT 1025.440 37.780 1025.700 38.040 ;
        RECT 1145.500 37.780 1145.760 38.040 ;
      LAYER met2 ;
        RECT 1145.630 510.340 1145.910 514.000 ;
        RECT 1145.560 510.000 1145.910 510.340 ;
        RECT 1145.560 38.070 1145.700 510.000 ;
        RECT 1025.440 37.750 1025.700 38.070 ;
        RECT 1145.500 37.750 1145.760 38.070 ;
        RECT 1025.500 2.400 1025.640 37.750 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1154.285 427.805 1154.455 435.115 ;
        RECT 1153.365 96.645 1153.535 110.755 ;
      LAYER mcon ;
        RECT 1154.285 434.945 1154.455 435.115 ;
        RECT 1153.365 110.585 1153.535 110.755 ;
      LAYER met1 ;
        RECT 1154.210 476.240 1154.530 476.300 ;
        RECT 1158.350 476.240 1158.670 476.300 ;
        RECT 1154.210 476.100 1158.670 476.240 ;
        RECT 1154.210 476.040 1154.530 476.100 ;
        RECT 1158.350 476.040 1158.670 476.100 ;
        RECT 1154.210 435.100 1154.530 435.160 ;
        RECT 1154.015 434.960 1154.530 435.100 ;
        RECT 1154.210 434.900 1154.530 434.960 ;
        RECT 1154.210 427.960 1154.530 428.020 ;
        RECT 1154.015 427.820 1154.530 427.960 ;
        RECT 1154.210 427.760 1154.530 427.820 ;
        RECT 1154.210 383.220 1154.530 383.480 ;
        RECT 1154.300 382.800 1154.440 383.220 ;
        RECT 1154.210 382.540 1154.530 382.800 ;
        RECT 1153.290 331.060 1153.610 331.120 ;
        RECT 1153.750 331.060 1154.070 331.120 ;
        RECT 1153.290 330.920 1154.070 331.060 ;
        RECT 1153.290 330.860 1153.610 330.920 ;
        RECT 1153.750 330.860 1154.070 330.920 ;
        RECT 1153.750 193.360 1154.070 193.420 ;
        RECT 1154.210 193.360 1154.530 193.420 ;
        RECT 1153.750 193.220 1154.530 193.360 ;
        RECT 1153.750 193.160 1154.070 193.220 ;
        RECT 1154.210 193.160 1154.530 193.220 ;
        RECT 1153.305 110.740 1153.595 110.785 ;
        RECT 1153.750 110.740 1154.070 110.800 ;
        RECT 1153.305 110.600 1154.070 110.740 ;
        RECT 1153.305 110.555 1153.595 110.600 ;
        RECT 1153.750 110.540 1154.070 110.600 ;
        RECT 1153.290 96.800 1153.610 96.860 ;
        RECT 1153.095 96.660 1153.610 96.800 ;
        RECT 1153.290 96.600 1153.610 96.660 ;
        RECT 1043.350 44.780 1043.670 44.840 ;
        RECT 1153.750 44.780 1154.070 44.840 ;
        RECT 1043.350 44.640 1154.070 44.780 ;
        RECT 1043.350 44.580 1043.670 44.640 ;
        RECT 1153.750 44.580 1154.070 44.640 ;
      LAYER via ;
        RECT 1154.240 476.040 1154.500 476.300 ;
        RECT 1158.380 476.040 1158.640 476.300 ;
        RECT 1154.240 434.900 1154.500 435.160 ;
        RECT 1154.240 427.760 1154.500 428.020 ;
        RECT 1154.240 383.220 1154.500 383.480 ;
        RECT 1154.240 382.540 1154.500 382.800 ;
        RECT 1153.320 330.860 1153.580 331.120 ;
        RECT 1153.780 330.860 1154.040 331.120 ;
        RECT 1153.780 193.160 1154.040 193.420 ;
        RECT 1154.240 193.160 1154.500 193.420 ;
        RECT 1153.780 110.540 1154.040 110.800 ;
        RECT 1153.320 96.600 1153.580 96.860 ;
        RECT 1043.380 44.580 1043.640 44.840 ;
        RECT 1153.780 44.580 1154.040 44.840 ;
      LAYER met2 ;
        RECT 1158.510 510.340 1158.790 514.000 ;
        RECT 1158.440 510.000 1158.790 510.340 ;
        RECT 1158.440 476.330 1158.580 510.000 ;
        RECT 1154.240 476.010 1154.500 476.330 ;
        RECT 1158.380 476.010 1158.640 476.330 ;
        RECT 1154.300 435.190 1154.440 476.010 ;
        RECT 1154.240 434.870 1154.500 435.190 ;
        RECT 1154.240 427.730 1154.500 428.050 ;
        RECT 1154.300 383.510 1154.440 427.730 ;
        RECT 1154.240 383.190 1154.500 383.510 ;
        RECT 1154.240 382.510 1154.500 382.830 ;
        RECT 1154.300 338.485 1154.440 382.510 ;
        RECT 1153.310 338.115 1153.590 338.485 ;
        RECT 1154.230 338.115 1154.510 338.485 ;
        RECT 1153.380 331.150 1153.520 338.115 ;
        RECT 1153.320 330.830 1153.580 331.150 ;
        RECT 1153.780 330.830 1154.040 331.150 ;
        RECT 1153.840 265.610 1153.980 330.830 ;
        RECT 1153.840 265.470 1154.440 265.610 ;
        RECT 1154.300 193.450 1154.440 265.470 ;
        RECT 1153.780 193.130 1154.040 193.450 ;
        RECT 1154.240 193.130 1154.500 193.450 ;
        RECT 1153.840 110.830 1153.980 193.130 ;
        RECT 1153.780 110.510 1154.040 110.830 ;
        RECT 1153.320 96.570 1153.580 96.890 ;
        RECT 1153.380 62.290 1153.520 96.570 ;
        RECT 1153.380 62.150 1153.980 62.290 ;
        RECT 1153.840 44.870 1153.980 62.150 ;
        RECT 1043.380 44.550 1043.640 44.870 ;
        RECT 1153.780 44.550 1154.040 44.870 ;
        RECT 1043.440 2.400 1043.580 44.550 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1153.310 338.160 1153.590 338.440 ;
        RECT 1154.230 338.160 1154.510 338.440 ;
      LAYER met3 ;
        RECT 1153.285 338.450 1153.615 338.465 ;
        RECT 1154.205 338.450 1154.535 338.465 ;
        RECT 1153.285 338.150 1154.535 338.450 ;
        RECT 1153.285 338.135 1153.615 338.150 ;
        RECT 1154.205 338.135 1154.535 338.150 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 472.840 1166.950 472.900 ;
        RECT 1169.390 472.840 1169.710 472.900 ;
        RECT 1166.630 472.700 1169.710 472.840 ;
        RECT 1166.630 472.640 1166.950 472.700 ;
        RECT 1169.390 472.640 1169.710 472.700 ;
        RECT 1061.290 51.580 1061.610 51.640 ;
        RECT 1166.630 51.580 1166.950 51.640 ;
        RECT 1061.290 51.440 1166.950 51.580 ;
        RECT 1061.290 51.380 1061.610 51.440 ;
        RECT 1166.630 51.380 1166.950 51.440 ;
      LAYER via ;
        RECT 1166.660 472.640 1166.920 472.900 ;
        RECT 1169.420 472.640 1169.680 472.900 ;
        RECT 1061.320 51.380 1061.580 51.640 ;
        RECT 1166.660 51.380 1166.920 51.640 ;
      LAYER met2 ;
        RECT 1171.390 510.410 1171.670 514.000 ;
        RECT 1169.480 510.270 1171.670 510.410 ;
        RECT 1169.480 472.930 1169.620 510.270 ;
        RECT 1171.390 510.000 1171.670 510.270 ;
        RECT 1166.660 472.610 1166.920 472.930 ;
        RECT 1169.420 472.610 1169.680 472.930 ;
        RECT 1166.720 51.670 1166.860 472.610 ;
        RECT 1061.320 51.350 1061.580 51.670 ;
        RECT 1166.660 51.350 1166.920 51.670 ;
        RECT 1061.380 2.400 1061.520 51.350 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.430 472.840 1180.750 472.900 ;
        RECT 1182.270 472.840 1182.590 472.900 ;
        RECT 1180.430 472.700 1182.590 472.840 ;
        RECT 1180.430 472.640 1180.750 472.700 ;
        RECT 1182.270 472.640 1182.590 472.700 ;
        RECT 1079.230 58.720 1079.550 58.780 ;
        RECT 1180.430 58.720 1180.750 58.780 ;
        RECT 1079.230 58.580 1180.750 58.720 ;
        RECT 1079.230 58.520 1079.550 58.580 ;
        RECT 1180.430 58.520 1180.750 58.580 ;
      LAYER via ;
        RECT 1180.460 472.640 1180.720 472.900 ;
        RECT 1182.300 472.640 1182.560 472.900 ;
        RECT 1079.260 58.520 1079.520 58.780 ;
        RECT 1180.460 58.520 1180.720 58.780 ;
      LAYER met2 ;
        RECT 1184.270 510.410 1184.550 514.000 ;
        RECT 1182.360 510.270 1184.550 510.410 ;
        RECT 1182.360 472.930 1182.500 510.270 ;
        RECT 1184.270 510.000 1184.550 510.270 ;
        RECT 1180.460 472.610 1180.720 472.930 ;
        RECT 1182.300 472.610 1182.560 472.930 ;
        RECT 1180.520 58.810 1180.660 472.610 ;
        RECT 1079.260 58.490 1079.520 58.810 ;
        RECT 1180.460 58.490 1180.720 58.810 ;
        RECT 1079.320 2.400 1079.460 58.490 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 65.520 1097.030 65.580 ;
        RECT 1193.770 65.520 1194.090 65.580 ;
        RECT 1096.710 65.380 1194.090 65.520 ;
        RECT 1096.710 65.320 1097.030 65.380 ;
        RECT 1193.770 65.320 1194.090 65.380 ;
      LAYER via ;
        RECT 1096.740 65.320 1097.000 65.580 ;
        RECT 1193.800 65.320 1194.060 65.580 ;
      LAYER met2 ;
        RECT 1197.150 510.410 1197.430 514.000 ;
        RECT 1193.860 510.270 1197.430 510.410 ;
        RECT 1193.860 65.610 1194.000 510.270 ;
        RECT 1197.150 510.000 1197.430 510.270 ;
        RECT 1096.740 65.290 1097.000 65.610 ;
        RECT 1193.800 65.290 1194.060 65.610 ;
        RECT 1096.800 2.400 1096.940 65.290 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 496.980 1197.310 497.040 ;
        RECT 1209.870 496.980 1210.190 497.040 ;
        RECT 1196.990 496.840 1210.190 496.980 ;
        RECT 1196.990 496.780 1197.310 496.840 ;
        RECT 1209.870 496.780 1210.190 496.840 ;
        RECT 1114.650 30.840 1114.970 30.900 ;
        RECT 1196.990 30.840 1197.310 30.900 ;
        RECT 1114.650 30.700 1197.310 30.840 ;
        RECT 1114.650 30.640 1114.970 30.700 ;
        RECT 1196.990 30.640 1197.310 30.700 ;
      LAYER via ;
        RECT 1197.020 496.780 1197.280 497.040 ;
        RECT 1209.900 496.780 1210.160 497.040 ;
        RECT 1114.680 30.640 1114.940 30.900 ;
        RECT 1197.020 30.640 1197.280 30.900 ;
      LAYER met2 ;
        RECT 1210.030 510.340 1210.310 514.000 ;
        RECT 1209.960 510.000 1210.310 510.340 ;
        RECT 1209.960 497.070 1210.100 510.000 ;
        RECT 1197.020 496.750 1197.280 497.070 ;
        RECT 1209.900 496.750 1210.160 497.070 ;
        RECT 1197.080 30.930 1197.220 496.750 ;
        RECT 1114.680 30.610 1114.940 30.930 ;
        RECT 1197.020 30.610 1197.280 30.930 ;
        RECT 1114.740 2.400 1114.880 30.610 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.590 24.040 1132.910 24.100 ;
        RECT 1221.830 24.040 1222.150 24.100 ;
        RECT 1132.590 23.900 1222.150 24.040 ;
        RECT 1132.590 23.840 1132.910 23.900 ;
        RECT 1221.830 23.840 1222.150 23.900 ;
      LAYER via ;
        RECT 1132.620 23.840 1132.880 24.100 ;
        RECT 1221.860 23.840 1222.120 24.100 ;
      LAYER met2 ;
        RECT 1222.450 510.410 1222.730 514.000 ;
        RECT 1221.920 510.270 1222.730 510.410 ;
        RECT 1221.920 24.130 1222.060 510.270 ;
        RECT 1222.450 510.000 1222.730 510.270 ;
        RECT 1132.620 23.810 1132.880 24.130 ;
        RECT 1221.860 23.810 1222.120 24.130 ;
        RECT 1132.680 2.400 1132.820 23.810 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 37.980 1150.850 38.040 ;
        RECT 1235.630 37.980 1235.950 38.040 ;
        RECT 1150.530 37.840 1235.950 37.980 ;
        RECT 1150.530 37.780 1150.850 37.840 ;
        RECT 1235.630 37.780 1235.950 37.840 ;
      LAYER via ;
        RECT 1150.560 37.780 1150.820 38.040 ;
        RECT 1235.660 37.780 1235.920 38.040 ;
      LAYER met2 ;
        RECT 1235.330 510.340 1235.610 514.000 ;
        RECT 1235.260 510.000 1235.610 510.340 ;
        RECT 1235.260 473.690 1235.400 510.000 ;
        RECT 1235.260 473.550 1235.860 473.690 ;
        RECT 1235.720 38.070 1235.860 473.550 ;
        RECT 1150.560 37.750 1150.820 38.070 ;
        RECT 1235.660 37.750 1235.920 38.070 ;
        RECT 1150.620 2.400 1150.760 37.750 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 883.805 138.125 883.975 173.315 ;
        RECT 883.805 51.425 883.975 62.475 ;
      LAYER mcon ;
        RECT 883.805 173.145 883.975 173.315 ;
        RECT 883.805 62.305 883.975 62.475 ;
      LAYER met1 ;
        RECT 883.270 400.420 883.590 400.480 ;
        RECT 885.570 400.420 885.890 400.480 ;
        RECT 883.270 400.280 885.890 400.420 ;
        RECT 883.270 400.220 883.590 400.280 ;
        RECT 885.570 400.220 885.890 400.280 ;
        RECT 884.190 349.220 884.510 349.480 ;
        RECT 884.280 348.800 884.420 349.220 ;
        RECT 884.190 348.540 884.510 348.800 ;
        RECT 884.190 304.200 884.510 304.260 ;
        RECT 883.820 304.060 884.510 304.200 ;
        RECT 883.820 303.920 883.960 304.060 ;
        RECT 884.190 304.000 884.510 304.060 ;
        RECT 883.730 303.660 884.050 303.920 ;
        RECT 883.270 241.640 883.590 241.700 ;
        RECT 884.650 241.640 884.970 241.700 ;
        RECT 883.270 241.500 884.970 241.640 ;
        RECT 883.270 241.440 883.590 241.500 ;
        RECT 884.650 241.440 884.970 241.500 ;
        RECT 884.650 193.700 884.970 193.760 ;
        RECT 884.280 193.560 884.970 193.700 ;
        RECT 884.280 193.420 884.420 193.560 ;
        RECT 884.650 193.500 884.970 193.560 ;
        RECT 884.190 193.160 884.510 193.420 ;
        RECT 883.730 173.300 884.050 173.360 ;
        RECT 883.535 173.160 884.050 173.300 ;
        RECT 883.730 173.100 884.050 173.160 ;
        RECT 883.745 138.280 884.035 138.325 ;
        RECT 884.650 138.280 884.970 138.340 ;
        RECT 883.745 138.140 884.970 138.280 ;
        RECT 883.745 138.095 884.035 138.140 ;
        RECT 884.650 138.080 884.970 138.140 ;
        RECT 884.650 110.740 884.970 110.800 ;
        RECT 883.820 110.600 884.970 110.740 ;
        RECT 883.820 110.460 883.960 110.600 ;
        RECT 884.650 110.540 884.970 110.600 ;
        RECT 883.730 110.200 884.050 110.460 ;
        RECT 883.730 62.460 884.050 62.520 ;
        RECT 883.535 62.320 884.050 62.460 ;
        RECT 883.730 62.260 884.050 62.320 ;
        RECT 668.910 51.580 669.230 51.640 ;
        RECT 883.745 51.580 884.035 51.625 ;
        RECT 668.910 51.440 884.035 51.580 ;
        RECT 668.910 51.380 669.230 51.440 ;
        RECT 883.745 51.395 884.035 51.440 ;
      LAYER via ;
        RECT 883.300 400.220 883.560 400.480 ;
        RECT 885.600 400.220 885.860 400.480 ;
        RECT 884.220 349.220 884.480 349.480 ;
        RECT 884.220 348.540 884.480 348.800 ;
        RECT 884.220 304.000 884.480 304.260 ;
        RECT 883.760 303.660 884.020 303.920 ;
        RECT 883.300 241.440 883.560 241.700 ;
        RECT 884.680 241.440 884.940 241.700 ;
        RECT 884.680 193.500 884.940 193.760 ;
        RECT 884.220 193.160 884.480 193.420 ;
        RECT 883.760 173.100 884.020 173.360 ;
        RECT 884.680 138.080 884.940 138.340 ;
        RECT 884.680 110.540 884.940 110.800 ;
        RECT 883.760 110.200 884.020 110.460 ;
        RECT 883.760 62.260 884.020 62.520 ;
        RECT 668.940 51.380 669.200 51.640 ;
      LAYER met2 ;
        RECT 889.870 510.410 890.150 514.000 ;
        RECT 886.580 510.270 890.150 510.410 ;
        RECT 886.580 449.210 886.720 510.270 ;
        RECT 889.870 510.000 890.150 510.270 ;
        RECT 886.120 449.070 886.720 449.210 ;
        RECT 886.120 400.930 886.260 449.070 ;
        RECT 885.660 400.790 886.260 400.930 ;
        RECT 883.360 400.510 883.500 400.665 ;
        RECT 885.660 400.510 885.800 400.790 ;
        RECT 883.300 400.250 883.560 400.510 ;
        RECT 883.300 400.190 884.420 400.250 ;
        RECT 885.600 400.190 885.860 400.510 ;
        RECT 883.360 400.110 884.420 400.190 ;
        RECT 884.280 349.510 884.420 400.110 ;
        RECT 884.220 349.190 884.480 349.510 ;
        RECT 884.220 348.510 884.480 348.830 ;
        RECT 884.280 304.290 884.420 348.510 ;
        RECT 884.220 303.970 884.480 304.290 ;
        RECT 883.760 303.630 884.020 303.950 ;
        RECT 883.820 265.610 883.960 303.630 ;
        RECT 883.360 265.470 883.960 265.610 ;
        RECT 883.360 241.730 883.500 265.470 ;
        RECT 883.300 241.410 883.560 241.730 ;
        RECT 884.680 241.410 884.940 241.730 ;
        RECT 884.740 193.790 884.880 241.410 ;
        RECT 884.680 193.470 884.940 193.790 ;
        RECT 884.220 193.130 884.480 193.450 ;
        RECT 884.280 192.850 884.420 193.130 ;
        RECT 883.820 192.710 884.420 192.850 ;
        RECT 883.820 173.390 883.960 192.710 ;
        RECT 883.760 173.070 884.020 173.390 ;
        RECT 884.680 138.050 884.940 138.370 ;
        RECT 884.740 110.830 884.880 138.050 ;
        RECT 884.680 110.510 884.940 110.830 ;
        RECT 883.760 110.170 884.020 110.490 ;
        RECT 883.820 62.550 883.960 110.170 ;
        RECT 883.760 62.230 884.020 62.550 ;
        RECT 668.940 51.350 669.200 51.670 ;
        RECT 669.000 2.400 669.140 51.350 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1244.445 386.325 1244.615 400.775 ;
        RECT 1243.065 338.045 1243.235 352.155 ;
        RECT 1244.905 186.405 1245.075 234.515 ;
        RECT 1243.065 51.425 1243.235 96.475 ;
      LAYER mcon ;
        RECT 1244.445 400.605 1244.615 400.775 ;
        RECT 1243.065 351.985 1243.235 352.155 ;
        RECT 1244.905 234.345 1245.075 234.515 ;
        RECT 1243.065 96.305 1243.235 96.475 ;
      LAYER met1 ;
        RECT 1244.370 435.100 1244.690 435.160 ;
        RECT 1244.830 435.100 1245.150 435.160 ;
        RECT 1244.370 434.960 1245.150 435.100 ;
        RECT 1244.370 434.900 1244.690 434.960 ;
        RECT 1244.830 434.900 1245.150 434.960 ;
        RECT 1244.370 400.760 1244.690 400.820 ;
        RECT 1244.175 400.620 1244.690 400.760 ;
        RECT 1244.370 400.560 1244.690 400.620 ;
        RECT 1242.990 386.480 1243.310 386.540 ;
        RECT 1244.385 386.480 1244.675 386.525 ;
        RECT 1242.990 386.340 1244.675 386.480 ;
        RECT 1242.990 386.280 1243.310 386.340 ;
        RECT 1244.385 386.295 1244.675 386.340 ;
        RECT 1242.990 352.140 1243.310 352.200 ;
        RECT 1242.795 352.000 1243.310 352.140 ;
        RECT 1242.990 351.940 1243.310 352.000 ;
        RECT 1242.990 338.200 1243.310 338.260 ;
        RECT 1242.795 338.060 1243.310 338.200 ;
        RECT 1242.990 338.000 1243.310 338.060 ;
        RECT 1243.450 303.660 1243.770 303.920 ;
        RECT 1243.540 303.240 1243.680 303.660 ;
        RECT 1243.450 302.980 1243.770 303.240 ;
        RECT 1244.830 234.500 1245.150 234.560 ;
        RECT 1244.635 234.360 1245.150 234.500 ;
        RECT 1244.830 234.300 1245.150 234.360 ;
        RECT 1244.830 186.560 1245.150 186.620 ;
        RECT 1244.635 186.420 1245.150 186.560 ;
        RECT 1244.830 186.360 1245.150 186.420 ;
        RECT 1243.450 145.080 1243.770 145.140 ;
        RECT 1244.830 145.080 1245.150 145.140 ;
        RECT 1243.450 144.940 1245.150 145.080 ;
        RECT 1243.450 144.880 1243.770 144.940 ;
        RECT 1244.830 144.880 1245.150 144.940 ;
        RECT 1242.990 96.460 1243.310 96.520 ;
        RECT 1242.795 96.320 1243.310 96.460 ;
        RECT 1242.990 96.260 1243.310 96.320 ;
        RECT 1168.470 51.580 1168.790 51.640 ;
        RECT 1243.005 51.580 1243.295 51.625 ;
        RECT 1168.470 51.440 1243.295 51.580 ;
        RECT 1168.470 51.380 1168.790 51.440 ;
        RECT 1243.005 51.395 1243.295 51.440 ;
      LAYER via ;
        RECT 1244.400 434.900 1244.660 435.160 ;
        RECT 1244.860 434.900 1245.120 435.160 ;
        RECT 1244.400 400.560 1244.660 400.820 ;
        RECT 1243.020 386.280 1243.280 386.540 ;
        RECT 1243.020 351.940 1243.280 352.200 ;
        RECT 1243.020 338.000 1243.280 338.260 ;
        RECT 1243.480 303.660 1243.740 303.920 ;
        RECT 1243.480 302.980 1243.740 303.240 ;
        RECT 1244.860 234.300 1245.120 234.560 ;
        RECT 1244.860 186.360 1245.120 186.620 ;
        RECT 1243.480 144.880 1243.740 145.140 ;
        RECT 1244.860 144.880 1245.120 145.140 ;
        RECT 1243.020 96.260 1243.280 96.520 ;
        RECT 1168.500 51.380 1168.760 51.640 ;
      LAYER met2 ;
        RECT 1248.210 511.090 1248.490 514.000 ;
        RECT 1244.920 510.950 1248.490 511.090 ;
        RECT 1244.920 435.190 1245.060 510.950 ;
        RECT 1248.210 510.000 1248.490 510.950 ;
        RECT 1244.400 434.870 1244.660 435.190 ;
        RECT 1244.860 434.870 1245.120 435.190 ;
        RECT 1244.460 400.850 1244.600 434.870 ;
        RECT 1244.400 400.530 1244.660 400.850 ;
        RECT 1243.020 386.250 1243.280 386.570 ;
        RECT 1243.080 352.230 1243.220 386.250 ;
        RECT 1243.020 351.910 1243.280 352.230 ;
        RECT 1243.020 337.970 1243.280 338.290 ;
        RECT 1243.080 337.690 1243.220 337.970 ;
        RECT 1243.080 337.550 1243.680 337.690 ;
        RECT 1243.540 303.950 1243.680 337.550 ;
        RECT 1243.480 303.630 1243.740 303.950 ;
        RECT 1243.480 302.950 1243.740 303.270 ;
        RECT 1243.540 241.245 1243.680 302.950 ;
        RECT 1243.470 240.875 1243.750 241.245 ;
        RECT 1244.850 240.875 1245.130 241.245 ;
        RECT 1244.920 234.590 1245.060 240.875 ;
        RECT 1244.860 234.270 1245.120 234.590 ;
        RECT 1244.860 186.330 1245.120 186.650 ;
        RECT 1244.920 145.170 1245.060 186.330 ;
        RECT 1243.480 144.850 1243.740 145.170 ;
        RECT 1244.860 144.850 1245.120 145.170 ;
        RECT 1243.540 110.570 1243.680 144.850 ;
        RECT 1243.080 110.430 1243.680 110.570 ;
        RECT 1243.080 96.550 1243.220 110.430 ;
        RECT 1243.020 96.230 1243.280 96.550 ;
        RECT 1168.500 51.350 1168.760 51.670 ;
        RECT 1168.560 2.400 1168.700 51.350 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
      LAYER via2 ;
        RECT 1243.470 240.920 1243.750 241.200 ;
        RECT 1244.850 240.920 1245.130 241.200 ;
      LAYER met3 ;
        RECT 1243.445 241.210 1243.775 241.225 ;
        RECT 1244.825 241.210 1245.155 241.225 ;
        RECT 1243.445 240.910 1245.155 241.210 ;
        RECT 1243.445 240.895 1243.775 240.910 ;
        RECT 1244.825 240.895 1245.155 240.910 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1257.325 421.005 1257.495 469.115 ;
      LAYER mcon ;
        RECT 1257.325 468.945 1257.495 469.115 ;
      LAYER met1 ;
        RECT 1257.265 469.100 1257.555 469.145 ;
        RECT 1257.710 469.100 1258.030 469.160 ;
        RECT 1257.265 468.960 1258.030 469.100 ;
        RECT 1257.265 468.915 1257.555 468.960 ;
        RECT 1257.710 468.900 1258.030 468.960 ;
        RECT 1257.250 421.160 1257.570 421.220 ;
        RECT 1257.055 421.020 1257.570 421.160 ;
        RECT 1257.250 420.960 1257.570 421.020 ;
        RECT 1256.790 337.660 1257.110 337.920 ;
        RECT 1256.880 337.520 1257.020 337.660 ;
        RECT 1257.250 337.520 1257.570 337.580 ;
        RECT 1256.880 337.380 1257.570 337.520 ;
        RECT 1257.250 337.320 1257.570 337.380 ;
        RECT 1256.790 62.460 1257.110 62.520 ;
        RECT 1256.420 62.320 1257.110 62.460 ;
        RECT 1256.420 62.180 1256.560 62.320 ;
        RECT 1256.790 62.260 1257.110 62.320 ;
        RECT 1256.330 61.920 1256.650 62.180 ;
        RECT 1185.950 44.780 1186.270 44.840 ;
        RECT 1256.330 44.780 1256.650 44.840 ;
        RECT 1185.950 44.640 1256.650 44.780 ;
        RECT 1185.950 44.580 1186.270 44.640 ;
        RECT 1256.330 44.580 1256.650 44.640 ;
      LAYER via ;
        RECT 1257.740 468.900 1258.000 469.160 ;
        RECT 1257.280 420.960 1257.540 421.220 ;
        RECT 1256.820 337.660 1257.080 337.920 ;
        RECT 1257.280 337.320 1257.540 337.580 ;
        RECT 1256.820 62.260 1257.080 62.520 ;
        RECT 1256.360 61.920 1256.620 62.180 ;
        RECT 1185.980 44.580 1186.240 44.840 ;
        RECT 1256.360 44.580 1256.620 44.840 ;
      LAYER met2 ;
        RECT 1261.090 511.090 1261.370 514.000 ;
        RECT 1257.800 510.950 1261.370 511.090 ;
        RECT 1257.800 469.190 1257.940 510.950 ;
        RECT 1261.090 510.000 1261.370 510.950 ;
        RECT 1257.740 468.870 1258.000 469.190 ;
        RECT 1257.280 420.930 1257.540 421.250 ;
        RECT 1257.340 362.170 1257.480 420.930 ;
        RECT 1256.880 362.030 1257.480 362.170 ;
        RECT 1256.880 337.950 1257.020 362.030 ;
        RECT 1256.820 337.630 1257.080 337.950 ;
        RECT 1257.280 337.290 1257.540 337.610 ;
        RECT 1257.340 110.570 1257.480 337.290 ;
        RECT 1256.880 110.430 1257.480 110.570 ;
        RECT 1256.880 62.550 1257.020 110.430 ;
        RECT 1256.820 62.230 1257.080 62.550 ;
        RECT 1256.360 61.890 1256.620 62.210 ;
        RECT 1256.420 44.870 1256.560 61.890 ;
        RECT 1185.980 44.550 1186.240 44.870 ;
        RECT 1256.360 44.550 1256.620 44.870 ;
        RECT 1186.040 2.400 1186.180 44.550 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.590 111.220 1270.910 111.480 ;
        RECT 1270.680 110.800 1270.820 111.220 ;
        RECT 1270.590 110.540 1270.910 110.800 ;
        RECT 1203.890 30.840 1204.210 30.900 ;
        RECT 1270.590 30.840 1270.910 30.900 ;
        RECT 1203.890 30.700 1270.910 30.840 ;
        RECT 1203.890 30.640 1204.210 30.700 ;
        RECT 1270.590 30.640 1270.910 30.700 ;
      LAYER via ;
        RECT 1270.620 111.220 1270.880 111.480 ;
        RECT 1270.620 110.540 1270.880 110.800 ;
        RECT 1203.920 30.640 1204.180 30.900 ;
        RECT 1270.620 30.640 1270.880 30.900 ;
      LAYER met2 ;
        RECT 1273.970 510.410 1274.250 514.000 ;
        RECT 1270.220 510.270 1274.250 510.410 ;
        RECT 1270.220 313.890 1270.360 510.270 ;
        RECT 1273.970 510.000 1274.250 510.270 ;
        RECT 1270.220 313.750 1270.820 313.890 ;
        RECT 1270.680 111.510 1270.820 313.750 ;
        RECT 1270.620 111.190 1270.880 111.510 ;
        RECT 1270.620 110.510 1270.880 110.830 ;
        RECT 1270.680 60.250 1270.820 110.510 ;
        RECT 1270.680 60.110 1271.280 60.250 ;
        RECT 1271.140 58.890 1271.280 60.110 ;
        RECT 1270.680 58.750 1271.280 58.890 ;
        RECT 1270.680 30.930 1270.820 58.750 ;
        RECT 1203.920 30.610 1204.180 30.930 ;
        RECT 1270.620 30.610 1270.880 30.930 ;
        RECT 1203.980 2.400 1204.120 30.610 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1222.290 24.040 1222.610 24.100 ;
        RECT 1283.470 24.040 1283.790 24.100 ;
        RECT 1222.290 23.900 1283.790 24.040 ;
        RECT 1222.290 23.840 1222.610 23.900 ;
        RECT 1283.470 23.840 1283.790 23.900 ;
      LAYER via ;
        RECT 1222.320 23.840 1222.580 24.100 ;
        RECT 1283.500 23.840 1283.760 24.100 ;
      LAYER met2 ;
        RECT 1286.850 510.410 1287.130 514.000 ;
        RECT 1283.560 510.270 1287.130 510.410 ;
        RECT 1283.560 24.130 1283.700 510.270 ;
        RECT 1286.850 510.000 1287.130 510.270 ;
        RECT 1222.320 23.810 1222.580 24.130 ;
        RECT 1283.500 23.810 1283.760 24.130 ;
        RECT 1222.380 11.970 1222.520 23.810 ;
        RECT 1221.920 11.830 1222.520 11.970 ;
        RECT 1221.920 2.400 1222.060 11.830 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1239.770 19.960 1240.090 20.020 ;
        RECT 1297.730 19.960 1298.050 20.020 ;
        RECT 1239.770 19.820 1298.050 19.960 ;
        RECT 1239.770 19.760 1240.090 19.820 ;
        RECT 1297.730 19.760 1298.050 19.820 ;
      LAYER via ;
        RECT 1239.800 19.760 1240.060 20.020 ;
        RECT 1297.760 19.760 1298.020 20.020 ;
      LAYER met2 ;
        RECT 1299.270 510.410 1299.550 514.000 ;
        RECT 1297.820 510.270 1299.550 510.410 ;
        RECT 1297.820 20.050 1297.960 510.270 ;
        RECT 1299.270 510.000 1299.550 510.270 ;
        RECT 1239.800 19.730 1240.060 20.050 ;
        RECT 1297.760 19.730 1298.020 20.050 ;
        RECT 1239.860 2.400 1240.000 19.730 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 17.920 1257.570 17.980 ;
        RECT 1311.530 17.920 1311.850 17.980 ;
        RECT 1257.250 17.780 1311.850 17.920 ;
        RECT 1257.250 17.720 1257.570 17.780 ;
        RECT 1311.530 17.720 1311.850 17.780 ;
      LAYER via ;
        RECT 1257.280 17.720 1257.540 17.980 ;
        RECT 1311.560 17.720 1311.820 17.980 ;
      LAYER met2 ;
        RECT 1312.150 510.410 1312.430 514.000 ;
        RECT 1311.620 510.270 1312.430 510.410 ;
        RECT 1311.620 18.010 1311.760 510.270 ;
        RECT 1312.150 510.000 1312.430 510.270 ;
        RECT 1257.280 17.690 1257.540 18.010 ;
        RECT 1311.560 17.690 1311.820 18.010 ;
        RECT 1257.340 2.400 1257.480 17.690 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1275.190 17.240 1275.510 17.300 ;
        RECT 1325.330 17.240 1325.650 17.300 ;
        RECT 1275.190 17.100 1325.650 17.240 ;
        RECT 1275.190 17.040 1275.510 17.100 ;
        RECT 1325.330 17.040 1325.650 17.100 ;
      LAYER via ;
        RECT 1275.220 17.040 1275.480 17.300 ;
        RECT 1325.360 17.040 1325.620 17.300 ;
      LAYER met2 ;
        RECT 1325.030 510.340 1325.310 514.000 ;
        RECT 1324.960 510.000 1325.310 510.340 ;
        RECT 1324.960 473.690 1325.100 510.000 ;
        RECT 1324.960 473.550 1325.560 473.690 ;
        RECT 1325.420 17.330 1325.560 473.550 ;
        RECT 1275.220 17.010 1275.480 17.330 ;
        RECT 1325.360 17.010 1325.620 17.330 ;
        RECT 1275.280 2.400 1275.420 17.010 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1332.305 241.485 1332.475 289.595 ;
      LAYER mcon ;
        RECT 1332.305 289.425 1332.475 289.595 ;
      LAYER met1 ;
        RECT 1333.150 304.200 1333.470 304.260 ;
        RECT 1332.780 304.060 1333.470 304.200 ;
        RECT 1332.780 303.920 1332.920 304.060 ;
        RECT 1333.150 304.000 1333.470 304.060 ;
        RECT 1332.690 303.660 1333.010 303.920 ;
        RECT 1332.245 289.580 1332.535 289.625 ;
        RECT 1332.690 289.580 1333.010 289.640 ;
        RECT 1332.245 289.440 1333.010 289.580 ;
        RECT 1332.245 289.395 1332.535 289.440 ;
        RECT 1332.690 289.380 1333.010 289.440 ;
        RECT 1332.230 241.640 1332.550 241.700 ;
        RECT 1332.035 241.500 1332.550 241.640 ;
        RECT 1332.230 241.440 1332.550 241.500 ;
        RECT 1332.230 193.360 1332.550 193.420 ;
        RECT 1332.690 193.360 1333.010 193.420 ;
        RECT 1332.230 193.220 1333.010 193.360 ;
        RECT 1332.230 193.160 1332.550 193.220 ;
        RECT 1332.690 193.160 1333.010 193.220 ;
        RECT 1293.130 16.560 1293.450 16.620 ;
        RECT 1332.690 16.560 1333.010 16.620 ;
        RECT 1293.130 16.420 1333.010 16.560 ;
        RECT 1293.130 16.360 1293.450 16.420 ;
        RECT 1332.690 16.360 1333.010 16.420 ;
      LAYER via ;
        RECT 1333.180 304.000 1333.440 304.260 ;
        RECT 1332.720 303.660 1332.980 303.920 ;
        RECT 1332.720 289.380 1332.980 289.640 ;
        RECT 1332.260 241.440 1332.520 241.700 ;
        RECT 1332.260 193.160 1332.520 193.420 ;
        RECT 1332.720 193.160 1332.980 193.420 ;
        RECT 1293.160 16.360 1293.420 16.620 ;
        RECT 1332.720 16.360 1332.980 16.620 ;
      LAYER met2 ;
        RECT 1337.910 510.410 1338.190 514.000 ;
        RECT 1335.080 510.270 1338.190 510.410 ;
        RECT 1335.080 449.210 1335.220 510.270 ;
        RECT 1337.910 510.000 1338.190 510.270 ;
        RECT 1334.160 449.070 1335.220 449.210 ;
        RECT 1334.160 400.080 1334.300 449.070 ;
        RECT 1333.240 399.940 1334.300 400.080 ;
        RECT 1333.240 304.290 1333.380 399.940 ;
        RECT 1333.180 303.970 1333.440 304.290 ;
        RECT 1332.720 303.630 1332.980 303.950 ;
        RECT 1332.780 289.670 1332.920 303.630 ;
        RECT 1332.720 289.350 1332.980 289.670 ;
        RECT 1332.260 241.410 1332.520 241.730 ;
        RECT 1332.320 193.450 1332.460 241.410 ;
        RECT 1332.260 193.130 1332.520 193.450 ;
        RECT 1332.720 193.130 1332.980 193.450 ;
        RECT 1332.780 110.570 1332.920 193.130 ;
        RECT 1332.320 110.430 1332.920 110.570 ;
        RECT 1332.320 109.890 1332.460 110.430 ;
        RECT 1332.320 109.750 1332.920 109.890 ;
        RECT 1332.780 16.650 1332.920 109.750 ;
        RECT 1293.160 16.330 1293.420 16.650 ;
        RECT 1332.720 16.330 1332.980 16.650 ;
        RECT 1293.220 2.400 1293.360 16.330 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 19.280 1311.390 19.340 ;
        RECT 1346.490 19.280 1346.810 19.340 ;
        RECT 1311.070 19.140 1346.810 19.280 ;
        RECT 1311.070 19.080 1311.390 19.140 ;
        RECT 1346.490 19.080 1346.810 19.140 ;
      LAYER via ;
        RECT 1311.100 19.080 1311.360 19.340 ;
        RECT 1346.520 19.080 1346.780 19.340 ;
      LAYER met2 ;
        RECT 1350.790 510.410 1351.070 514.000 ;
        RECT 1348.880 510.270 1351.070 510.410 ;
        RECT 1348.880 449.210 1349.020 510.270 ;
        RECT 1350.790 510.000 1351.070 510.270 ;
        RECT 1347.960 449.070 1349.020 449.210 ;
        RECT 1347.960 400.080 1348.100 449.070 ;
        RECT 1347.040 399.940 1348.100 400.080 ;
        RECT 1347.040 304.370 1347.180 399.940 ;
        RECT 1346.580 304.230 1347.180 304.370 ;
        RECT 1346.580 303.690 1346.720 304.230 ;
        RECT 1346.120 303.550 1346.720 303.690 ;
        RECT 1346.120 303.010 1346.260 303.550 ;
        RECT 1346.120 302.870 1346.720 303.010 ;
        RECT 1346.580 207.130 1346.720 302.870 ;
        RECT 1346.120 206.990 1346.720 207.130 ;
        RECT 1346.120 206.450 1346.260 206.990 ;
        RECT 1346.120 206.310 1346.720 206.450 ;
        RECT 1346.580 110.570 1346.720 206.310 ;
        RECT 1346.120 110.430 1346.720 110.570 ;
        RECT 1346.120 109.890 1346.260 110.430 ;
        RECT 1346.120 109.750 1346.720 109.890 ;
        RECT 1346.580 19.370 1346.720 109.750 ;
        RECT 1311.100 19.050 1311.360 19.370 ;
        RECT 1346.520 19.050 1346.780 19.370 ;
        RECT 1311.160 2.400 1311.300 19.050 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1360.365 386.325 1360.535 401.115 ;
        RECT 1359.905 96.645 1360.075 144.755 ;
        RECT 1359.905 15.725 1360.075 48.195 ;
      LAYER mcon ;
        RECT 1360.365 400.945 1360.535 401.115 ;
        RECT 1359.905 144.585 1360.075 144.755 ;
        RECT 1359.905 48.025 1360.075 48.195 ;
      LAYER met1 ;
        RECT 1360.305 401.100 1360.595 401.145 ;
        RECT 1360.750 401.100 1361.070 401.160 ;
        RECT 1360.305 400.960 1361.070 401.100 ;
        RECT 1360.305 400.915 1360.595 400.960 ;
        RECT 1360.750 400.900 1361.070 400.960 ;
        RECT 1360.290 386.480 1360.610 386.540 ;
        RECT 1360.095 386.340 1360.610 386.480 ;
        RECT 1360.290 386.280 1360.610 386.340 ;
        RECT 1359.830 289.920 1360.150 289.980 ;
        RECT 1360.290 289.920 1360.610 289.980 ;
        RECT 1359.830 289.780 1360.610 289.920 ;
        RECT 1359.830 289.720 1360.150 289.780 ;
        RECT 1360.290 289.720 1360.610 289.780 ;
        RECT 1359.830 241.640 1360.150 241.700 ;
        RECT 1360.290 241.640 1360.610 241.700 ;
        RECT 1359.830 241.500 1360.610 241.640 ;
        RECT 1359.830 241.440 1360.150 241.500 ;
        RECT 1360.290 241.440 1360.610 241.500 ;
        RECT 1359.830 217.500 1360.150 217.560 ;
        RECT 1361.210 217.500 1361.530 217.560 ;
        RECT 1359.830 217.360 1361.530 217.500 ;
        RECT 1359.830 217.300 1360.150 217.360 ;
        RECT 1361.210 217.300 1361.530 217.360 ;
        RECT 1358.910 193.020 1359.230 193.080 ;
        RECT 1359.830 193.020 1360.150 193.080 ;
        RECT 1358.910 192.880 1360.150 193.020 ;
        RECT 1358.910 192.820 1359.230 192.880 ;
        RECT 1359.830 192.820 1360.150 192.880 ;
        RECT 1359.830 144.740 1360.150 144.800 ;
        RECT 1359.635 144.600 1360.150 144.740 ;
        RECT 1359.830 144.540 1360.150 144.600 ;
        RECT 1359.830 96.800 1360.150 96.860 ;
        RECT 1359.635 96.660 1360.150 96.800 ;
        RECT 1359.830 96.600 1360.150 96.660 ;
        RECT 1359.830 48.180 1360.150 48.240 ;
        RECT 1359.635 48.040 1360.150 48.180 ;
        RECT 1359.830 47.980 1360.150 48.040 ;
        RECT 1329.010 15.880 1329.330 15.940 ;
        RECT 1359.845 15.880 1360.135 15.925 ;
        RECT 1329.010 15.740 1360.135 15.880 ;
        RECT 1329.010 15.680 1329.330 15.740 ;
        RECT 1359.845 15.695 1360.135 15.740 ;
      LAYER via ;
        RECT 1360.780 400.900 1361.040 401.160 ;
        RECT 1360.320 386.280 1360.580 386.540 ;
        RECT 1359.860 289.720 1360.120 289.980 ;
        RECT 1360.320 289.720 1360.580 289.980 ;
        RECT 1359.860 241.440 1360.120 241.700 ;
        RECT 1360.320 241.440 1360.580 241.700 ;
        RECT 1359.860 217.300 1360.120 217.560 ;
        RECT 1361.240 217.300 1361.500 217.560 ;
        RECT 1358.940 192.820 1359.200 193.080 ;
        RECT 1359.860 192.820 1360.120 193.080 ;
        RECT 1359.860 144.540 1360.120 144.800 ;
        RECT 1359.860 96.600 1360.120 96.860 ;
        RECT 1359.860 47.980 1360.120 48.240 ;
        RECT 1329.040 15.680 1329.300 15.940 ;
      LAYER met2 ;
        RECT 1363.670 510.410 1363.950 514.000 ;
        RECT 1361.300 510.270 1363.950 510.410 ;
        RECT 1361.300 449.210 1361.440 510.270 ;
        RECT 1363.670 510.000 1363.950 510.270 ;
        RECT 1360.840 449.070 1361.440 449.210 ;
        RECT 1360.840 401.190 1360.980 449.070 ;
        RECT 1360.780 400.870 1361.040 401.190 ;
        RECT 1360.320 386.250 1360.580 386.570 ;
        RECT 1360.380 290.010 1360.520 386.250 ;
        RECT 1359.860 289.690 1360.120 290.010 ;
        RECT 1360.320 289.690 1360.580 290.010 ;
        RECT 1359.920 289.410 1360.060 289.690 ;
        RECT 1359.920 289.270 1360.520 289.410 ;
        RECT 1360.380 241.730 1360.520 289.270 ;
        RECT 1359.860 241.410 1360.120 241.730 ;
        RECT 1360.320 241.410 1360.580 241.730 ;
        RECT 1359.920 217.590 1360.060 241.410 ;
        RECT 1359.860 217.270 1360.120 217.590 ;
        RECT 1361.240 217.270 1361.500 217.590 ;
        RECT 1361.300 193.645 1361.440 217.270 ;
        RECT 1360.310 193.530 1360.590 193.645 ;
        RECT 1359.920 193.390 1360.590 193.530 ;
        RECT 1359.920 193.110 1360.060 193.390 ;
        RECT 1360.310 193.275 1360.590 193.390 ;
        RECT 1361.230 193.275 1361.510 193.645 ;
        RECT 1358.940 192.790 1359.200 193.110 ;
        RECT 1359.860 192.790 1360.120 193.110 ;
        RECT 1359.000 145.365 1359.140 192.790 ;
        RECT 1358.930 144.995 1359.210 145.365 ;
        RECT 1359.850 144.995 1360.130 145.365 ;
        RECT 1359.920 144.830 1360.060 144.995 ;
        RECT 1359.860 144.510 1360.120 144.830 ;
        RECT 1359.860 96.570 1360.120 96.890 ;
        RECT 1359.920 48.270 1360.060 96.570 ;
        RECT 1359.860 47.950 1360.120 48.270 ;
        RECT 1329.040 15.650 1329.300 15.970 ;
        RECT 1329.100 2.400 1329.240 15.650 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1360.310 193.320 1360.590 193.600 ;
        RECT 1361.230 193.320 1361.510 193.600 ;
        RECT 1358.930 145.040 1359.210 145.320 ;
        RECT 1359.850 145.040 1360.130 145.320 ;
      LAYER met3 ;
        RECT 1360.285 193.610 1360.615 193.625 ;
        RECT 1361.205 193.610 1361.535 193.625 ;
        RECT 1360.285 193.310 1361.535 193.610 ;
        RECT 1360.285 193.295 1360.615 193.310 ;
        RECT 1361.205 193.295 1361.535 193.310 ;
        RECT 1358.905 145.330 1359.235 145.345 ;
        RECT 1359.825 145.330 1360.155 145.345 ;
        RECT 1358.905 145.030 1360.155 145.330 ;
        RECT 1358.905 145.015 1359.235 145.030 ;
        RECT 1359.825 145.015 1360.155 145.030 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.070 461.960 897.390 462.020 ;
        RECT 900.750 461.960 901.070 462.020 ;
        RECT 897.070 461.820 901.070 461.960 ;
        RECT 897.070 461.760 897.390 461.820 ;
        RECT 900.750 461.760 901.070 461.820 ;
        RECT 689.610 58.720 689.930 58.780 ;
        RECT 897.070 58.720 897.390 58.780 ;
        RECT 689.610 58.580 897.390 58.720 ;
        RECT 689.610 58.520 689.930 58.580 ;
        RECT 897.070 58.520 897.390 58.580 ;
        RECT 686.390 16.900 686.710 16.960 ;
        RECT 689.610 16.900 689.930 16.960 ;
        RECT 686.390 16.760 689.930 16.900 ;
        RECT 686.390 16.700 686.710 16.760 ;
        RECT 689.610 16.700 689.930 16.760 ;
      LAYER via ;
        RECT 897.100 461.760 897.360 462.020 ;
        RECT 900.780 461.760 901.040 462.020 ;
        RECT 689.640 58.520 689.900 58.780 ;
        RECT 897.100 58.520 897.360 58.780 ;
        RECT 686.420 16.700 686.680 16.960 ;
        RECT 689.640 16.700 689.900 16.960 ;
      LAYER met2 ;
        RECT 902.750 510.410 903.030 514.000 ;
        RECT 900.840 510.270 903.030 510.410 ;
        RECT 900.840 462.050 900.980 510.270 ;
        RECT 902.750 510.000 903.030 510.270 ;
        RECT 897.100 461.730 897.360 462.050 ;
        RECT 900.780 461.730 901.040 462.050 ;
        RECT 897.160 58.810 897.300 461.730 ;
        RECT 689.640 58.490 689.900 58.810 ;
        RECT 897.100 58.490 897.360 58.810 ;
        RECT 689.700 16.990 689.840 58.490 ;
        RECT 686.420 16.670 686.680 16.990 ;
        RECT 689.640 16.670 689.900 16.990 ;
        RECT 686.480 2.400 686.620 16.670 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 18.600 1346.810 18.660 ;
        RECT 1373.170 18.600 1373.490 18.660 ;
        RECT 1346.490 18.460 1373.490 18.600 ;
        RECT 1346.490 18.400 1346.810 18.460 ;
        RECT 1373.170 18.400 1373.490 18.460 ;
      LAYER via ;
        RECT 1346.520 18.400 1346.780 18.660 ;
        RECT 1373.200 18.400 1373.460 18.660 ;
      LAYER met2 ;
        RECT 1376.090 510.410 1376.370 514.000 ;
        RECT 1373.260 510.270 1376.370 510.410 ;
        RECT 1373.260 18.690 1373.400 510.270 ;
        RECT 1376.090 510.000 1376.370 510.270 ;
        RECT 1346.520 18.370 1346.780 18.690 ;
        RECT 1373.200 18.370 1373.460 18.690 ;
        RECT 1346.580 2.400 1346.720 18.370 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1364.430 17.580 1364.750 17.640 ;
        RECT 1386.970 17.580 1387.290 17.640 ;
        RECT 1364.430 17.440 1387.290 17.580 ;
        RECT 1364.430 17.380 1364.750 17.440 ;
        RECT 1386.970 17.380 1387.290 17.440 ;
      LAYER via ;
        RECT 1364.460 17.380 1364.720 17.640 ;
        RECT 1387.000 17.380 1387.260 17.640 ;
      LAYER met2 ;
        RECT 1388.970 510.410 1389.250 514.000 ;
        RECT 1387.060 510.270 1389.250 510.410 ;
        RECT 1387.060 17.670 1387.200 510.270 ;
        RECT 1388.970 510.000 1389.250 510.270 ;
        RECT 1364.460 17.350 1364.720 17.670 ;
        RECT 1387.000 17.350 1387.260 17.670 ;
        RECT 1364.520 2.400 1364.660 17.350 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1382.370 18.940 1382.690 19.000 ;
        RECT 1400.770 18.940 1401.090 19.000 ;
        RECT 1382.370 18.800 1401.090 18.940 ;
        RECT 1382.370 18.740 1382.690 18.800 ;
        RECT 1400.770 18.740 1401.090 18.800 ;
      LAYER via ;
        RECT 1382.400 18.740 1382.660 19.000 ;
        RECT 1400.800 18.740 1401.060 19.000 ;
      LAYER met2 ;
        RECT 1401.850 510.410 1402.130 514.000 ;
        RECT 1400.860 510.270 1402.130 510.410 ;
        RECT 1400.860 19.030 1401.000 510.270 ;
        RECT 1401.850 510.000 1402.130 510.270 ;
        RECT 1382.400 18.710 1382.660 19.030 ;
        RECT 1400.800 18.710 1401.060 19.030 ;
        RECT 1382.460 2.400 1382.600 18.710 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 17.240 1400.630 17.300 ;
        RECT 1414.570 17.240 1414.890 17.300 ;
        RECT 1400.310 17.100 1414.890 17.240 ;
        RECT 1400.310 17.040 1400.630 17.100 ;
        RECT 1414.570 17.040 1414.890 17.100 ;
      LAYER via ;
        RECT 1400.340 17.040 1400.600 17.300 ;
        RECT 1414.600 17.040 1414.860 17.300 ;
      LAYER met2 ;
        RECT 1414.730 510.340 1415.010 514.000 ;
        RECT 1414.660 510.000 1415.010 510.340 ;
        RECT 1414.660 17.330 1414.800 510.000 ;
        RECT 1400.340 17.010 1400.600 17.330 ;
        RECT 1414.600 17.010 1414.860 17.330 ;
        RECT 1400.400 2.400 1400.540 17.010 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1422.465 145.265 1422.635 193.035 ;
        RECT 1422.465 96.645 1422.635 144.755 ;
      LAYER mcon ;
        RECT 1422.465 192.865 1422.635 193.035 ;
        RECT 1422.465 144.585 1422.635 144.755 ;
      LAYER met1 ;
        RECT 1422.850 427.960 1423.170 428.020 ;
        RECT 1423.770 427.960 1424.090 428.020 ;
        RECT 1422.850 427.820 1424.090 427.960 ;
        RECT 1422.850 427.760 1423.170 427.820 ;
        RECT 1423.770 427.760 1424.090 427.820 ;
        RECT 1422.850 386.820 1423.170 386.880 ;
        RECT 1422.020 386.680 1423.170 386.820 ;
        RECT 1422.020 386.200 1422.160 386.680 ;
        RECT 1422.850 386.620 1423.170 386.680 ;
        RECT 1421.930 385.940 1422.250 386.200 ;
        RECT 1421.930 338.200 1422.250 338.260 ;
        RECT 1422.390 338.200 1422.710 338.260 ;
        RECT 1421.930 338.060 1422.710 338.200 ;
        RECT 1421.930 338.000 1422.250 338.060 ;
        RECT 1422.390 338.000 1422.710 338.060 ;
        RECT 1422.390 193.020 1422.710 193.080 ;
        RECT 1422.195 192.880 1422.710 193.020 ;
        RECT 1422.390 192.820 1422.710 192.880 ;
        RECT 1422.390 145.420 1422.710 145.480 ;
        RECT 1422.195 145.280 1422.710 145.420 ;
        RECT 1422.390 145.220 1422.710 145.280 ;
        RECT 1422.390 144.740 1422.710 144.800 ;
        RECT 1422.195 144.600 1422.710 144.740 ;
        RECT 1422.390 144.540 1422.710 144.600 ;
        RECT 1422.390 96.800 1422.710 96.860 ;
        RECT 1422.195 96.660 1422.710 96.800 ;
        RECT 1422.390 96.600 1422.710 96.660 ;
        RECT 1418.250 48.180 1418.570 48.240 ;
        RECT 1422.390 48.180 1422.710 48.240 ;
        RECT 1418.250 48.040 1422.710 48.180 ;
        RECT 1418.250 47.980 1418.570 48.040 ;
        RECT 1422.390 47.980 1422.710 48.040 ;
      LAYER via ;
        RECT 1422.880 427.760 1423.140 428.020 ;
        RECT 1423.800 427.760 1424.060 428.020 ;
        RECT 1422.880 386.620 1423.140 386.880 ;
        RECT 1421.960 385.940 1422.220 386.200 ;
        RECT 1421.960 338.000 1422.220 338.260 ;
        RECT 1422.420 338.000 1422.680 338.260 ;
        RECT 1422.420 192.820 1422.680 193.080 ;
        RECT 1422.420 145.220 1422.680 145.480 ;
        RECT 1422.420 144.540 1422.680 144.800 ;
        RECT 1422.420 96.600 1422.680 96.860 ;
        RECT 1418.280 47.980 1418.540 48.240 ;
        RECT 1422.420 47.980 1422.680 48.240 ;
      LAYER met2 ;
        RECT 1427.610 511.090 1427.890 514.000 ;
        RECT 1423.860 510.950 1427.890 511.090 ;
        RECT 1423.860 428.050 1424.000 510.950 ;
        RECT 1427.610 510.000 1427.890 510.950 ;
        RECT 1422.880 427.730 1423.140 428.050 ;
        RECT 1423.800 427.730 1424.060 428.050 ;
        RECT 1422.940 386.910 1423.080 427.730 ;
        RECT 1422.880 386.590 1423.140 386.910 ;
        RECT 1421.960 385.910 1422.220 386.230 ;
        RECT 1422.020 338.290 1422.160 385.910 ;
        RECT 1421.960 337.970 1422.220 338.290 ;
        RECT 1422.420 337.970 1422.680 338.290 ;
        RECT 1422.480 207.130 1422.620 337.970 ;
        RECT 1422.480 206.990 1423.080 207.130 ;
        RECT 1422.940 193.530 1423.080 206.990 ;
        RECT 1422.480 193.390 1423.080 193.530 ;
        RECT 1422.480 193.110 1422.620 193.390 ;
        RECT 1422.420 192.790 1422.680 193.110 ;
        RECT 1422.420 145.190 1422.680 145.510 ;
        RECT 1422.480 144.830 1422.620 145.190 ;
        RECT 1422.420 144.510 1422.680 144.830 ;
        RECT 1422.420 96.570 1422.680 96.890 ;
        RECT 1422.480 48.270 1422.620 96.570 ;
        RECT 1418.280 47.950 1418.540 48.270 ;
        RECT 1422.420 47.950 1422.680 48.270 ;
        RECT 1418.340 2.400 1418.480 47.950 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1436.725 386.325 1436.895 401.115 ;
        RECT 1436.265 282.965 1436.435 331.075 ;
        RECT 1436.265 198.985 1436.435 241.315 ;
        RECT 1436.265 96.645 1436.435 144.755 ;
      LAYER mcon ;
        RECT 1436.725 400.945 1436.895 401.115 ;
        RECT 1436.265 330.905 1436.435 331.075 ;
        RECT 1436.265 241.145 1436.435 241.315 ;
        RECT 1436.265 144.585 1436.435 144.755 ;
      LAYER met1 ;
        RECT 1436.665 401.100 1436.955 401.145 ;
        RECT 1437.110 401.100 1437.430 401.160 ;
        RECT 1436.665 400.960 1437.430 401.100 ;
        RECT 1436.665 400.915 1436.955 400.960 ;
        RECT 1437.110 400.900 1437.430 400.960 ;
        RECT 1436.650 386.480 1436.970 386.540 ;
        RECT 1436.455 386.340 1436.970 386.480 ;
        RECT 1436.650 386.280 1436.970 386.340 ;
        RECT 1436.205 331.060 1436.495 331.105 ;
        RECT 1436.650 331.060 1436.970 331.120 ;
        RECT 1436.205 330.920 1436.970 331.060 ;
        RECT 1436.205 330.875 1436.495 330.920 ;
        RECT 1436.650 330.860 1436.970 330.920 ;
        RECT 1436.190 283.120 1436.510 283.180 ;
        RECT 1435.995 282.980 1436.510 283.120 ;
        RECT 1436.190 282.920 1436.510 282.980 ;
        RECT 1436.190 241.300 1436.510 241.360 ;
        RECT 1435.995 241.160 1436.510 241.300 ;
        RECT 1436.190 241.100 1436.510 241.160 ;
        RECT 1436.190 199.140 1436.510 199.200 ;
        RECT 1435.995 199.000 1436.510 199.140 ;
        RECT 1436.190 198.940 1436.510 199.000 ;
        RECT 1436.190 144.740 1436.510 144.800 ;
        RECT 1435.995 144.600 1436.510 144.740 ;
        RECT 1436.190 144.540 1436.510 144.600 ;
        RECT 1436.205 96.800 1436.495 96.845 ;
        RECT 1436.650 96.800 1436.970 96.860 ;
        RECT 1436.205 96.660 1436.970 96.800 ;
        RECT 1436.205 96.615 1436.495 96.660 ;
        RECT 1436.650 96.600 1436.970 96.660 ;
        RECT 1435.730 2.960 1436.050 3.020 ;
        RECT 1436.650 2.960 1436.970 3.020 ;
        RECT 1435.730 2.820 1436.970 2.960 ;
        RECT 1435.730 2.760 1436.050 2.820 ;
        RECT 1436.650 2.760 1436.970 2.820 ;
      LAYER via ;
        RECT 1437.140 400.900 1437.400 401.160 ;
        RECT 1436.680 386.280 1436.940 386.540 ;
        RECT 1436.680 330.860 1436.940 331.120 ;
        RECT 1436.220 282.920 1436.480 283.180 ;
        RECT 1436.220 241.100 1436.480 241.360 ;
        RECT 1436.220 198.940 1436.480 199.200 ;
        RECT 1436.220 144.540 1436.480 144.800 ;
        RECT 1436.680 96.600 1436.940 96.860 ;
        RECT 1435.760 2.760 1436.020 3.020 ;
        RECT 1436.680 2.760 1436.940 3.020 ;
      LAYER met2 ;
        RECT 1440.490 510.410 1440.770 514.000 ;
        RECT 1439.040 510.270 1440.770 510.410 ;
        RECT 1439.040 449.210 1439.180 510.270 ;
        RECT 1440.490 510.000 1440.770 510.270 ;
        RECT 1437.200 449.070 1439.180 449.210 ;
        RECT 1437.200 401.190 1437.340 449.070 ;
        RECT 1437.140 400.870 1437.400 401.190 ;
        RECT 1436.680 386.250 1436.940 386.570 ;
        RECT 1436.740 331.150 1436.880 386.250 ;
        RECT 1436.680 330.830 1436.940 331.150 ;
        RECT 1436.220 282.890 1436.480 283.210 ;
        RECT 1436.280 241.390 1436.420 282.890 ;
        RECT 1436.220 241.070 1436.480 241.390 ;
        RECT 1436.220 198.910 1436.480 199.230 ;
        RECT 1436.280 144.830 1436.420 198.910 ;
        RECT 1436.220 144.510 1436.480 144.830 ;
        RECT 1436.680 96.570 1436.940 96.890 ;
        RECT 1436.740 3.050 1436.880 96.570 ;
        RECT 1435.760 2.730 1436.020 3.050 ;
        RECT 1436.680 2.730 1436.940 3.050 ;
        RECT 1435.820 2.400 1435.960 2.730 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1450.065 386.325 1450.235 434.775 ;
      LAYER mcon ;
        RECT 1450.065 434.605 1450.235 434.775 ;
      LAYER met1 ;
        RECT 1450.005 434.760 1450.295 434.805 ;
        RECT 1450.450 434.760 1450.770 434.820 ;
        RECT 1450.005 434.620 1450.770 434.760 ;
        RECT 1450.005 434.575 1450.295 434.620 ;
        RECT 1450.450 434.560 1450.770 434.620 ;
        RECT 1449.990 386.480 1450.310 386.540 ;
        RECT 1449.795 386.340 1450.310 386.480 ;
        RECT 1449.990 386.280 1450.310 386.340 ;
        RECT 1449.530 20.640 1449.850 20.700 ;
        RECT 1453.670 20.640 1453.990 20.700 ;
        RECT 1449.530 20.500 1453.990 20.640 ;
        RECT 1449.530 20.440 1449.850 20.500 ;
        RECT 1453.670 20.440 1453.990 20.500 ;
      LAYER via ;
        RECT 1450.480 434.560 1450.740 434.820 ;
        RECT 1450.020 386.280 1450.280 386.540 ;
        RECT 1449.560 20.440 1449.820 20.700 ;
        RECT 1453.700 20.440 1453.960 20.700 ;
      LAYER met2 ;
        RECT 1452.910 510.410 1453.190 514.000 ;
        RECT 1451.000 510.270 1453.190 510.410 ;
        RECT 1451.000 449.210 1451.140 510.270 ;
        RECT 1452.910 510.000 1453.190 510.270 ;
        RECT 1450.540 449.070 1451.140 449.210 ;
        RECT 1450.540 434.850 1450.680 449.070 ;
        RECT 1450.480 434.530 1450.740 434.850 ;
        RECT 1450.020 386.250 1450.280 386.570 ;
        RECT 1450.080 304.370 1450.220 386.250 ;
        RECT 1449.620 304.230 1450.220 304.370 ;
        RECT 1449.620 303.690 1449.760 304.230 ;
        RECT 1449.160 303.550 1449.760 303.690 ;
        RECT 1449.160 303.010 1449.300 303.550 ;
        RECT 1449.160 302.870 1449.760 303.010 ;
        RECT 1449.620 207.130 1449.760 302.870 ;
        RECT 1449.160 206.990 1449.760 207.130 ;
        RECT 1449.160 206.450 1449.300 206.990 ;
        RECT 1449.160 206.310 1449.760 206.450 ;
        RECT 1449.620 110.570 1449.760 206.310 ;
        RECT 1449.160 110.430 1449.760 110.570 ;
        RECT 1449.160 109.890 1449.300 110.430 ;
        RECT 1449.160 109.750 1449.760 109.890 ;
        RECT 1449.620 20.730 1449.760 109.750 ;
        RECT 1449.560 20.410 1449.820 20.730 ;
        RECT 1453.700 20.410 1453.960 20.730 ;
        RECT 1453.760 2.400 1453.900 20.410 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1465.630 496.980 1465.950 497.040 ;
        RECT 1469.310 496.980 1469.630 497.040 ;
        RECT 1465.630 496.840 1469.630 496.980 ;
        RECT 1465.630 496.780 1465.950 496.840 ;
        RECT 1469.310 496.780 1469.630 496.840 ;
        RECT 1469.310 15.880 1469.630 15.940 ;
        RECT 1471.610 15.880 1471.930 15.940 ;
        RECT 1469.310 15.740 1471.930 15.880 ;
        RECT 1469.310 15.680 1469.630 15.740 ;
        RECT 1471.610 15.680 1471.930 15.740 ;
      LAYER via ;
        RECT 1465.660 496.780 1465.920 497.040 ;
        RECT 1469.340 496.780 1469.600 497.040 ;
        RECT 1469.340 15.680 1469.600 15.940 ;
        RECT 1471.640 15.680 1471.900 15.940 ;
      LAYER met2 ;
        RECT 1465.790 510.340 1466.070 514.000 ;
        RECT 1465.720 510.000 1466.070 510.340 ;
        RECT 1465.720 497.070 1465.860 510.000 ;
        RECT 1465.660 496.750 1465.920 497.070 ;
        RECT 1469.340 496.750 1469.600 497.070 ;
        RECT 1469.400 15.970 1469.540 496.750 ;
        RECT 1469.340 15.650 1469.600 15.970 ;
        RECT 1471.640 15.650 1471.900 15.970 ;
        RECT 1471.700 2.400 1471.840 15.650 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1478.510 496.980 1478.830 497.040 ;
        RECT 1483.110 496.980 1483.430 497.040 ;
        RECT 1478.510 496.840 1483.430 496.980 ;
        RECT 1478.510 496.780 1478.830 496.840 ;
        RECT 1483.110 496.780 1483.430 496.840 ;
        RECT 1483.110 20.300 1483.430 20.360 ;
        RECT 1489.550 20.300 1489.870 20.360 ;
        RECT 1483.110 20.160 1489.870 20.300 ;
        RECT 1483.110 20.100 1483.430 20.160 ;
        RECT 1489.550 20.100 1489.870 20.160 ;
      LAYER via ;
        RECT 1478.540 496.780 1478.800 497.040 ;
        RECT 1483.140 496.780 1483.400 497.040 ;
        RECT 1483.140 20.100 1483.400 20.360 ;
        RECT 1489.580 20.100 1489.840 20.360 ;
      LAYER met2 ;
        RECT 1478.670 510.340 1478.950 514.000 ;
        RECT 1478.600 510.000 1478.950 510.340 ;
        RECT 1478.600 497.070 1478.740 510.000 ;
        RECT 1478.540 496.750 1478.800 497.070 ;
        RECT 1483.140 496.750 1483.400 497.070 ;
        RECT 1483.200 20.390 1483.340 496.750 ;
        RECT 1483.140 20.070 1483.400 20.390 ;
        RECT 1489.580 20.070 1489.840 20.390 ;
        RECT 1489.640 2.400 1489.780 20.070 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1491.390 496.980 1491.710 497.040 ;
        RECT 1496.910 496.980 1497.230 497.040 ;
        RECT 1491.390 496.840 1497.230 496.980 ;
        RECT 1491.390 496.780 1491.710 496.840 ;
        RECT 1496.910 496.780 1497.230 496.840 ;
        RECT 1496.910 15.200 1497.230 15.260 ;
        RECT 1507.030 15.200 1507.350 15.260 ;
        RECT 1496.910 15.060 1507.350 15.200 ;
        RECT 1496.910 15.000 1497.230 15.060 ;
        RECT 1507.030 15.000 1507.350 15.060 ;
      LAYER via ;
        RECT 1491.420 496.780 1491.680 497.040 ;
        RECT 1496.940 496.780 1497.200 497.040 ;
        RECT 1496.940 15.000 1497.200 15.260 ;
        RECT 1507.060 15.000 1507.320 15.260 ;
      LAYER met2 ;
        RECT 1491.550 510.340 1491.830 514.000 ;
        RECT 1491.480 510.000 1491.830 510.340 ;
        RECT 1491.480 497.070 1491.620 510.000 ;
        RECT 1491.420 496.750 1491.680 497.070 ;
        RECT 1496.940 496.750 1497.200 497.070 ;
        RECT 1497.000 15.290 1497.140 496.750 ;
        RECT 1496.940 14.970 1497.200 15.290 ;
        RECT 1507.060 14.970 1507.320 15.290 ;
        RECT 1507.120 2.400 1507.260 14.970 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 910.870 472.840 911.190 472.900 ;
        RECT 913.630 472.840 913.950 472.900 ;
        RECT 910.870 472.700 913.950 472.840 ;
        RECT 910.870 472.640 911.190 472.700 ;
        RECT 913.630 472.640 913.950 472.700 ;
        RECT 709.850 65.520 710.170 65.580 ;
        RECT 910.870 65.520 911.190 65.580 ;
        RECT 709.850 65.380 911.190 65.520 ;
        RECT 709.850 65.320 710.170 65.380 ;
        RECT 910.870 65.320 911.190 65.380 ;
        RECT 704.330 16.900 704.650 16.960 ;
        RECT 709.850 16.900 710.170 16.960 ;
        RECT 704.330 16.760 710.170 16.900 ;
        RECT 704.330 16.700 704.650 16.760 ;
        RECT 709.850 16.700 710.170 16.760 ;
      LAYER via ;
        RECT 910.900 472.640 911.160 472.900 ;
        RECT 913.660 472.640 913.920 472.900 ;
        RECT 709.880 65.320 710.140 65.580 ;
        RECT 910.900 65.320 911.160 65.580 ;
        RECT 704.360 16.700 704.620 16.960 ;
        RECT 709.880 16.700 710.140 16.960 ;
      LAYER met2 ;
        RECT 915.170 510.410 915.450 514.000 ;
        RECT 913.720 510.270 915.450 510.410 ;
        RECT 913.720 472.930 913.860 510.270 ;
        RECT 915.170 510.000 915.450 510.270 ;
        RECT 910.900 472.610 911.160 472.930 ;
        RECT 913.660 472.610 913.920 472.930 ;
        RECT 910.960 65.610 911.100 472.610 ;
        RECT 709.880 65.290 710.140 65.610 ;
        RECT 910.900 65.290 911.160 65.610 ;
        RECT 709.940 16.990 710.080 65.290 ;
        RECT 704.360 16.670 704.620 16.990 ;
        RECT 709.880 16.670 710.140 16.990 ;
        RECT 704.420 2.400 704.560 16.670 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1504.270 496.980 1504.590 497.040 ;
        RECT 1510.710 496.980 1511.030 497.040 ;
        RECT 1504.270 496.840 1511.030 496.980 ;
        RECT 1504.270 496.780 1504.590 496.840 ;
        RECT 1510.710 496.780 1511.030 496.840 ;
        RECT 1510.710 15.880 1511.030 15.940 ;
        RECT 1524.970 15.880 1525.290 15.940 ;
        RECT 1510.710 15.740 1525.290 15.880 ;
        RECT 1510.710 15.680 1511.030 15.740 ;
        RECT 1524.970 15.680 1525.290 15.740 ;
      LAYER via ;
        RECT 1504.300 496.780 1504.560 497.040 ;
        RECT 1510.740 496.780 1511.000 497.040 ;
        RECT 1510.740 15.680 1511.000 15.940 ;
        RECT 1525.000 15.680 1525.260 15.940 ;
      LAYER met2 ;
        RECT 1504.430 510.340 1504.710 514.000 ;
        RECT 1504.360 510.000 1504.710 510.340 ;
        RECT 1504.360 497.070 1504.500 510.000 ;
        RECT 1504.300 496.750 1504.560 497.070 ;
        RECT 1510.740 496.750 1511.000 497.070 ;
        RECT 1510.800 15.970 1510.940 496.750 ;
        RECT 1510.740 15.650 1511.000 15.970 ;
        RECT 1525.000 15.650 1525.260 15.970 ;
        RECT 1525.060 2.400 1525.200 15.650 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 19.620 1517.470 19.680 ;
        RECT 1542.910 19.620 1543.230 19.680 ;
        RECT 1517.150 19.480 1543.230 19.620 ;
        RECT 1517.150 19.420 1517.470 19.480 ;
        RECT 1542.910 19.420 1543.230 19.480 ;
      LAYER via ;
        RECT 1517.180 19.420 1517.440 19.680 ;
        RECT 1542.940 19.420 1543.200 19.680 ;
      LAYER met2 ;
        RECT 1517.310 510.340 1517.590 514.000 ;
        RECT 1517.240 510.000 1517.590 510.340 ;
        RECT 1517.240 19.710 1517.380 510.000 ;
        RECT 1517.180 19.390 1517.440 19.710 ;
        RECT 1542.940 19.390 1543.200 19.710 ;
        RECT 1543.000 2.400 1543.140 19.390 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1560.850 17.580 1561.170 17.640 ;
        RECT 1530.950 17.440 1561.170 17.580 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
        RECT 1560.850 17.380 1561.170 17.440 ;
      LAYER via ;
        RECT 1530.980 17.380 1531.240 17.640 ;
        RECT 1560.880 17.380 1561.140 17.640 ;
      LAYER met2 ;
        RECT 1529.730 510.410 1530.010 514.000 ;
        RECT 1529.730 510.270 1531.180 510.410 ;
        RECT 1529.730 510.000 1530.010 510.270 ;
        RECT 1531.040 17.670 1531.180 510.270 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1560.880 17.350 1561.140 17.670 ;
        RECT 1560.940 2.400 1561.080 17.350 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 15.200 1545.530 15.260 ;
        RECT 1578.790 15.200 1579.110 15.260 ;
        RECT 1545.210 15.060 1579.110 15.200 ;
        RECT 1545.210 15.000 1545.530 15.060 ;
        RECT 1578.790 15.000 1579.110 15.060 ;
      LAYER via ;
        RECT 1545.240 15.000 1545.500 15.260 ;
        RECT 1578.820 15.000 1579.080 15.260 ;
      LAYER met2 ;
        RECT 1542.610 510.410 1542.890 514.000 ;
        RECT 1542.610 510.270 1545.440 510.410 ;
        RECT 1542.610 510.000 1542.890 510.270 ;
        RECT 1545.300 15.290 1545.440 510.270 ;
        RECT 1545.240 14.970 1545.500 15.290 ;
        RECT 1578.820 14.970 1579.080 15.290 ;
        RECT 1578.880 2.400 1579.020 14.970 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 19.620 1559.330 19.680 ;
        RECT 1596.270 19.620 1596.590 19.680 ;
        RECT 1559.010 19.480 1596.590 19.620 ;
        RECT 1559.010 19.420 1559.330 19.480 ;
        RECT 1596.270 19.420 1596.590 19.480 ;
      LAYER via ;
        RECT 1559.040 19.420 1559.300 19.680 ;
        RECT 1596.300 19.420 1596.560 19.680 ;
      LAYER met2 ;
        RECT 1555.490 510.410 1555.770 514.000 ;
        RECT 1555.490 510.270 1559.240 510.410 ;
        RECT 1555.490 510.000 1555.770 510.270 ;
        RECT 1559.100 19.710 1559.240 510.270 ;
        RECT 1559.040 19.390 1559.300 19.710 ;
        RECT 1596.300 19.390 1596.560 19.710 ;
        RECT 1596.360 2.400 1596.500 19.390 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1568.210 503.440 1568.530 503.500 ;
        RECT 1572.810 503.440 1573.130 503.500 ;
        RECT 1568.210 503.300 1573.130 503.440 ;
        RECT 1568.210 503.240 1568.530 503.300 ;
        RECT 1572.810 503.240 1573.130 503.300 ;
        RECT 1572.810 20.300 1573.130 20.360 ;
        RECT 1614.210 20.300 1614.530 20.360 ;
        RECT 1572.810 20.160 1614.530 20.300 ;
        RECT 1572.810 20.100 1573.130 20.160 ;
        RECT 1614.210 20.100 1614.530 20.160 ;
      LAYER via ;
        RECT 1568.240 503.240 1568.500 503.500 ;
        RECT 1572.840 503.240 1573.100 503.500 ;
        RECT 1572.840 20.100 1573.100 20.360 ;
        RECT 1614.240 20.100 1614.500 20.360 ;
      LAYER met2 ;
        RECT 1568.370 510.340 1568.650 514.000 ;
        RECT 1568.300 510.000 1568.650 510.340 ;
        RECT 1568.300 503.530 1568.440 510.000 ;
        RECT 1568.240 503.210 1568.500 503.530 ;
        RECT 1572.840 503.210 1573.100 503.530 ;
        RECT 1572.900 20.390 1573.040 503.210 ;
        RECT 1572.840 20.070 1573.100 20.390 ;
        RECT 1614.240 20.070 1614.500 20.390 ;
        RECT 1614.300 2.400 1614.440 20.070 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.090 503.440 1581.410 503.500 ;
        RECT 1586.150 503.440 1586.470 503.500 ;
        RECT 1581.090 503.300 1586.470 503.440 ;
        RECT 1581.090 503.240 1581.410 503.300 ;
        RECT 1586.150 503.240 1586.470 503.300 ;
        RECT 1586.150 23.700 1586.470 23.760 ;
        RECT 1632.150 23.700 1632.470 23.760 ;
        RECT 1586.150 23.560 1632.470 23.700 ;
        RECT 1586.150 23.500 1586.470 23.560 ;
        RECT 1632.150 23.500 1632.470 23.560 ;
      LAYER via ;
        RECT 1581.120 503.240 1581.380 503.500 ;
        RECT 1586.180 503.240 1586.440 503.500 ;
        RECT 1586.180 23.500 1586.440 23.760 ;
        RECT 1632.180 23.500 1632.440 23.760 ;
      LAYER met2 ;
        RECT 1581.250 510.340 1581.530 514.000 ;
        RECT 1581.180 510.000 1581.530 510.340 ;
        RECT 1581.180 503.530 1581.320 510.000 ;
        RECT 1581.120 503.210 1581.380 503.530 ;
        RECT 1586.180 503.210 1586.440 503.530 ;
        RECT 1586.240 23.790 1586.380 503.210 ;
        RECT 1586.180 23.470 1586.440 23.790 ;
        RECT 1632.180 23.470 1632.440 23.790 ;
        RECT 1632.240 2.400 1632.380 23.470 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.970 497.320 1594.290 497.380 ;
        RECT 1631.690 497.320 1632.010 497.380 ;
        RECT 1593.970 497.180 1632.010 497.320 ;
        RECT 1593.970 497.120 1594.290 497.180 ;
        RECT 1631.690 497.120 1632.010 497.180 ;
        RECT 1631.690 27.440 1632.010 27.500 ;
        RECT 1650.090 27.440 1650.410 27.500 ;
        RECT 1631.690 27.300 1650.410 27.440 ;
        RECT 1631.690 27.240 1632.010 27.300 ;
        RECT 1650.090 27.240 1650.410 27.300 ;
      LAYER via ;
        RECT 1594.000 497.120 1594.260 497.380 ;
        RECT 1631.720 497.120 1631.980 497.380 ;
        RECT 1631.720 27.240 1631.980 27.500 ;
        RECT 1650.120 27.240 1650.380 27.500 ;
      LAYER met2 ;
        RECT 1594.130 510.340 1594.410 514.000 ;
        RECT 1594.060 510.000 1594.410 510.340 ;
        RECT 1594.060 497.410 1594.200 510.000 ;
        RECT 1594.000 497.090 1594.260 497.410 ;
        RECT 1631.720 497.090 1631.980 497.410 ;
        RECT 1631.780 27.530 1631.920 497.090 ;
        RECT 1631.720 27.210 1631.980 27.530 ;
        RECT 1650.120 27.210 1650.380 27.530 ;
        RECT 1650.180 2.400 1650.320 27.210 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1605.545 276.165 1605.715 324.275 ;
        RECT 1605.545 138.125 1605.715 186.235 ;
        RECT 1605.545 89.845 1605.715 110.755 ;
        RECT 1605.545 30.685 1605.715 47.855 ;
      LAYER mcon ;
        RECT 1605.545 324.105 1605.715 324.275 ;
        RECT 1605.545 186.065 1605.715 186.235 ;
        RECT 1605.545 110.585 1605.715 110.755 ;
        RECT 1605.545 47.685 1605.715 47.855 ;
      LAYER met1 ;
        RECT 1605.930 476.240 1606.250 476.300 ;
        RECT 1606.850 476.240 1607.170 476.300 ;
        RECT 1605.930 476.100 1607.170 476.240 ;
        RECT 1605.930 476.040 1606.250 476.100 ;
        RECT 1606.850 476.040 1607.170 476.100 ;
        RECT 1605.930 427.960 1606.250 428.020 ;
        RECT 1606.390 427.960 1606.710 428.020 ;
        RECT 1605.930 427.820 1606.710 427.960 ;
        RECT 1605.930 427.760 1606.250 427.820 ;
        RECT 1606.390 427.760 1606.710 427.820 ;
        RECT 1605.930 355.540 1606.250 355.600 ;
        RECT 1606.850 355.540 1607.170 355.600 ;
        RECT 1605.930 355.400 1607.170 355.540 ;
        RECT 1605.930 355.340 1606.250 355.400 ;
        RECT 1606.850 355.340 1607.170 355.400 ;
        RECT 1605.470 324.260 1605.790 324.320 ;
        RECT 1605.275 324.120 1605.790 324.260 ;
        RECT 1605.470 324.060 1605.790 324.120 ;
        RECT 1605.485 276.320 1605.775 276.365 ;
        RECT 1605.930 276.320 1606.250 276.380 ;
        RECT 1605.485 276.180 1606.250 276.320 ;
        RECT 1605.485 276.135 1605.775 276.180 ;
        RECT 1605.930 276.120 1606.250 276.180 ;
        RECT 1605.930 255.580 1606.250 255.640 ;
        RECT 1605.560 255.440 1606.250 255.580 ;
        RECT 1605.560 255.300 1605.700 255.440 ;
        RECT 1605.930 255.380 1606.250 255.440 ;
        RECT 1605.470 255.040 1605.790 255.300 ;
        RECT 1605.485 186.220 1605.775 186.265 ;
        RECT 1605.930 186.220 1606.250 186.280 ;
        RECT 1605.485 186.080 1606.250 186.220 ;
        RECT 1605.485 186.035 1605.775 186.080 ;
        RECT 1605.930 186.020 1606.250 186.080 ;
        RECT 1605.470 138.280 1605.790 138.340 ;
        RECT 1605.275 138.140 1605.790 138.280 ;
        RECT 1605.470 138.080 1605.790 138.140 ;
        RECT 1605.470 110.740 1605.790 110.800 ;
        RECT 1605.275 110.600 1605.790 110.740 ;
        RECT 1605.470 110.540 1605.790 110.600 ;
        RECT 1605.470 90.000 1605.790 90.060 ;
        RECT 1605.275 89.860 1605.790 90.000 ;
        RECT 1605.470 89.800 1605.790 89.860 ;
        RECT 1605.470 47.840 1605.790 47.900 ;
        RECT 1605.275 47.700 1605.790 47.840 ;
        RECT 1605.470 47.640 1605.790 47.700 ;
        RECT 1605.485 30.840 1605.775 30.885 ;
        RECT 1605.485 30.700 1656.300 30.840 ;
        RECT 1605.485 30.655 1605.775 30.700 ;
        RECT 1656.160 30.160 1656.300 30.700 ;
        RECT 1668.030 30.160 1668.350 30.220 ;
        RECT 1656.160 30.020 1668.350 30.160 ;
        RECT 1668.030 29.960 1668.350 30.020 ;
      LAYER via ;
        RECT 1605.960 476.040 1606.220 476.300 ;
        RECT 1606.880 476.040 1607.140 476.300 ;
        RECT 1605.960 427.760 1606.220 428.020 ;
        RECT 1606.420 427.760 1606.680 428.020 ;
        RECT 1605.960 355.340 1606.220 355.600 ;
        RECT 1606.880 355.340 1607.140 355.600 ;
        RECT 1605.500 324.060 1605.760 324.320 ;
        RECT 1605.960 276.120 1606.220 276.380 ;
        RECT 1605.960 255.380 1606.220 255.640 ;
        RECT 1605.500 255.040 1605.760 255.300 ;
        RECT 1605.960 186.020 1606.220 186.280 ;
        RECT 1605.500 138.080 1605.760 138.340 ;
        RECT 1605.500 110.540 1605.760 110.800 ;
        RECT 1605.500 89.800 1605.760 90.060 ;
        RECT 1605.500 47.640 1605.760 47.900 ;
        RECT 1668.060 29.960 1668.320 30.220 ;
      LAYER met2 ;
        RECT 1606.550 510.410 1606.830 514.000 ;
        RECT 1606.020 510.270 1606.830 510.410 ;
        RECT 1606.020 476.330 1606.160 510.270 ;
        RECT 1606.550 510.000 1606.830 510.270 ;
        RECT 1605.960 476.010 1606.220 476.330 ;
        RECT 1606.880 476.010 1607.140 476.330 ;
        RECT 1606.940 475.730 1607.080 476.010 ;
        RECT 1606.020 475.590 1607.080 475.730 ;
        RECT 1606.020 428.050 1606.160 475.590 ;
        RECT 1605.960 427.730 1606.220 428.050 ;
        RECT 1606.420 427.730 1606.680 428.050 ;
        RECT 1606.480 403.650 1606.620 427.730 ;
        RECT 1606.020 403.510 1606.620 403.650 ;
        RECT 1606.020 355.630 1606.160 403.510 ;
        RECT 1605.960 355.310 1606.220 355.630 ;
        RECT 1606.880 355.310 1607.140 355.630 ;
        RECT 1606.940 331.685 1607.080 355.310 ;
        RECT 1605.950 331.570 1606.230 331.685 ;
        RECT 1605.560 331.430 1606.230 331.570 ;
        RECT 1605.560 324.350 1605.700 331.430 ;
        RECT 1605.950 331.315 1606.230 331.430 ;
        RECT 1606.870 331.315 1607.150 331.685 ;
        RECT 1605.500 324.030 1605.760 324.350 ;
        RECT 1605.960 276.090 1606.220 276.410 ;
        RECT 1606.020 255.670 1606.160 276.090 ;
        RECT 1605.960 255.350 1606.220 255.670 ;
        RECT 1605.500 255.010 1605.760 255.330 ;
        RECT 1605.560 234.330 1605.700 255.010 ;
        RECT 1605.950 234.330 1606.230 234.445 ;
        RECT 1605.560 234.190 1606.230 234.330 ;
        RECT 1605.950 234.075 1606.230 234.190 ;
        RECT 1605.950 186.475 1606.230 186.845 ;
        RECT 1606.020 186.310 1606.160 186.475 ;
        RECT 1605.960 185.990 1606.220 186.310 ;
        RECT 1605.500 138.050 1605.760 138.370 ;
        RECT 1605.560 110.830 1605.700 138.050 ;
        RECT 1605.500 110.510 1605.760 110.830 ;
        RECT 1605.500 89.770 1605.760 90.090 ;
        RECT 1605.560 47.930 1605.700 89.770 ;
        RECT 1605.500 47.610 1605.760 47.930 ;
        RECT 1668.060 29.930 1668.320 30.250 ;
        RECT 1668.120 2.400 1668.260 29.930 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
      LAYER via2 ;
        RECT 1605.950 331.360 1606.230 331.640 ;
        RECT 1606.870 331.360 1607.150 331.640 ;
        RECT 1605.950 234.120 1606.230 234.400 ;
        RECT 1605.950 186.520 1606.230 186.800 ;
      LAYER met3 ;
        RECT 1605.925 331.650 1606.255 331.665 ;
        RECT 1606.845 331.650 1607.175 331.665 ;
        RECT 1605.925 331.350 1607.175 331.650 ;
        RECT 1605.925 331.335 1606.255 331.350 ;
        RECT 1606.845 331.335 1607.175 331.350 ;
        RECT 1605.925 234.410 1606.255 234.425 ;
        RECT 1606.590 234.410 1606.970 234.420 ;
        RECT 1605.925 234.110 1606.970 234.410 ;
        RECT 1605.925 234.095 1606.255 234.110 ;
        RECT 1606.590 234.100 1606.970 234.110 ;
        RECT 1605.925 186.810 1606.255 186.825 ;
        RECT 1606.590 186.810 1606.970 186.820 ;
        RECT 1605.925 186.510 1606.970 186.810 ;
        RECT 1605.925 186.495 1606.255 186.510 ;
        RECT 1606.590 186.500 1606.970 186.510 ;
      LAYER via3 ;
        RECT 1606.620 234.100 1606.940 234.420 ;
        RECT 1606.620 186.500 1606.940 186.820 ;
      LAYER met4 ;
        RECT 1606.615 234.095 1606.945 234.425 ;
        RECT 1606.630 186.825 1606.930 234.095 ;
        RECT 1606.615 186.495 1606.945 186.825 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1620.650 37.980 1620.970 38.040 ;
        RECT 1685.510 37.980 1685.830 38.040 ;
        RECT 1620.650 37.840 1685.830 37.980 ;
        RECT 1620.650 37.780 1620.970 37.840 ;
        RECT 1685.510 37.780 1685.830 37.840 ;
      LAYER via ;
        RECT 1620.680 37.780 1620.940 38.040 ;
        RECT 1685.540 37.780 1685.800 38.040 ;
      LAYER met2 ;
        RECT 1619.430 510.410 1619.710 514.000 ;
        RECT 1619.430 510.270 1620.880 510.410 ;
        RECT 1619.430 510.000 1619.710 510.270 ;
        RECT 1620.740 38.070 1620.880 510.270 ;
        RECT 1620.680 37.750 1620.940 38.070 ;
        RECT 1685.540 37.750 1685.800 38.070 ;
        RECT 1685.600 2.400 1685.740 37.750 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 72.320 724.430 72.380 ;
        RECT 924.670 72.320 924.990 72.380 ;
        RECT 724.110 72.180 924.990 72.320 ;
        RECT 724.110 72.120 724.430 72.180 ;
        RECT 924.670 72.120 924.990 72.180 ;
      LAYER via ;
        RECT 724.140 72.120 724.400 72.380 ;
        RECT 924.700 72.120 924.960 72.380 ;
      LAYER met2 ;
        RECT 928.050 510.410 928.330 514.000 ;
        RECT 924.760 510.270 928.330 510.410 ;
        RECT 924.760 72.410 924.900 510.270 ;
        RECT 928.050 510.000 928.330 510.270 ;
        RECT 724.140 72.090 724.400 72.410 ;
        RECT 924.700 72.090 924.960 72.410 ;
        RECT 724.200 16.900 724.340 72.090 ;
        RECT 722.360 16.760 724.340 16.900 ;
        RECT 722.360 2.400 722.500 16.760 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1632.150 500.040 1632.470 500.100 ;
        RECT 1686.890 500.040 1687.210 500.100 ;
        RECT 1632.150 499.900 1687.210 500.040 ;
        RECT 1632.150 499.840 1632.470 499.900 ;
        RECT 1686.890 499.840 1687.210 499.900 ;
        RECT 1686.890 42.740 1687.210 42.800 ;
        RECT 1703.450 42.740 1703.770 42.800 ;
        RECT 1686.890 42.600 1703.770 42.740 ;
        RECT 1686.890 42.540 1687.210 42.600 ;
        RECT 1703.450 42.540 1703.770 42.600 ;
      LAYER via ;
        RECT 1632.180 499.840 1632.440 500.100 ;
        RECT 1686.920 499.840 1687.180 500.100 ;
        RECT 1686.920 42.540 1687.180 42.800 ;
        RECT 1703.480 42.540 1703.740 42.800 ;
      LAYER met2 ;
        RECT 1632.310 510.340 1632.590 514.000 ;
        RECT 1632.240 510.000 1632.590 510.340 ;
        RECT 1632.240 500.130 1632.380 510.000 ;
        RECT 1632.180 499.810 1632.440 500.130 ;
        RECT 1686.920 499.810 1687.180 500.130 ;
        RECT 1686.980 42.830 1687.120 499.810 ;
        RECT 1686.920 42.510 1687.180 42.830 ;
        RECT 1703.480 42.510 1703.740 42.830 ;
        RECT 1703.540 2.400 1703.680 42.510 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1645.030 503.440 1645.350 503.500 ;
        RECT 1648.710 503.440 1649.030 503.500 ;
        RECT 1645.030 503.300 1649.030 503.440 ;
        RECT 1645.030 503.240 1645.350 503.300 ;
        RECT 1648.710 503.240 1649.030 503.300 ;
        RECT 1648.710 51.580 1649.030 51.640 ;
        RECT 1718.170 51.580 1718.490 51.640 ;
        RECT 1648.710 51.440 1718.490 51.580 ;
        RECT 1648.710 51.380 1649.030 51.440 ;
        RECT 1718.170 51.380 1718.490 51.440 ;
      LAYER via ;
        RECT 1645.060 503.240 1645.320 503.500 ;
        RECT 1648.740 503.240 1649.000 503.500 ;
        RECT 1648.740 51.380 1649.000 51.640 ;
        RECT 1718.200 51.380 1718.460 51.640 ;
      LAYER met2 ;
        RECT 1645.190 510.340 1645.470 514.000 ;
        RECT 1645.120 510.000 1645.470 510.340 ;
        RECT 1645.120 503.530 1645.260 510.000 ;
        RECT 1645.060 503.210 1645.320 503.530 ;
        RECT 1648.740 503.210 1649.000 503.530 ;
        RECT 1648.800 51.670 1648.940 503.210 ;
        RECT 1648.740 51.350 1649.000 51.670 ;
        RECT 1718.200 51.350 1718.460 51.670 ;
        RECT 1718.260 16.730 1718.400 51.350 ;
        RECT 1718.260 16.590 1721.620 16.730 ;
        RECT 1721.480 2.400 1721.620 16.590 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1657.910 503.440 1658.230 503.500 ;
        RECT 1666.190 503.440 1666.510 503.500 ;
        RECT 1657.910 503.300 1666.510 503.440 ;
        RECT 1657.910 503.240 1658.230 503.300 ;
        RECT 1666.190 503.240 1666.510 503.300 ;
        RECT 1666.190 30.840 1666.510 30.900 ;
        RECT 1739.330 30.840 1739.650 30.900 ;
        RECT 1666.190 30.700 1739.650 30.840 ;
        RECT 1666.190 30.640 1666.510 30.700 ;
        RECT 1739.330 30.640 1739.650 30.700 ;
      LAYER via ;
        RECT 1657.940 503.240 1658.200 503.500 ;
        RECT 1666.220 503.240 1666.480 503.500 ;
        RECT 1666.220 30.640 1666.480 30.900 ;
        RECT 1739.360 30.640 1739.620 30.900 ;
      LAYER met2 ;
        RECT 1658.070 510.340 1658.350 514.000 ;
        RECT 1658.000 510.000 1658.350 510.340 ;
        RECT 1658.000 503.530 1658.140 510.000 ;
        RECT 1657.940 503.210 1658.200 503.530 ;
        RECT 1666.220 503.210 1666.480 503.530 ;
        RECT 1666.280 30.930 1666.420 503.210 ;
        RECT 1666.220 30.610 1666.480 30.930 ;
        RECT 1739.360 30.610 1739.620 30.930 ;
        RECT 1739.420 2.400 1739.560 30.610 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1670.790 503.440 1671.110 503.500 ;
        RECT 1676.310 503.440 1676.630 503.500 ;
        RECT 1670.790 503.300 1676.630 503.440 ;
        RECT 1670.790 503.240 1671.110 503.300 ;
        RECT 1676.310 503.240 1676.630 503.300 ;
        RECT 1676.310 24.040 1676.630 24.100 ;
        RECT 1756.810 24.040 1757.130 24.100 ;
        RECT 1676.310 23.900 1757.130 24.040 ;
        RECT 1676.310 23.840 1676.630 23.900 ;
        RECT 1756.810 23.840 1757.130 23.900 ;
      LAYER via ;
        RECT 1670.820 503.240 1671.080 503.500 ;
        RECT 1676.340 503.240 1676.600 503.500 ;
        RECT 1676.340 23.840 1676.600 24.100 ;
        RECT 1756.840 23.840 1757.100 24.100 ;
      LAYER met2 ;
        RECT 1670.950 510.340 1671.230 514.000 ;
        RECT 1670.880 510.000 1671.230 510.340 ;
        RECT 1670.880 503.530 1671.020 510.000 ;
        RECT 1670.820 503.210 1671.080 503.530 ;
        RECT 1676.340 503.210 1676.600 503.530 ;
        RECT 1676.400 24.130 1676.540 503.210 ;
        RECT 1676.340 23.810 1676.600 24.130 ;
        RECT 1756.840 23.810 1757.100 24.130 ;
        RECT 1756.900 2.400 1757.040 23.810 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 493.240 1683.530 493.300 ;
        RECT 1773.370 493.240 1773.690 493.300 ;
        RECT 1683.210 493.100 1773.690 493.240 ;
        RECT 1683.210 493.040 1683.530 493.100 ;
        RECT 1773.370 493.040 1773.690 493.100 ;
      LAYER via ;
        RECT 1683.240 493.040 1683.500 493.300 ;
        RECT 1773.400 493.040 1773.660 493.300 ;
      LAYER met2 ;
        RECT 1683.370 510.340 1683.650 514.000 ;
        RECT 1683.300 510.000 1683.650 510.340 ;
        RECT 1683.300 493.330 1683.440 510.000 ;
        RECT 1683.240 493.010 1683.500 493.330 ;
        RECT 1773.400 493.010 1773.660 493.330 ;
        RECT 1773.460 5.170 1773.600 493.010 ;
        RECT 1773.460 5.030 1774.980 5.170 ;
        RECT 1774.840 2.400 1774.980 5.030 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1792.765 2.805 1792.935 48.195 ;
      LAYER mcon ;
        RECT 1792.765 48.025 1792.935 48.195 ;
      LAYER met1 ;
        RECT 1696.090 497.660 1696.410 497.720 ;
        RECT 1721.390 497.660 1721.710 497.720 ;
        RECT 1696.090 497.520 1721.710 497.660 ;
        RECT 1696.090 497.460 1696.410 497.520 ;
        RECT 1721.390 497.460 1721.710 497.520 ;
        RECT 1721.390 72.320 1721.710 72.380 ;
        RECT 1787.170 72.320 1787.490 72.380 ;
        RECT 1721.390 72.180 1787.490 72.320 ;
        RECT 1721.390 72.120 1721.710 72.180 ;
        RECT 1787.170 72.120 1787.490 72.180 ;
        RECT 1787.170 48.180 1787.490 48.240 ;
        RECT 1792.705 48.180 1792.995 48.225 ;
        RECT 1787.170 48.040 1792.995 48.180 ;
        RECT 1787.170 47.980 1787.490 48.040 ;
        RECT 1792.705 47.995 1792.995 48.040 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1792.495 2.820 1793.010 2.960 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
      LAYER via ;
        RECT 1696.120 497.460 1696.380 497.720 ;
        RECT 1721.420 497.460 1721.680 497.720 ;
        RECT 1721.420 72.120 1721.680 72.380 ;
        RECT 1787.200 72.120 1787.460 72.380 ;
        RECT 1787.200 47.980 1787.460 48.240 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
      LAYER met2 ;
        RECT 1696.250 510.340 1696.530 514.000 ;
        RECT 1696.180 510.000 1696.530 510.340 ;
        RECT 1696.180 497.750 1696.320 510.000 ;
        RECT 1696.120 497.430 1696.380 497.750 ;
        RECT 1721.420 497.430 1721.680 497.750 ;
        RECT 1721.480 72.410 1721.620 497.430 ;
        RECT 1721.420 72.090 1721.680 72.410 ;
        RECT 1787.200 72.090 1787.460 72.410 ;
        RECT 1787.260 48.270 1787.400 72.090 ;
        RECT 1787.200 47.950 1787.460 48.270 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.350 369.140 1710.670 369.200 ;
        RECT 1807.870 369.140 1808.190 369.200 ;
        RECT 1710.350 369.000 1808.190 369.140 ;
        RECT 1710.350 368.940 1710.670 369.000 ;
        RECT 1807.870 368.940 1808.190 369.000 ;
      LAYER via ;
        RECT 1710.380 368.940 1710.640 369.200 ;
        RECT 1807.900 368.940 1808.160 369.200 ;
      LAYER met2 ;
        RECT 1709.130 510.410 1709.410 514.000 ;
        RECT 1709.130 510.270 1710.580 510.410 ;
        RECT 1709.130 510.000 1709.410 510.270 ;
        RECT 1710.440 369.230 1710.580 510.270 ;
        RECT 1710.380 368.910 1710.640 369.230 ;
        RECT 1807.900 368.910 1808.160 369.230 ;
        RECT 1807.960 16.050 1808.100 368.910 ;
        RECT 1807.960 15.910 1810.860 16.050 ;
        RECT 1810.720 2.400 1810.860 15.910 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 37.980 1724.930 38.040 ;
        RECT 1829.030 37.980 1829.350 38.040 ;
        RECT 1724.610 37.840 1829.350 37.980 ;
        RECT 1724.610 37.780 1724.930 37.840 ;
        RECT 1829.030 37.780 1829.350 37.840 ;
      LAYER via ;
        RECT 1724.640 37.780 1724.900 38.040 ;
        RECT 1829.060 37.780 1829.320 38.040 ;
      LAYER met2 ;
        RECT 1722.010 510.410 1722.290 514.000 ;
        RECT 1722.010 510.270 1724.840 510.410 ;
        RECT 1722.010 510.000 1722.290 510.270 ;
        RECT 1724.700 38.070 1724.840 510.270 ;
        RECT 1724.640 37.750 1724.900 38.070 ;
        RECT 1829.060 37.750 1829.320 38.070 ;
        RECT 1829.120 17.410 1829.260 37.750 ;
        RECT 1828.660 17.270 1829.260 17.410 ;
        RECT 1828.660 2.400 1828.800 17.270 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1734.730 500.040 1735.050 500.100 ;
        RECT 1842.830 500.040 1843.150 500.100 ;
        RECT 1734.730 499.900 1843.150 500.040 ;
        RECT 1734.730 499.840 1735.050 499.900 ;
        RECT 1842.830 499.840 1843.150 499.900 ;
      LAYER via ;
        RECT 1734.760 499.840 1735.020 500.100 ;
        RECT 1842.860 499.840 1843.120 500.100 ;
      LAYER met2 ;
        RECT 1734.890 510.340 1735.170 514.000 ;
        RECT 1734.820 510.000 1735.170 510.340 ;
        RECT 1734.820 500.130 1734.960 510.000 ;
        RECT 1734.760 499.810 1735.020 500.130 ;
        RECT 1842.860 499.810 1843.120 500.130 ;
        RECT 1842.920 17.410 1843.060 499.810 ;
        RECT 1842.920 17.270 1846.280 17.410 ;
        RECT 1846.140 2.400 1846.280 17.270 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1747.610 486.440 1747.930 486.500 ;
        RECT 1747.610 486.300 1833.400 486.440 ;
        RECT 1747.610 486.240 1747.930 486.300 ;
        RECT 1833.260 486.100 1833.400 486.300 ;
        RECT 1863.070 486.100 1863.390 486.160 ;
        RECT 1833.260 485.960 1863.390 486.100 ;
        RECT 1863.070 485.900 1863.390 485.960 ;
      LAYER via ;
        RECT 1747.640 486.240 1747.900 486.500 ;
        RECT 1863.100 485.900 1863.360 486.160 ;
      LAYER met2 ;
        RECT 1747.770 510.340 1748.050 514.000 ;
        RECT 1747.700 510.000 1748.050 510.340 ;
        RECT 1747.700 486.530 1747.840 510.000 ;
        RECT 1747.640 486.210 1747.900 486.530 ;
        RECT 1863.100 485.870 1863.360 486.190 ;
        RECT 1863.160 17.410 1863.300 485.870 ;
        RECT 1863.160 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 927.890 496.980 928.210 497.040 ;
        RECT 940.770 496.980 941.090 497.040 ;
        RECT 927.890 496.840 941.090 496.980 ;
        RECT 927.890 496.780 928.210 496.840 ;
        RECT 940.770 496.780 941.090 496.840 ;
        RECT 744.810 79.460 745.130 79.520 ;
        RECT 927.890 79.460 928.210 79.520 ;
        RECT 744.810 79.320 928.210 79.460 ;
        RECT 744.810 79.260 745.130 79.320 ;
        RECT 927.890 79.260 928.210 79.320 ;
        RECT 740.210 15.880 740.530 15.940 ;
        RECT 744.810 15.880 745.130 15.940 ;
        RECT 740.210 15.740 745.130 15.880 ;
        RECT 740.210 15.680 740.530 15.740 ;
        RECT 744.810 15.680 745.130 15.740 ;
      LAYER via ;
        RECT 927.920 496.780 928.180 497.040 ;
        RECT 940.800 496.780 941.060 497.040 ;
        RECT 744.840 79.260 745.100 79.520 ;
        RECT 927.920 79.260 928.180 79.520 ;
        RECT 740.240 15.680 740.500 15.940 ;
        RECT 744.840 15.680 745.100 15.940 ;
      LAYER met2 ;
        RECT 940.930 510.340 941.210 514.000 ;
        RECT 940.860 510.000 941.210 510.340 ;
        RECT 940.860 497.070 941.000 510.000 ;
        RECT 927.920 496.750 928.180 497.070 ;
        RECT 940.800 496.750 941.060 497.070 ;
        RECT 927.980 79.550 928.120 496.750 ;
        RECT 744.840 79.230 745.100 79.550 ;
        RECT 927.920 79.230 928.180 79.550 ;
        RECT 744.900 15.970 745.040 79.230 ;
        RECT 740.240 15.650 740.500 15.970 ;
        RECT 744.840 15.650 745.100 15.970 ;
        RECT 740.300 2.400 740.440 15.650 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1760.030 503.100 1760.350 503.160 ;
        RECT 1766.010 503.100 1766.330 503.160 ;
        RECT 1760.030 502.960 1766.330 503.100 ;
        RECT 1760.030 502.900 1760.350 502.960 ;
        RECT 1766.010 502.900 1766.330 502.960 ;
        RECT 1766.010 24.040 1766.330 24.100 ;
        RECT 1881.930 24.040 1882.250 24.100 ;
        RECT 1766.010 23.900 1882.250 24.040 ;
        RECT 1766.010 23.840 1766.330 23.900 ;
        RECT 1881.930 23.840 1882.250 23.900 ;
      LAYER via ;
        RECT 1760.060 502.900 1760.320 503.160 ;
        RECT 1766.040 502.900 1766.300 503.160 ;
        RECT 1766.040 23.840 1766.300 24.100 ;
        RECT 1881.960 23.840 1882.220 24.100 ;
      LAYER met2 ;
        RECT 1760.190 510.340 1760.470 514.000 ;
        RECT 1760.120 510.000 1760.470 510.340 ;
        RECT 1760.120 503.190 1760.260 510.000 ;
        RECT 1760.060 502.870 1760.320 503.190 ;
        RECT 1766.040 502.870 1766.300 503.190 ;
        RECT 1766.100 24.130 1766.240 502.870 ;
        RECT 1766.040 23.810 1766.300 24.130 ;
        RECT 1881.960 23.810 1882.220 24.130 ;
        RECT 1882.020 2.400 1882.160 23.810 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.450 479.640 1772.770 479.700 ;
        RECT 1897.570 479.640 1897.890 479.700 ;
        RECT 1772.450 479.500 1897.890 479.640 ;
        RECT 1772.450 479.440 1772.770 479.500 ;
        RECT 1897.570 479.440 1897.890 479.500 ;
      LAYER via ;
        RECT 1772.480 479.440 1772.740 479.700 ;
        RECT 1897.600 479.440 1897.860 479.700 ;
      LAYER met2 ;
        RECT 1773.070 510.410 1773.350 514.000 ;
        RECT 1772.540 510.270 1773.350 510.410 ;
        RECT 1772.540 479.730 1772.680 510.270 ;
        RECT 1773.070 510.000 1773.350 510.270 ;
        RECT 1772.480 479.410 1772.740 479.730 ;
        RECT 1897.600 479.410 1897.860 479.730 ;
        RECT 1897.660 16.730 1897.800 479.410 ;
        RECT 1897.660 16.590 1900.100 16.730 ;
        RECT 1899.960 2.400 1900.100 16.590 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1784.945 282.965 1785.115 331.075 ;
        RECT 1785.405 158.525 1785.575 186.235 ;
        RECT 1785.865 89.845 1786.035 137.955 ;
      LAYER mcon ;
        RECT 1784.945 330.905 1785.115 331.075 ;
        RECT 1785.405 186.065 1785.575 186.235 ;
        RECT 1785.865 137.785 1786.035 137.955 ;
      LAYER met1 ;
        RECT 1784.410 483.380 1784.730 483.440 ;
        RECT 1784.870 483.380 1785.190 483.440 ;
        RECT 1784.410 483.240 1785.190 483.380 ;
        RECT 1784.410 483.180 1784.730 483.240 ;
        RECT 1784.870 483.180 1785.190 483.240 ;
        RECT 1785.330 400.900 1785.650 401.160 ;
        RECT 1785.420 400.140 1785.560 400.900 ;
        RECT 1785.330 399.880 1785.650 400.140 ;
        RECT 1784.870 331.060 1785.190 331.120 ;
        RECT 1784.675 330.920 1785.190 331.060 ;
        RECT 1784.870 330.860 1785.190 330.920 ;
        RECT 1784.885 283.120 1785.175 283.165 ;
        RECT 1785.330 283.120 1785.650 283.180 ;
        RECT 1784.885 282.980 1785.650 283.120 ;
        RECT 1784.885 282.935 1785.175 282.980 ;
        RECT 1785.330 282.920 1785.650 282.980 ;
        RECT 1784.870 207.100 1785.190 207.360 ;
        RECT 1784.960 206.620 1785.100 207.100 ;
        RECT 1785.330 206.620 1785.650 206.680 ;
        RECT 1784.960 206.480 1785.650 206.620 ;
        RECT 1785.330 206.420 1785.650 206.480 ;
        RECT 1785.330 186.220 1785.650 186.280 ;
        RECT 1785.135 186.080 1785.650 186.220 ;
        RECT 1785.330 186.020 1785.650 186.080 ;
        RECT 1785.330 158.680 1785.650 158.740 ;
        RECT 1785.135 158.540 1785.650 158.680 ;
        RECT 1785.330 158.480 1785.650 158.540 ;
        RECT 1785.790 137.940 1786.110 138.000 ;
        RECT 1785.595 137.800 1786.110 137.940 ;
        RECT 1785.790 137.740 1786.110 137.800 ;
        RECT 1785.805 90.000 1786.095 90.045 ;
        RECT 1786.250 90.000 1786.570 90.060 ;
        RECT 1785.805 89.860 1786.570 90.000 ;
        RECT 1785.805 89.815 1786.095 89.860 ;
        RECT 1786.250 89.800 1786.570 89.860 ;
        RECT 1785.790 30.840 1786.110 30.900 ;
        RECT 1917.350 30.840 1917.670 30.900 ;
        RECT 1785.790 30.700 1917.670 30.840 ;
        RECT 1785.790 30.640 1786.110 30.700 ;
        RECT 1917.350 30.640 1917.670 30.700 ;
      LAYER via ;
        RECT 1784.440 483.180 1784.700 483.440 ;
        RECT 1784.900 483.180 1785.160 483.440 ;
        RECT 1785.360 400.900 1785.620 401.160 ;
        RECT 1785.360 399.880 1785.620 400.140 ;
        RECT 1784.900 330.860 1785.160 331.120 ;
        RECT 1785.360 282.920 1785.620 283.180 ;
        RECT 1784.900 207.100 1785.160 207.360 ;
        RECT 1785.360 206.420 1785.620 206.680 ;
        RECT 1785.360 186.020 1785.620 186.280 ;
        RECT 1785.360 158.480 1785.620 158.740 ;
        RECT 1785.820 137.740 1786.080 138.000 ;
        RECT 1786.280 89.800 1786.540 90.060 ;
        RECT 1785.820 30.640 1786.080 30.900 ;
        RECT 1917.380 30.640 1917.640 30.900 ;
      LAYER met2 ;
        RECT 1785.950 511.090 1786.230 514.000 ;
        RECT 1784.500 510.950 1786.230 511.090 ;
        RECT 1784.500 483.470 1784.640 510.950 ;
        RECT 1785.950 510.000 1786.230 510.950 ;
        RECT 1784.440 483.150 1784.700 483.470 ;
        RECT 1784.900 483.150 1785.160 483.470 ;
        RECT 1784.960 448.530 1785.100 483.150 ;
        RECT 1784.960 448.390 1785.560 448.530 ;
        RECT 1785.420 401.190 1785.560 448.390 ;
        RECT 1785.360 400.870 1785.620 401.190 ;
        RECT 1785.360 399.850 1785.620 400.170 ;
        RECT 1785.420 338.370 1785.560 399.850 ;
        RECT 1784.960 338.230 1785.560 338.370 ;
        RECT 1784.960 331.150 1785.100 338.230 ;
        RECT 1784.900 330.830 1785.160 331.150 ;
        RECT 1785.360 282.890 1785.620 283.210 ;
        RECT 1785.420 254.730 1785.560 282.890 ;
        RECT 1784.960 254.590 1785.560 254.730 ;
        RECT 1784.960 207.390 1785.100 254.590 ;
        RECT 1784.900 207.070 1785.160 207.390 ;
        RECT 1785.360 206.390 1785.620 206.710 ;
        RECT 1785.420 186.310 1785.560 206.390 ;
        RECT 1785.360 185.990 1785.620 186.310 ;
        RECT 1785.360 158.450 1785.620 158.770 ;
        RECT 1785.420 138.450 1785.560 158.450 ;
        RECT 1785.420 138.310 1786.020 138.450 ;
        RECT 1785.880 138.030 1786.020 138.310 ;
        RECT 1785.820 137.710 1786.080 138.030 ;
        RECT 1786.280 89.770 1786.540 90.090 ;
        RECT 1786.340 62.290 1786.480 89.770 ;
        RECT 1785.880 62.150 1786.480 62.290 ;
        RECT 1785.880 30.930 1786.020 62.150 ;
        RECT 1785.820 30.610 1786.080 30.930 ;
        RECT 1917.380 30.610 1917.640 30.930 ;
        RECT 1917.440 30.330 1917.580 30.610 ;
        RECT 1917.440 30.190 1918.040 30.330 ;
        RECT 1917.900 2.400 1918.040 30.190 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.050 44.780 1800.370 44.840 ;
        RECT 1935.290 44.780 1935.610 44.840 ;
        RECT 1800.050 44.640 1935.610 44.780 ;
        RECT 1800.050 44.580 1800.370 44.640 ;
        RECT 1935.290 44.580 1935.610 44.640 ;
      LAYER via ;
        RECT 1800.080 44.580 1800.340 44.840 ;
        RECT 1935.320 44.580 1935.580 44.840 ;
      LAYER met2 ;
        RECT 1798.830 510.410 1799.110 514.000 ;
        RECT 1798.830 510.270 1800.280 510.410 ;
        RECT 1798.830 510.000 1799.110 510.270 ;
        RECT 1800.140 44.870 1800.280 510.270 ;
        RECT 1800.080 44.550 1800.340 44.870 ;
        RECT 1935.320 44.550 1935.580 44.870 ;
        RECT 1935.380 2.400 1935.520 44.550 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 51.580 1814.630 51.640 ;
        RECT 1953.230 51.580 1953.550 51.640 ;
        RECT 1814.310 51.440 1953.550 51.580 ;
        RECT 1814.310 51.380 1814.630 51.440 ;
        RECT 1953.230 51.380 1953.550 51.440 ;
      LAYER via ;
        RECT 1814.340 51.380 1814.600 51.640 ;
        RECT 1953.260 51.380 1953.520 51.640 ;
      LAYER met2 ;
        RECT 1811.710 510.410 1811.990 514.000 ;
        RECT 1811.710 510.270 1814.540 510.410 ;
        RECT 1811.710 510.000 1811.990 510.270 ;
        RECT 1814.400 51.670 1814.540 510.270 ;
        RECT 1814.340 51.350 1814.600 51.670 ;
        RECT 1953.260 51.350 1953.520 51.670 ;
        RECT 1953.320 2.400 1953.460 51.350 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.430 496.980 1824.750 497.040 ;
        RECT 1828.110 496.980 1828.430 497.040 ;
        RECT 1824.430 496.840 1828.430 496.980 ;
        RECT 1824.430 496.780 1824.750 496.840 ;
        RECT 1828.110 496.780 1828.430 496.840 ;
        RECT 1828.110 58.720 1828.430 58.780 ;
        RECT 1971.170 58.720 1971.490 58.780 ;
        RECT 1828.110 58.580 1971.490 58.720 ;
        RECT 1828.110 58.520 1828.430 58.580 ;
        RECT 1971.170 58.520 1971.490 58.580 ;
      LAYER via ;
        RECT 1824.460 496.780 1824.720 497.040 ;
        RECT 1828.140 496.780 1828.400 497.040 ;
        RECT 1828.140 58.520 1828.400 58.780 ;
        RECT 1971.200 58.520 1971.460 58.780 ;
      LAYER met2 ;
        RECT 1824.590 510.340 1824.870 514.000 ;
        RECT 1824.520 510.000 1824.870 510.340 ;
        RECT 1824.520 497.070 1824.660 510.000 ;
        RECT 1824.460 496.750 1824.720 497.070 ;
        RECT 1828.140 496.750 1828.400 497.070 ;
        RECT 1828.200 58.810 1828.340 496.750 ;
        RECT 1828.140 58.490 1828.400 58.810 ;
        RECT 1971.200 58.490 1971.460 58.810 ;
        RECT 1971.260 2.400 1971.400 58.490 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1837.310 493.240 1837.630 493.300 ;
        RECT 1987.270 493.240 1987.590 493.300 ;
        RECT 1837.310 493.100 1987.590 493.240 ;
        RECT 1837.310 493.040 1837.630 493.100 ;
        RECT 1987.270 493.040 1987.590 493.100 ;
        RECT 1987.730 61.780 1988.050 61.840 ;
        RECT 1989.110 61.780 1989.430 61.840 ;
        RECT 1987.730 61.640 1989.430 61.780 ;
        RECT 1987.730 61.580 1988.050 61.640 ;
        RECT 1989.110 61.580 1989.430 61.640 ;
        RECT 1989.110 47.980 1989.430 48.240 ;
        RECT 1989.200 47.560 1989.340 47.980 ;
        RECT 1989.110 47.300 1989.430 47.560 ;
      LAYER via ;
        RECT 1837.340 493.040 1837.600 493.300 ;
        RECT 1987.300 493.040 1987.560 493.300 ;
        RECT 1987.760 61.580 1988.020 61.840 ;
        RECT 1989.140 61.580 1989.400 61.840 ;
        RECT 1989.140 47.980 1989.400 48.240 ;
        RECT 1989.140 47.300 1989.400 47.560 ;
      LAYER met2 ;
        RECT 1837.470 510.340 1837.750 514.000 ;
        RECT 1837.400 510.000 1837.750 510.340 ;
        RECT 1837.400 493.330 1837.540 510.000 ;
        RECT 1837.340 493.010 1837.600 493.330 ;
        RECT 1987.300 493.010 1987.560 493.330 ;
        RECT 1987.360 72.490 1987.500 493.010 ;
        RECT 1987.360 72.350 1987.960 72.490 ;
        RECT 1987.820 61.870 1987.960 72.350 ;
        RECT 1987.760 61.550 1988.020 61.870 ;
        RECT 1989.140 61.550 1989.400 61.870 ;
        RECT 1989.200 48.270 1989.340 61.550 ;
        RECT 1989.140 47.950 1989.400 48.270 ;
        RECT 1989.140 47.270 1989.400 47.590 ;
        RECT 1989.200 2.400 1989.340 47.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1849.730 502.760 1850.050 502.820 ;
        RECT 1880.090 502.760 1880.410 502.820 ;
        RECT 1849.730 502.620 1880.410 502.760 ;
        RECT 1849.730 502.560 1850.050 502.620 ;
        RECT 1880.090 502.560 1880.410 502.620 ;
        RECT 1880.090 24.380 1880.410 24.440 ;
        RECT 2006.590 24.380 2006.910 24.440 ;
        RECT 1880.090 24.240 2006.910 24.380 ;
        RECT 1880.090 24.180 1880.410 24.240 ;
        RECT 2006.590 24.180 2006.910 24.240 ;
      LAYER via ;
        RECT 1849.760 502.560 1850.020 502.820 ;
        RECT 1880.120 502.560 1880.380 502.820 ;
        RECT 1880.120 24.180 1880.380 24.440 ;
        RECT 2006.620 24.180 2006.880 24.440 ;
      LAYER met2 ;
        RECT 1849.890 510.340 1850.170 514.000 ;
        RECT 1849.820 510.000 1850.170 510.340 ;
        RECT 1849.820 502.850 1849.960 510.000 ;
        RECT 1849.760 502.530 1850.020 502.850 ;
        RECT 1880.120 502.530 1880.380 502.850 ;
        RECT 1880.180 24.470 1880.320 502.530 ;
        RECT 1880.120 24.150 1880.380 24.470 ;
        RECT 2006.620 24.150 2006.880 24.470 ;
        RECT 2006.680 2.400 2006.820 24.150 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1863.070 486.580 1863.390 486.840 ;
        RECT 1863.160 486.440 1863.300 486.580 ;
        RECT 2021.770 486.440 2022.090 486.500 ;
        RECT 1863.160 486.300 2022.090 486.440 ;
        RECT 2021.770 486.240 2022.090 486.300 ;
        RECT 2021.770 62.120 2022.090 62.180 ;
        RECT 2024.530 62.120 2024.850 62.180 ;
        RECT 2021.770 61.980 2024.850 62.120 ;
        RECT 2021.770 61.920 2022.090 61.980 ;
        RECT 2024.530 61.920 2024.850 61.980 ;
      LAYER via ;
        RECT 1863.100 486.580 1863.360 486.840 ;
        RECT 2021.800 486.240 2022.060 486.500 ;
        RECT 2021.800 61.920 2022.060 62.180 ;
        RECT 2024.560 61.920 2024.820 62.180 ;
      LAYER met2 ;
        RECT 1862.770 510.340 1863.050 514.000 ;
        RECT 1862.700 510.000 1863.050 510.340 ;
        RECT 1862.700 503.610 1862.840 510.000 ;
        RECT 1862.700 503.470 1863.300 503.610 ;
        RECT 1863.160 486.870 1863.300 503.470 ;
        RECT 1863.100 486.550 1863.360 486.870 ;
        RECT 2021.800 486.210 2022.060 486.530 ;
        RECT 2021.860 62.210 2022.000 486.210 ;
        RECT 2021.800 61.890 2022.060 62.210 ;
        RECT 2024.560 61.890 2024.820 62.210 ;
        RECT 2024.620 2.400 2024.760 61.890 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 65.860 1876.730 65.920 ;
        RECT 2042.930 65.860 2043.250 65.920 ;
        RECT 1876.410 65.720 2043.250 65.860 ;
        RECT 1876.410 65.660 1876.730 65.720 ;
        RECT 2042.930 65.660 2043.250 65.720 ;
      LAYER via ;
        RECT 1876.440 65.660 1876.700 65.920 ;
        RECT 2042.960 65.660 2043.220 65.920 ;
      LAYER met2 ;
        RECT 1875.650 510.410 1875.930 514.000 ;
        RECT 1875.650 510.270 1876.640 510.410 ;
        RECT 1875.650 510.000 1875.930 510.270 ;
        RECT 1876.500 65.950 1876.640 510.270 ;
        RECT 1876.440 65.630 1876.700 65.950 ;
        RECT 2042.960 65.630 2043.220 65.950 ;
        RECT 2043.020 37.810 2043.160 65.630 ;
        RECT 2042.560 37.670 2043.160 37.810 ;
        RECT 2042.560 2.400 2042.700 37.670 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 757.765 2.805 757.935 48.195 ;
      LAYER mcon ;
        RECT 757.765 48.025 757.935 48.195 ;
      LAYER met1 ;
        RECT 758.150 86.260 758.470 86.320 ;
        RECT 952.270 86.260 952.590 86.320 ;
        RECT 758.150 86.120 952.590 86.260 ;
        RECT 758.150 86.060 758.470 86.120 ;
        RECT 952.270 86.060 952.590 86.120 ;
        RECT 757.705 48.180 757.995 48.225 ;
        RECT 758.150 48.180 758.470 48.240 ;
        RECT 757.705 48.040 758.470 48.180 ;
        RECT 757.705 47.995 757.995 48.040 ;
        RECT 758.150 47.980 758.470 48.040 ;
        RECT 757.690 2.960 758.010 3.020 ;
        RECT 757.495 2.820 758.010 2.960 ;
        RECT 757.690 2.760 758.010 2.820 ;
      LAYER via ;
        RECT 758.180 86.060 758.440 86.320 ;
        RECT 952.300 86.060 952.560 86.320 ;
        RECT 758.180 47.980 758.440 48.240 ;
        RECT 757.720 2.760 757.980 3.020 ;
      LAYER met2 ;
        RECT 953.810 510.410 954.090 514.000 ;
        RECT 952.360 510.270 954.090 510.410 ;
        RECT 952.360 86.350 952.500 510.270 ;
        RECT 953.810 510.000 954.090 510.270 ;
        RECT 758.180 86.030 758.440 86.350 ;
        RECT 952.300 86.030 952.560 86.350 ;
        RECT 758.240 48.270 758.380 86.030 ;
        RECT 758.180 47.950 758.440 48.270 ;
        RECT 757.720 2.730 757.980 3.050 ;
        RECT 757.780 2.400 757.920 2.730 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1888.370 500.040 1888.690 500.100 ;
        RECT 2056.730 500.040 2057.050 500.100 ;
        RECT 1888.370 499.900 2057.050 500.040 ;
        RECT 1888.370 499.840 1888.690 499.900 ;
        RECT 2056.730 499.840 2057.050 499.900 ;
        RECT 2056.730 62.120 2057.050 62.180 ;
        RECT 2060.410 62.120 2060.730 62.180 ;
        RECT 2056.730 61.980 2060.730 62.120 ;
        RECT 2056.730 61.920 2057.050 61.980 ;
        RECT 2060.410 61.920 2060.730 61.980 ;
      LAYER via ;
        RECT 1888.400 499.840 1888.660 500.100 ;
        RECT 2056.760 499.840 2057.020 500.100 ;
        RECT 2056.760 61.920 2057.020 62.180 ;
        RECT 2060.440 61.920 2060.700 62.180 ;
      LAYER met2 ;
        RECT 1888.530 510.340 1888.810 514.000 ;
        RECT 1888.460 510.000 1888.810 510.340 ;
        RECT 1888.460 500.130 1888.600 510.000 ;
        RECT 1888.400 499.810 1888.660 500.130 ;
        RECT 2056.760 499.810 2057.020 500.130 ;
        RECT 2056.820 62.210 2056.960 499.810 ;
        RECT 2056.760 61.890 2057.020 62.210 ;
        RECT 2060.440 61.890 2060.700 62.210 ;
        RECT 2060.500 2.400 2060.640 61.890 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 37.980 1904.330 38.040 ;
        RECT 2078.350 37.980 2078.670 38.040 ;
        RECT 1904.010 37.840 2078.670 37.980 ;
        RECT 1904.010 37.780 1904.330 37.840 ;
        RECT 2078.350 37.780 2078.670 37.840 ;
      LAYER via ;
        RECT 1904.040 37.780 1904.300 38.040 ;
        RECT 2078.380 37.780 2078.640 38.040 ;
      LAYER met2 ;
        RECT 1901.410 510.410 1901.690 514.000 ;
        RECT 1901.410 510.270 1904.240 510.410 ;
        RECT 1901.410 510.000 1901.690 510.270 ;
        RECT 1904.100 38.070 1904.240 510.270 ;
        RECT 1904.040 37.750 1904.300 38.070 ;
        RECT 2078.380 37.750 2078.640 38.070 ;
        RECT 2078.440 2.400 2078.580 37.750 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 30.840 1918.130 30.900 ;
        RECT 2095.830 30.840 2096.150 30.900 ;
        RECT 1917.810 30.700 2096.150 30.840 ;
        RECT 1917.810 30.640 1918.130 30.700 ;
        RECT 2095.830 30.640 2096.150 30.700 ;
      LAYER via ;
        RECT 1917.840 30.640 1918.100 30.900 ;
        RECT 2095.860 30.640 2096.120 30.900 ;
      LAYER met2 ;
        RECT 1914.290 510.410 1914.570 514.000 ;
        RECT 1914.290 510.270 1918.040 510.410 ;
        RECT 1914.290 510.000 1914.570 510.270 ;
        RECT 1917.900 30.930 1918.040 510.270 ;
        RECT 1917.840 30.610 1918.100 30.930 ;
        RECT 2095.860 30.610 2096.120 30.930 ;
        RECT 2095.920 2.400 2096.060 30.610 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2111.545 48.365 2111.715 137.955 ;
      LAYER mcon ;
        RECT 2111.545 137.785 2111.715 137.955 ;
      LAYER met1 ;
        RECT 1926.550 479.640 1926.870 479.700 ;
        RECT 2111.470 479.640 2111.790 479.700 ;
        RECT 1926.550 479.500 2111.790 479.640 ;
        RECT 1926.550 479.440 1926.870 479.500 ;
        RECT 2111.470 479.440 2111.790 479.500 ;
        RECT 2111.470 289.580 2111.790 289.640 ;
        RECT 2111.930 289.580 2112.250 289.640 ;
        RECT 2111.470 289.440 2112.250 289.580 ;
        RECT 2111.470 289.380 2111.790 289.440 ;
        RECT 2111.930 289.380 2112.250 289.440 ;
        RECT 2111.470 193.020 2111.790 193.080 ;
        RECT 2111.930 193.020 2112.250 193.080 ;
        RECT 2111.470 192.880 2112.250 193.020 ;
        RECT 2111.470 192.820 2111.790 192.880 ;
        RECT 2111.930 192.820 2112.250 192.880 ;
        RECT 2111.470 137.940 2111.790 138.000 ;
        RECT 2111.275 137.800 2111.790 137.940 ;
        RECT 2111.470 137.740 2111.790 137.800 ;
        RECT 2111.485 48.520 2111.775 48.565 ;
        RECT 2113.770 48.520 2114.090 48.580 ;
        RECT 2111.485 48.380 2114.090 48.520 ;
        RECT 2111.485 48.335 2111.775 48.380 ;
        RECT 2113.770 48.320 2114.090 48.380 ;
      LAYER via ;
        RECT 1926.580 479.440 1926.840 479.700 ;
        RECT 2111.500 479.440 2111.760 479.700 ;
        RECT 2111.500 289.380 2111.760 289.640 ;
        RECT 2111.960 289.380 2112.220 289.640 ;
        RECT 2111.500 192.820 2111.760 193.080 ;
        RECT 2111.960 192.820 2112.220 193.080 ;
        RECT 2111.500 137.740 2111.760 138.000 ;
        RECT 2113.800 48.320 2114.060 48.580 ;
      LAYER met2 ;
        RECT 1926.710 510.340 1926.990 514.000 ;
        RECT 1926.640 510.000 1926.990 510.340 ;
        RECT 1926.640 479.730 1926.780 510.000 ;
        RECT 1926.580 479.410 1926.840 479.730 ;
        RECT 2111.500 479.410 2111.760 479.730 ;
        RECT 2111.560 289.670 2111.700 479.410 ;
        RECT 2111.500 289.350 2111.760 289.670 ;
        RECT 2111.960 289.350 2112.220 289.670 ;
        RECT 2112.020 241.810 2112.160 289.350 ;
        RECT 2111.560 241.670 2112.160 241.810 ;
        RECT 2111.560 193.110 2111.700 241.670 ;
        RECT 2111.500 192.790 2111.760 193.110 ;
        RECT 2111.960 192.790 2112.220 193.110 ;
        RECT 2112.020 145.250 2112.160 192.790 ;
        RECT 2111.560 145.110 2112.160 145.250 ;
        RECT 2111.560 138.030 2111.700 145.110 ;
        RECT 2111.500 137.710 2111.760 138.030 ;
        RECT 2113.800 48.290 2114.060 48.610 ;
        RECT 2113.860 2.400 2114.000 48.290 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1939.430 503.100 1939.750 503.160 ;
        RECT 1945.410 503.100 1945.730 503.160 ;
        RECT 1939.430 502.960 1945.730 503.100 ;
        RECT 1939.430 502.900 1939.750 502.960 ;
        RECT 1945.410 502.900 1945.730 502.960 ;
        RECT 1945.410 44.780 1945.730 44.840 ;
        RECT 2131.710 44.780 2132.030 44.840 ;
        RECT 1945.410 44.640 2132.030 44.780 ;
        RECT 1945.410 44.580 1945.730 44.640 ;
        RECT 2131.710 44.580 2132.030 44.640 ;
      LAYER via ;
        RECT 1939.460 502.900 1939.720 503.160 ;
        RECT 1945.440 502.900 1945.700 503.160 ;
        RECT 1945.440 44.580 1945.700 44.840 ;
        RECT 2131.740 44.580 2132.000 44.840 ;
      LAYER met2 ;
        RECT 1939.590 510.340 1939.870 514.000 ;
        RECT 1939.520 510.000 1939.870 510.340 ;
        RECT 1939.520 503.190 1939.660 510.000 ;
        RECT 1939.460 502.870 1939.720 503.190 ;
        RECT 1945.440 502.870 1945.700 503.190 ;
        RECT 1945.500 44.870 1945.640 502.870 ;
        RECT 1945.440 44.550 1945.700 44.870 ;
        RECT 2131.740 44.550 2132.000 44.870 ;
        RECT 2131.800 2.400 2131.940 44.550 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 496.980 1952.630 497.040 ;
        RECT 1955.990 496.980 1956.310 497.040 ;
        RECT 1952.310 496.840 1956.310 496.980 ;
        RECT 1952.310 496.780 1952.630 496.840 ;
        RECT 1955.990 496.780 1956.310 496.840 ;
        RECT 1955.990 272.580 1956.310 272.640 ;
        RECT 2145.970 272.580 2146.290 272.640 ;
        RECT 1955.990 272.440 2146.290 272.580 ;
        RECT 1955.990 272.380 1956.310 272.440 ;
        RECT 2145.970 272.380 2146.290 272.440 ;
        RECT 2145.970 62.120 2146.290 62.180 ;
        RECT 2149.650 62.120 2149.970 62.180 ;
        RECT 2145.970 61.980 2149.970 62.120 ;
        RECT 2145.970 61.920 2146.290 61.980 ;
        RECT 2149.650 61.920 2149.970 61.980 ;
      LAYER via ;
        RECT 1952.340 496.780 1952.600 497.040 ;
        RECT 1956.020 496.780 1956.280 497.040 ;
        RECT 1956.020 272.380 1956.280 272.640 ;
        RECT 2146.000 272.380 2146.260 272.640 ;
        RECT 2146.000 61.920 2146.260 62.180 ;
        RECT 2149.680 61.920 2149.940 62.180 ;
      LAYER met2 ;
        RECT 1952.470 510.340 1952.750 514.000 ;
        RECT 1952.400 510.000 1952.750 510.340 ;
        RECT 1952.400 497.070 1952.540 510.000 ;
        RECT 1952.340 496.750 1952.600 497.070 ;
        RECT 1956.020 496.750 1956.280 497.070 ;
        RECT 1956.080 272.670 1956.220 496.750 ;
        RECT 1956.020 272.350 1956.280 272.670 ;
        RECT 2146.000 272.350 2146.260 272.670 ;
        RECT 2146.060 62.210 2146.200 272.350 ;
        RECT 2146.000 61.890 2146.260 62.210 ;
        RECT 2149.680 61.890 2149.940 62.210 ;
        RECT 2149.740 2.400 2149.880 61.890 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 51.580 1966.430 51.640 ;
        RECT 2167.590 51.580 2167.910 51.640 ;
        RECT 1966.110 51.440 2167.910 51.580 ;
        RECT 1966.110 51.380 1966.430 51.440 ;
        RECT 2167.590 51.380 2167.910 51.440 ;
      LAYER via ;
        RECT 1966.140 51.380 1966.400 51.640 ;
        RECT 2167.620 51.380 2167.880 51.640 ;
      LAYER met2 ;
        RECT 1965.350 510.410 1965.630 514.000 ;
        RECT 1965.350 510.270 1966.340 510.410 ;
        RECT 1965.350 510.000 1965.630 510.270 ;
        RECT 1966.200 51.670 1966.340 510.270 ;
        RECT 1966.140 51.350 1966.400 51.670 ;
        RECT 2167.620 51.350 2167.880 51.670 ;
        RECT 2167.680 2.400 2167.820 51.350 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 58.720 1980.230 58.780 ;
        RECT 2185.070 58.720 2185.390 58.780 ;
        RECT 1979.910 58.580 2185.390 58.720 ;
        RECT 1979.910 58.520 1980.230 58.580 ;
        RECT 2185.070 58.520 2185.390 58.580 ;
      LAYER via ;
        RECT 1979.940 58.520 1980.200 58.780 ;
        RECT 2185.100 58.520 2185.360 58.780 ;
      LAYER met2 ;
        RECT 1978.230 510.410 1978.510 514.000 ;
        RECT 1978.230 510.270 1980.140 510.410 ;
        RECT 1978.230 510.000 1978.510 510.270 ;
        RECT 1980.000 58.810 1980.140 510.270 ;
        RECT 1979.940 58.490 1980.200 58.810 ;
        RECT 2185.100 58.490 2185.360 58.810 ;
        RECT 2185.160 2.400 2185.300 58.490 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 72.320 1994.030 72.380 ;
        RECT 2201.170 72.320 2201.490 72.380 ;
        RECT 1993.710 72.180 2201.490 72.320 ;
        RECT 1993.710 72.120 1994.030 72.180 ;
        RECT 2201.170 72.120 2201.490 72.180 ;
      LAYER via ;
        RECT 1993.740 72.120 1994.000 72.380 ;
        RECT 2201.200 72.120 2201.460 72.380 ;
      LAYER met2 ;
        RECT 1991.110 510.410 1991.390 514.000 ;
        RECT 1991.110 510.270 1993.940 510.410 ;
        RECT 1991.110 510.000 1991.390 510.270 ;
        RECT 1993.800 72.410 1993.940 510.270 ;
        RECT 1993.740 72.090 1994.000 72.410 ;
        RECT 2201.200 72.090 2201.460 72.410 ;
        RECT 2201.260 17.410 2201.400 72.090 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2003.370 496.980 2003.690 497.040 ;
        RECT 2007.510 496.980 2007.830 497.040 ;
        RECT 2003.370 496.840 2007.830 496.980 ;
        RECT 2003.370 496.780 2003.690 496.840 ;
        RECT 2007.510 496.780 2007.830 496.840 ;
        RECT 2007.510 79.460 2007.830 79.520 ;
        RECT 2215.430 79.460 2215.750 79.520 ;
        RECT 2007.510 79.320 2215.750 79.460 ;
        RECT 2007.510 79.260 2007.830 79.320 ;
        RECT 2215.430 79.260 2215.750 79.320 ;
      LAYER via ;
        RECT 2003.400 496.780 2003.660 497.040 ;
        RECT 2007.540 496.780 2007.800 497.040 ;
        RECT 2007.540 79.260 2007.800 79.520 ;
        RECT 2215.460 79.260 2215.720 79.520 ;
      LAYER met2 ;
        RECT 2003.530 510.340 2003.810 514.000 ;
        RECT 2003.460 510.000 2003.810 510.340 ;
        RECT 2003.460 497.070 2003.600 510.000 ;
        RECT 2003.400 496.750 2003.660 497.070 ;
        RECT 2007.540 496.750 2007.800 497.070 ;
        RECT 2007.600 79.550 2007.740 496.750 ;
        RECT 2007.540 79.230 2007.800 79.550 ;
        RECT 2215.460 79.230 2215.720 79.550 ;
        RECT 2215.520 17.410 2215.660 79.230 ;
        RECT 2215.520 17.270 2221.180 17.410 ;
        RECT 2221.040 2.400 2221.180 17.270 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 93.060 779.630 93.120 ;
        RECT 966.070 93.060 966.390 93.120 ;
        RECT 779.310 92.920 966.390 93.060 ;
        RECT 779.310 92.860 779.630 92.920 ;
        RECT 966.070 92.860 966.390 92.920 ;
        RECT 775.630 15.880 775.950 15.940 ;
        RECT 779.310 15.880 779.630 15.940 ;
        RECT 775.630 15.740 779.630 15.880 ;
        RECT 775.630 15.680 775.950 15.740 ;
        RECT 779.310 15.680 779.630 15.740 ;
      LAYER via ;
        RECT 779.340 92.860 779.600 93.120 ;
        RECT 966.100 92.860 966.360 93.120 ;
        RECT 775.660 15.680 775.920 15.940 ;
        RECT 779.340 15.680 779.600 15.940 ;
      LAYER met2 ;
        RECT 966.690 510.410 966.970 514.000 ;
        RECT 966.160 510.270 966.970 510.410 ;
        RECT 966.160 93.150 966.300 510.270 ;
        RECT 966.690 510.000 966.970 510.270 ;
        RECT 779.340 92.830 779.600 93.150 ;
        RECT 966.100 92.830 966.360 93.150 ;
        RECT 779.400 15.970 779.540 92.830 ;
        RECT 775.660 15.650 775.920 15.970 ;
        RECT 779.340 15.650 779.600 15.970 ;
        RECT 775.720 2.400 775.860 15.650 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.250 496.980 2016.570 497.040 ;
        RECT 2020.850 496.980 2021.170 497.040 ;
        RECT 2016.250 496.840 2021.170 496.980 ;
        RECT 2016.250 496.780 2016.570 496.840 ;
        RECT 2020.850 496.780 2021.170 496.840 ;
        RECT 2020.850 86.260 2021.170 86.320 ;
        RECT 2235.670 86.260 2235.990 86.320 ;
        RECT 2020.850 86.120 2235.990 86.260 ;
        RECT 2020.850 86.060 2021.170 86.120 ;
        RECT 2235.670 86.060 2235.990 86.120 ;
      LAYER via ;
        RECT 2016.280 496.780 2016.540 497.040 ;
        RECT 2020.880 496.780 2021.140 497.040 ;
        RECT 2020.880 86.060 2021.140 86.320 ;
        RECT 2235.700 86.060 2235.960 86.320 ;
      LAYER met2 ;
        RECT 2016.410 510.340 2016.690 514.000 ;
        RECT 2016.340 510.000 2016.690 510.340 ;
        RECT 2016.340 497.070 2016.480 510.000 ;
        RECT 2016.280 496.750 2016.540 497.070 ;
        RECT 2020.880 496.750 2021.140 497.070 ;
        RECT 2020.940 86.350 2021.080 496.750 ;
        RECT 2020.880 86.030 2021.140 86.350 ;
        RECT 2235.700 86.030 2235.960 86.350 ;
        RECT 2235.760 17.410 2235.900 86.030 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2029.130 496.980 2029.450 497.040 ;
        RECT 2035.110 496.980 2035.430 497.040 ;
        RECT 2029.130 496.840 2035.430 496.980 ;
        RECT 2029.130 496.780 2029.450 496.840 ;
        RECT 2035.110 496.780 2035.430 496.840 ;
        RECT 2035.110 93.060 2035.430 93.120 ;
        RECT 2256.830 93.060 2257.150 93.120 ;
        RECT 2035.110 92.920 2257.150 93.060 ;
        RECT 2035.110 92.860 2035.430 92.920 ;
        RECT 2256.830 92.860 2257.150 92.920 ;
      LAYER via ;
        RECT 2029.160 496.780 2029.420 497.040 ;
        RECT 2035.140 496.780 2035.400 497.040 ;
        RECT 2035.140 92.860 2035.400 93.120 ;
        RECT 2256.860 92.860 2257.120 93.120 ;
      LAYER met2 ;
        RECT 2029.290 510.340 2029.570 514.000 ;
        RECT 2029.220 510.000 2029.570 510.340 ;
        RECT 2029.220 497.070 2029.360 510.000 ;
        RECT 2029.160 496.750 2029.420 497.070 ;
        RECT 2035.140 496.750 2035.400 497.070 ;
        RECT 2035.200 93.150 2035.340 496.750 ;
        RECT 2035.140 92.830 2035.400 93.150 ;
        RECT 2256.860 92.830 2257.120 93.150 ;
        RECT 2256.920 7.210 2257.060 92.830 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 496.980 2042.330 497.040 ;
        RECT 2045.690 496.980 2046.010 497.040 ;
        RECT 2042.010 496.840 2046.010 496.980 ;
        RECT 2042.010 496.780 2042.330 496.840 ;
        RECT 2045.690 496.780 2046.010 496.840 ;
        RECT 2045.690 99.860 2046.010 99.920 ;
        RECT 2270.170 99.860 2270.490 99.920 ;
        RECT 2045.690 99.720 2270.490 99.860 ;
        RECT 2045.690 99.660 2046.010 99.720 ;
        RECT 2270.170 99.660 2270.490 99.720 ;
      LAYER via ;
        RECT 2042.040 496.780 2042.300 497.040 ;
        RECT 2045.720 496.780 2045.980 497.040 ;
        RECT 2045.720 99.660 2045.980 99.920 ;
        RECT 2270.200 99.660 2270.460 99.920 ;
      LAYER met2 ;
        RECT 2042.170 510.340 2042.450 514.000 ;
        RECT 2042.100 510.000 2042.450 510.340 ;
        RECT 2042.100 497.070 2042.240 510.000 ;
        RECT 2042.040 496.750 2042.300 497.070 ;
        RECT 2045.720 496.750 2045.980 497.070 ;
        RECT 2045.780 99.950 2045.920 496.750 ;
        RECT 2045.720 99.630 2045.980 99.950 ;
        RECT 2270.200 99.630 2270.460 99.950 ;
        RECT 2270.260 17.410 2270.400 99.630 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2054.505 349.945 2054.675 372.555 ;
      LAYER mcon ;
        RECT 2054.505 372.385 2054.675 372.555 ;
      LAYER met1 ;
        RECT 2054.430 476.240 2054.750 476.300 ;
        RECT 2055.350 476.240 2055.670 476.300 ;
        RECT 2054.430 476.100 2055.670 476.240 ;
        RECT 2054.430 476.040 2054.750 476.100 ;
        RECT 2055.350 476.040 2055.670 476.100 ;
        RECT 2054.430 372.540 2054.750 372.600 ;
        RECT 2054.235 372.400 2054.750 372.540 ;
        RECT 2054.430 372.340 2054.750 372.400 ;
        RECT 2054.445 350.100 2054.735 350.145 ;
        RECT 2054.890 350.100 2055.210 350.160 ;
        RECT 2054.445 349.960 2055.210 350.100 ;
        RECT 2054.445 349.915 2054.735 349.960 ;
        RECT 2054.890 349.900 2055.210 349.960 ;
        RECT 2054.890 317.460 2055.210 317.520 ;
        RECT 2055.350 317.460 2055.670 317.520 ;
        RECT 2054.890 317.320 2055.670 317.460 ;
        RECT 2054.890 317.260 2055.210 317.320 ;
        RECT 2055.350 317.260 2055.670 317.320 ;
        RECT 2054.890 227.500 2055.210 227.760 ;
        RECT 2054.980 227.080 2055.120 227.500 ;
        RECT 2054.890 226.820 2055.210 227.080 ;
        RECT 2054.890 107.000 2055.210 107.060 ;
        RECT 2290.870 107.000 2291.190 107.060 ;
        RECT 2054.890 106.860 2291.190 107.000 ;
        RECT 2054.890 106.800 2055.210 106.860 ;
        RECT 2290.870 106.800 2291.190 106.860 ;
      LAYER via ;
        RECT 2054.460 476.040 2054.720 476.300 ;
        RECT 2055.380 476.040 2055.640 476.300 ;
        RECT 2054.460 372.340 2054.720 372.600 ;
        RECT 2054.920 349.900 2055.180 350.160 ;
        RECT 2054.920 317.260 2055.180 317.520 ;
        RECT 2055.380 317.260 2055.640 317.520 ;
        RECT 2054.920 227.500 2055.180 227.760 ;
        RECT 2054.920 226.820 2055.180 227.080 ;
        RECT 2054.920 106.800 2055.180 107.060 ;
        RECT 2290.900 106.800 2291.160 107.060 ;
      LAYER met2 ;
        RECT 2055.050 510.410 2055.330 514.000 ;
        RECT 2054.520 510.270 2055.330 510.410 ;
        RECT 2054.520 476.330 2054.660 510.270 ;
        RECT 2055.050 510.000 2055.330 510.270 ;
        RECT 2054.460 476.010 2054.720 476.330 ;
        RECT 2055.380 476.010 2055.640 476.330 ;
        RECT 2055.440 435.725 2055.580 476.010 ;
        RECT 2055.370 435.355 2055.650 435.725 ;
        RECT 2054.910 434.675 2055.190 435.045 ;
        RECT 2054.980 399.570 2055.120 434.675 ;
        RECT 2054.520 399.430 2055.120 399.570 ;
        RECT 2054.520 372.630 2054.660 399.430 ;
        RECT 2054.460 372.310 2054.720 372.630 ;
        RECT 2054.920 349.870 2055.180 350.190 ;
        RECT 2054.980 317.550 2055.120 349.870 ;
        RECT 2054.920 317.230 2055.180 317.550 ;
        RECT 2055.380 317.230 2055.640 317.550 ;
        RECT 2055.440 234.330 2055.580 317.230 ;
        RECT 2054.980 234.190 2055.580 234.330 ;
        RECT 2054.980 227.790 2055.120 234.190 ;
        RECT 2054.920 227.470 2055.180 227.790 ;
        RECT 2054.920 226.790 2055.180 227.110 ;
        RECT 2054.980 107.090 2055.120 226.790 ;
        RECT 2054.920 106.770 2055.180 107.090 ;
        RECT 2290.900 106.770 2291.160 107.090 ;
        RECT 2290.960 17.410 2291.100 106.770 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
      LAYER via2 ;
        RECT 2055.370 435.400 2055.650 435.680 ;
        RECT 2054.910 434.720 2055.190 435.000 ;
      LAYER met3 ;
        RECT 2055.345 435.690 2055.675 435.705 ;
        RECT 2054.670 435.390 2055.675 435.690 ;
        RECT 2054.670 435.025 2054.970 435.390 ;
        RECT 2055.345 435.375 2055.675 435.390 ;
        RECT 2054.670 434.710 2055.215 435.025 ;
        RECT 2054.885 434.695 2055.215 434.710 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2067.770 497.320 2068.090 497.380 ;
        RECT 2080.190 497.320 2080.510 497.380 ;
        RECT 2067.770 497.180 2080.510 497.320 ;
        RECT 2067.770 497.120 2068.090 497.180 ;
        RECT 2080.190 497.120 2080.510 497.180 ;
        RECT 2080.190 113.800 2080.510 113.860 ;
        RECT 2304.670 113.800 2304.990 113.860 ;
        RECT 2080.190 113.660 2304.990 113.800 ;
        RECT 2080.190 113.600 2080.510 113.660 ;
        RECT 2304.670 113.600 2304.990 113.660 ;
      LAYER via ;
        RECT 2067.800 497.120 2068.060 497.380 ;
        RECT 2080.220 497.120 2080.480 497.380 ;
        RECT 2080.220 113.600 2080.480 113.860 ;
        RECT 2304.700 113.600 2304.960 113.860 ;
      LAYER met2 ;
        RECT 2067.930 510.340 2068.210 514.000 ;
        RECT 2067.860 510.000 2068.210 510.340 ;
        RECT 2067.860 497.410 2068.000 510.000 ;
        RECT 2067.800 497.090 2068.060 497.410 ;
        RECT 2080.220 497.090 2080.480 497.410 ;
        RECT 2080.280 113.890 2080.420 497.090 ;
        RECT 2080.220 113.570 2080.480 113.890 ;
        RECT 2304.700 113.570 2304.960 113.890 ;
        RECT 2304.760 17.410 2304.900 113.570 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 120.600 2083.730 120.660 ;
        RECT 2325.370 120.600 2325.690 120.660 ;
        RECT 2083.410 120.460 2325.690 120.600 ;
        RECT 2083.410 120.400 2083.730 120.460 ;
        RECT 2325.370 120.400 2325.690 120.460 ;
      LAYER via ;
        RECT 2083.440 120.400 2083.700 120.660 ;
        RECT 2325.400 120.400 2325.660 120.660 ;
      LAYER met2 ;
        RECT 2080.350 510.410 2080.630 514.000 ;
        RECT 2080.350 510.270 2083.640 510.410 ;
        RECT 2080.350 510.000 2080.630 510.270 ;
        RECT 2083.500 120.690 2083.640 510.270 ;
        RECT 2083.440 120.370 2083.700 120.690 ;
        RECT 2325.400 120.370 2325.660 120.690 ;
        RECT 2325.460 17.410 2325.600 120.370 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2093.070 499.020 2093.390 499.080 ;
        RECT 2100.890 499.020 2101.210 499.080 ;
        RECT 2093.070 498.880 2101.210 499.020 ;
        RECT 2093.070 498.820 2093.390 498.880 ;
        RECT 2100.890 498.820 2101.210 498.880 ;
        RECT 2100.890 127.740 2101.210 127.800 ;
        RECT 2339.630 127.740 2339.950 127.800 ;
        RECT 2100.890 127.600 2339.950 127.740 ;
        RECT 2100.890 127.540 2101.210 127.600 ;
        RECT 2339.630 127.540 2339.950 127.600 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.610 16.900 2345.930 16.960 ;
        RECT 2339.630 16.760 2345.930 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.610 16.700 2345.930 16.760 ;
      LAYER via ;
        RECT 2093.100 498.820 2093.360 499.080 ;
        RECT 2100.920 498.820 2101.180 499.080 ;
        RECT 2100.920 127.540 2101.180 127.800 ;
        RECT 2339.660 127.540 2339.920 127.800 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.640 16.700 2345.900 16.960 ;
      LAYER met2 ;
        RECT 2093.230 510.340 2093.510 514.000 ;
        RECT 2093.160 510.000 2093.510 510.340 ;
        RECT 2093.160 499.110 2093.300 510.000 ;
        RECT 2093.100 498.790 2093.360 499.110 ;
        RECT 2100.920 498.790 2101.180 499.110 ;
        RECT 2100.980 127.830 2101.120 498.790 ;
        RECT 2100.920 127.510 2101.180 127.830 ;
        RECT 2339.660 127.510 2339.920 127.830 ;
        RECT 2339.720 16.990 2339.860 127.510 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.640 16.670 2345.900 16.990 ;
        RECT 2345.700 2.400 2345.840 16.670 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.950 503.440 2106.270 503.500 ;
        RECT 2111.010 503.440 2111.330 503.500 ;
        RECT 2105.950 503.300 2111.330 503.440 ;
        RECT 2105.950 503.240 2106.270 503.300 ;
        RECT 2111.010 503.240 2111.330 503.300 ;
        RECT 2111.010 134.540 2111.330 134.600 ;
        RECT 2359.870 134.540 2360.190 134.600 ;
        RECT 2111.010 134.400 2360.190 134.540 ;
        RECT 2111.010 134.340 2111.330 134.400 ;
        RECT 2359.870 134.340 2360.190 134.400 ;
      LAYER via ;
        RECT 2105.980 503.240 2106.240 503.500 ;
        RECT 2111.040 503.240 2111.300 503.500 ;
        RECT 2111.040 134.340 2111.300 134.600 ;
        RECT 2359.900 134.340 2360.160 134.600 ;
      LAYER met2 ;
        RECT 2106.110 510.340 2106.390 514.000 ;
        RECT 2106.040 510.000 2106.390 510.340 ;
        RECT 2106.040 503.530 2106.180 510.000 ;
        RECT 2105.980 503.210 2106.240 503.530 ;
        RECT 2111.040 503.210 2111.300 503.530 ;
        RECT 2111.100 134.630 2111.240 503.210 ;
        RECT 2111.040 134.310 2111.300 134.630 ;
        RECT 2359.900 134.310 2360.160 134.630 ;
        RECT 2359.960 16.730 2360.100 134.310 ;
        RECT 2359.960 16.590 2363.780 16.730 ;
        RECT 2363.640 2.400 2363.780 16.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2118.830 503.100 2119.150 503.160 ;
        RECT 2124.810 503.100 2125.130 503.160 ;
        RECT 2118.830 502.960 2125.130 503.100 ;
        RECT 2118.830 502.900 2119.150 502.960 ;
        RECT 2124.810 502.900 2125.130 502.960 ;
        RECT 2124.810 141.680 2125.130 141.740 ;
        RECT 2380.570 141.680 2380.890 141.740 ;
        RECT 2124.810 141.540 2380.890 141.680 ;
        RECT 2124.810 141.480 2125.130 141.540 ;
        RECT 2380.570 141.480 2380.890 141.540 ;
      LAYER via ;
        RECT 2118.860 502.900 2119.120 503.160 ;
        RECT 2124.840 502.900 2125.100 503.160 ;
        RECT 2124.840 141.480 2125.100 141.740 ;
        RECT 2380.600 141.480 2380.860 141.740 ;
      LAYER met2 ;
        RECT 2118.990 510.340 2119.270 514.000 ;
        RECT 2118.920 510.000 2119.270 510.340 ;
        RECT 2118.920 503.190 2119.060 510.000 ;
        RECT 2118.860 502.870 2119.120 503.190 ;
        RECT 2124.840 502.870 2125.100 503.190 ;
        RECT 2124.900 141.770 2125.040 502.870 ;
        RECT 2124.840 141.450 2125.100 141.770 ;
        RECT 2380.600 141.450 2380.860 141.770 ;
        RECT 2380.660 16.730 2380.800 141.450 ;
        RECT 2380.660 16.590 2381.720 16.730 ;
        RECT 2381.580 2.400 2381.720 16.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 503.440 2132.030 503.500 ;
        RECT 2135.390 503.440 2135.710 503.500 ;
        RECT 2131.710 503.300 2135.710 503.440 ;
        RECT 2131.710 503.240 2132.030 503.300 ;
        RECT 2135.390 503.240 2135.710 503.300 ;
        RECT 2135.390 155.280 2135.710 155.340 ;
        RECT 2394.370 155.280 2394.690 155.340 ;
        RECT 2135.390 155.140 2394.690 155.280 ;
        RECT 2135.390 155.080 2135.710 155.140 ;
        RECT 2394.370 155.080 2394.690 155.140 ;
      LAYER via ;
        RECT 2131.740 503.240 2132.000 503.500 ;
        RECT 2135.420 503.240 2135.680 503.500 ;
        RECT 2135.420 155.080 2135.680 155.340 ;
        RECT 2394.400 155.080 2394.660 155.340 ;
      LAYER met2 ;
        RECT 2131.870 510.340 2132.150 514.000 ;
        RECT 2131.800 510.000 2132.150 510.340 ;
        RECT 2131.800 503.530 2131.940 510.000 ;
        RECT 2131.740 503.210 2132.000 503.530 ;
        RECT 2135.420 503.210 2135.680 503.530 ;
        RECT 2135.480 155.370 2135.620 503.210 ;
        RECT 2135.420 155.050 2135.680 155.370 ;
        RECT 2394.400 155.050 2394.660 155.370 ;
        RECT 2394.460 16.730 2394.600 155.050 ;
        RECT 2394.460 16.590 2399.660 16.730 ;
        RECT 2399.520 2.400 2399.660 16.590 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.970 489.840 973.290 489.900 ;
        RECT 978.030 489.840 978.350 489.900 ;
        RECT 972.970 489.700 978.350 489.840 ;
        RECT 972.970 489.640 973.290 489.700 ;
        RECT 978.030 489.640 978.350 489.700 ;
        RECT 799.550 99.860 799.870 99.920 ;
        RECT 972.970 99.860 973.290 99.920 ;
        RECT 799.550 99.720 973.290 99.860 ;
        RECT 799.550 99.660 799.870 99.720 ;
        RECT 972.970 99.660 973.290 99.720 ;
        RECT 793.570 20.640 793.890 20.700 ;
        RECT 799.550 20.640 799.870 20.700 ;
        RECT 793.570 20.500 799.870 20.640 ;
        RECT 793.570 20.440 793.890 20.500 ;
        RECT 799.550 20.440 799.870 20.500 ;
      LAYER via ;
        RECT 973.000 489.640 973.260 489.900 ;
        RECT 978.060 489.640 978.320 489.900 ;
        RECT 799.580 99.660 799.840 99.920 ;
        RECT 973.000 99.660 973.260 99.920 ;
        RECT 793.600 20.440 793.860 20.700 ;
        RECT 799.580 20.440 799.840 20.700 ;
      LAYER met2 ;
        RECT 979.570 510.410 979.850 514.000 ;
        RECT 978.120 510.270 979.850 510.410 ;
        RECT 978.120 489.930 978.260 510.270 ;
        RECT 979.570 510.000 979.850 510.270 ;
        RECT 973.000 489.610 973.260 489.930 ;
        RECT 978.060 489.610 978.320 489.930 ;
        RECT 973.060 99.950 973.200 489.610 ;
        RECT 799.580 99.630 799.840 99.950 ;
        RECT 973.000 99.630 973.260 99.950 ;
        RECT 799.640 20.730 799.780 99.630 ;
        RECT 793.600 20.410 793.860 20.730 ;
        RECT 799.580 20.410 799.840 20.730 ;
        RECT 793.660 2.400 793.800 20.410 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 864.485 448.205 864.655 483.055 ;
        RECT 863.105 379.525 863.275 403.835 ;
        RECT 864.485 234.685 864.655 289.595 ;
      LAYER mcon ;
        RECT 864.485 482.885 864.655 483.055 ;
        RECT 863.105 403.665 863.275 403.835 ;
        RECT 864.485 289.425 864.655 289.595 ;
      LAYER met1 ;
        RECT 864.425 483.040 864.715 483.085 ;
        RECT 865.790 483.040 866.110 483.100 ;
        RECT 864.425 482.900 866.110 483.040 ;
        RECT 864.425 482.855 864.715 482.900 ;
        RECT 865.790 482.840 866.110 482.900 ;
        RECT 864.410 448.360 864.730 448.420 ;
        RECT 864.215 448.220 864.730 448.360 ;
        RECT 864.410 448.160 864.730 448.220 ;
        RECT 863.045 403.820 863.335 403.865 ;
        RECT 864.410 403.820 864.730 403.880 ;
        RECT 863.045 403.680 864.730 403.820 ;
        RECT 863.045 403.635 863.335 403.680 ;
        RECT 864.410 403.620 864.730 403.680 ;
        RECT 863.030 379.680 863.350 379.740 ;
        RECT 862.835 379.540 863.350 379.680 ;
        RECT 863.030 379.480 863.350 379.540 ;
        RECT 863.950 303.860 864.270 303.920 ;
        RECT 863.950 303.720 864.640 303.860 ;
        RECT 863.950 303.660 864.270 303.720 ;
        RECT 864.500 303.580 864.640 303.720 ;
        RECT 864.410 303.320 864.730 303.580 ;
        RECT 864.410 289.580 864.730 289.640 ;
        RECT 864.215 289.440 864.730 289.580 ;
        RECT 864.410 289.380 864.730 289.440 ;
        RECT 863.030 234.840 863.350 234.900 ;
        RECT 864.425 234.840 864.715 234.885 ;
        RECT 863.030 234.700 864.715 234.840 ;
        RECT 863.030 234.640 863.350 234.700 ;
        RECT 864.425 234.655 864.715 234.700 ;
        RECT 863.030 207.100 863.350 207.360 ;
        RECT 863.120 206.620 863.260 207.100 ;
        RECT 863.490 206.620 863.810 206.680 ;
        RECT 863.120 206.480 863.810 206.620 ;
        RECT 863.490 206.420 863.810 206.480 ;
        RECT 863.490 145.420 863.810 145.480 ;
        RECT 863.120 145.280 863.810 145.420 ;
        RECT 863.120 145.140 863.260 145.280 ;
        RECT 863.490 145.220 863.810 145.280 ;
        RECT 863.030 144.880 863.350 145.140 ;
        RECT 641.310 107.340 641.630 107.400 ;
        RECT 863.030 107.340 863.350 107.400 ;
        RECT 641.310 107.200 863.350 107.340 ;
        RECT 641.310 107.140 641.630 107.200 ;
        RECT 863.030 107.140 863.350 107.200 ;
        RECT 639.010 16.900 639.330 16.960 ;
        RECT 641.310 16.900 641.630 16.960 ;
        RECT 639.010 16.760 641.630 16.900 ;
        RECT 639.010 16.700 639.330 16.760 ;
        RECT 641.310 16.700 641.630 16.760 ;
      LAYER via ;
        RECT 865.820 482.840 866.080 483.100 ;
        RECT 864.440 448.160 864.700 448.420 ;
        RECT 864.440 403.620 864.700 403.880 ;
        RECT 863.060 379.480 863.320 379.740 ;
        RECT 863.980 303.660 864.240 303.920 ;
        RECT 864.440 303.320 864.700 303.580 ;
        RECT 864.440 289.380 864.700 289.640 ;
        RECT 863.060 234.640 863.320 234.900 ;
        RECT 863.060 207.100 863.320 207.360 ;
        RECT 863.520 206.420 863.780 206.680 ;
        RECT 863.520 145.220 863.780 145.480 ;
        RECT 863.060 144.880 863.320 145.140 ;
        RECT 641.340 107.140 641.600 107.400 ;
        RECT 863.060 107.140 863.320 107.400 ;
        RECT 639.040 16.700 639.300 16.960 ;
        RECT 641.340 16.700 641.600 16.960 ;
      LAYER met2 ;
        RECT 868.250 510.410 868.530 514.000 ;
        RECT 865.880 510.270 868.530 510.410 ;
        RECT 865.880 483.130 866.020 510.270 ;
        RECT 868.250 510.000 868.530 510.270 ;
        RECT 865.820 482.810 866.080 483.130 ;
        RECT 864.440 448.130 864.700 448.450 ;
        RECT 864.500 403.910 864.640 448.130 ;
        RECT 864.440 403.590 864.700 403.910 ;
        RECT 863.060 379.450 863.320 379.770 ;
        RECT 863.120 351.970 863.260 379.450 ;
        RECT 863.120 351.830 864.180 351.970 ;
        RECT 864.040 303.950 864.180 351.830 ;
        RECT 863.980 303.630 864.240 303.950 ;
        RECT 864.440 303.290 864.700 303.610 ;
        RECT 864.500 289.670 864.640 303.290 ;
        RECT 864.440 289.350 864.700 289.670 ;
        RECT 863.060 234.610 863.320 234.930 ;
        RECT 863.120 207.390 863.260 234.610 ;
        RECT 863.060 207.070 863.320 207.390 ;
        RECT 863.520 206.390 863.780 206.710 ;
        RECT 863.580 145.510 863.720 206.390 ;
        RECT 863.520 145.190 863.780 145.510 ;
        RECT 863.060 144.850 863.320 145.170 ;
        RECT 863.120 107.430 863.260 144.850 ;
        RECT 641.340 107.110 641.600 107.430 ;
        RECT 863.060 107.110 863.320 107.430 ;
        RECT 641.400 16.990 641.540 107.110 ;
        RECT 639.040 16.670 639.300 16.990 ;
        RECT 641.340 16.670 641.600 16.990 ;
        RECT 639.100 2.400 639.240 16.670 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2152.410 162.080 2152.730 162.140 ;
        RECT 2421.970 162.080 2422.290 162.140 ;
        RECT 2152.410 161.940 2422.290 162.080 ;
        RECT 2152.410 161.880 2152.730 161.940 ;
        RECT 2421.970 161.880 2422.290 161.940 ;
      LAYER via ;
        RECT 2152.440 161.880 2152.700 162.140 ;
        RECT 2422.000 161.880 2422.260 162.140 ;
      LAYER met2 ;
        RECT 2148.890 510.410 2149.170 514.000 ;
        RECT 2148.890 510.270 2152.640 510.410 ;
        RECT 2148.890 510.000 2149.170 510.270 ;
        RECT 2152.500 162.170 2152.640 510.270 ;
        RECT 2152.440 161.850 2152.700 162.170 ;
        RECT 2422.000 161.850 2422.260 162.170 ;
        RECT 2422.060 16.730 2422.200 161.850 ;
        RECT 2422.060 16.590 2423.120 16.730 ;
        RECT 2422.980 2.400 2423.120 16.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2161.610 503.440 2161.930 503.500 ;
        RECT 2169.890 503.440 2170.210 503.500 ;
        RECT 2161.610 503.300 2170.210 503.440 ;
        RECT 2161.610 503.240 2161.930 503.300 ;
        RECT 2169.890 503.240 2170.210 503.300 ;
        RECT 2169.890 237.900 2170.210 237.960 ;
        RECT 2435.770 237.900 2436.090 237.960 ;
        RECT 2169.890 237.760 2436.090 237.900 ;
        RECT 2169.890 237.700 2170.210 237.760 ;
        RECT 2435.770 237.700 2436.090 237.760 ;
      LAYER via ;
        RECT 2161.640 503.240 2161.900 503.500 ;
        RECT 2169.920 503.240 2170.180 503.500 ;
        RECT 2169.920 237.700 2170.180 237.960 ;
        RECT 2435.800 237.700 2436.060 237.960 ;
      LAYER met2 ;
        RECT 2161.770 510.340 2162.050 514.000 ;
        RECT 2161.700 510.000 2162.050 510.340 ;
        RECT 2161.700 503.530 2161.840 510.000 ;
        RECT 2161.640 503.210 2161.900 503.530 ;
        RECT 2169.920 503.210 2170.180 503.530 ;
        RECT 2169.980 237.990 2170.120 503.210 ;
        RECT 2169.920 237.670 2170.180 237.990 ;
        RECT 2435.800 237.670 2436.060 237.990 ;
        RECT 2435.860 16.730 2436.000 237.670 ;
        RECT 2435.860 16.590 2441.060 16.730 ;
        RECT 2440.920 2.400 2441.060 16.590 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2174.490 503.440 2174.810 503.500 ;
        RECT 2180.010 503.440 2180.330 503.500 ;
        RECT 2174.490 503.300 2180.330 503.440 ;
        RECT 2174.490 503.240 2174.810 503.300 ;
        RECT 2180.010 503.240 2180.330 503.300 ;
        RECT 2180.010 168.880 2180.330 168.940 ;
        RECT 2456.470 168.880 2456.790 168.940 ;
        RECT 2180.010 168.740 2456.790 168.880 ;
        RECT 2180.010 168.680 2180.330 168.740 ;
        RECT 2456.470 168.680 2456.790 168.740 ;
      LAYER via ;
        RECT 2174.520 503.240 2174.780 503.500 ;
        RECT 2180.040 503.240 2180.300 503.500 ;
        RECT 2180.040 168.680 2180.300 168.940 ;
        RECT 2456.500 168.680 2456.760 168.940 ;
      LAYER met2 ;
        RECT 2174.650 510.340 2174.930 514.000 ;
        RECT 2174.580 510.000 2174.930 510.340 ;
        RECT 2174.580 503.530 2174.720 510.000 ;
        RECT 2174.520 503.210 2174.780 503.530 ;
        RECT 2180.040 503.210 2180.300 503.530 ;
        RECT 2180.100 168.970 2180.240 503.210 ;
        RECT 2180.040 168.650 2180.300 168.970 ;
        RECT 2456.500 168.650 2456.760 168.970 ;
        RECT 2456.560 17.410 2456.700 168.650 ;
        RECT 2456.560 17.270 2459.000 17.410 ;
        RECT 2458.860 2.400 2459.000 17.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2186.910 176.020 2187.230 176.080 ;
        RECT 2470.270 176.020 2470.590 176.080 ;
        RECT 2186.910 175.880 2470.590 176.020 ;
        RECT 2186.910 175.820 2187.230 175.880 ;
        RECT 2470.270 175.820 2470.590 175.880 ;
        RECT 2470.270 17.580 2470.590 17.640 ;
        RECT 2476.710 17.580 2477.030 17.640 ;
        RECT 2470.270 17.440 2477.030 17.580 ;
        RECT 2470.270 17.380 2470.590 17.440 ;
        RECT 2476.710 17.380 2477.030 17.440 ;
      LAYER via ;
        RECT 2186.940 175.820 2187.200 176.080 ;
        RECT 2470.300 175.820 2470.560 176.080 ;
        RECT 2470.300 17.380 2470.560 17.640 ;
        RECT 2476.740 17.380 2477.000 17.640 ;
      LAYER met2 ;
        RECT 2187.070 510.340 2187.350 514.000 ;
        RECT 2187.000 510.000 2187.350 510.340 ;
        RECT 2187.000 176.110 2187.140 510.000 ;
        RECT 2186.940 175.790 2187.200 176.110 ;
        RECT 2470.300 175.790 2470.560 176.110 ;
        RECT 2470.360 17.670 2470.500 175.790 ;
        RECT 2470.300 17.350 2470.560 17.670 ;
        RECT 2476.740 17.350 2477.000 17.670 ;
        RECT 2476.800 2.400 2476.940 17.350 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2199.865 338.045 2200.035 386.155 ;
        RECT 2199.405 241.485 2199.575 289.255 ;
        RECT 2199.405 193.205 2199.575 207.315 ;
      LAYER mcon ;
        RECT 2199.865 385.985 2200.035 386.155 ;
        RECT 2199.405 289.085 2199.575 289.255 ;
        RECT 2199.405 207.145 2199.575 207.315 ;
      LAYER met1 ;
        RECT 2199.330 400.220 2199.650 400.480 ;
        RECT 2199.420 399.740 2199.560 400.220 ;
        RECT 2199.790 399.740 2200.110 399.800 ;
        RECT 2199.420 399.600 2200.110 399.740 ;
        RECT 2199.790 399.540 2200.110 399.600 ;
        RECT 2199.790 386.140 2200.110 386.200 ;
        RECT 2199.595 386.000 2200.110 386.140 ;
        RECT 2199.790 385.940 2200.110 386.000 ;
        RECT 2199.805 338.200 2200.095 338.245 ;
        RECT 2200.250 338.200 2200.570 338.260 ;
        RECT 2199.805 338.060 2200.570 338.200 ;
        RECT 2199.805 338.015 2200.095 338.060 ;
        RECT 2200.250 338.000 2200.570 338.060 ;
        RECT 2199.330 289.920 2199.650 289.980 ;
        RECT 2199.790 289.920 2200.110 289.980 ;
        RECT 2199.330 289.780 2200.110 289.920 ;
        RECT 2199.330 289.720 2199.650 289.780 ;
        RECT 2199.790 289.720 2200.110 289.780 ;
        RECT 2199.330 289.240 2199.650 289.300 ;
        RECT 2199.135 289.100 2199.650 289.240 ;
        RECT 2199.330 289.040 2199.650 289.100 ;
        RECT 2199.345 241.640 2199.635 241.685 ;
        RECT 2199.790 241.640 2200.110 241.700 ;
        RECT 2199.345 241.500 2200.110 241.640 ;
        RECT 2199.345 241.455 2199.635 241.500 ;
        RECT 2199.790 241.440 2200.110 241.500 ;
        RECT 2199.345 207.300 2199.635 207.345 ;
        RECT 2199.790 207.300 2200.110 207.360 ;
        RECT 2199.345 207.160 2200.110 207.300 ;
        RECT 2199.345 207.115 2199.635 207.160 ;
        RECT 2199.790 207.100 2200.110 207.160 ;
        RECT 2199.330 193.360 2199.650 193.420 ;
        RECT 2199.135 193.220 2199.650 193.360 ;
        RECT 2199.330 193.160 2199.650 193.220 ;
        RECT 2199.330 182.820 2199.650 182.880 ;
        RECT 2490.970 182.820 2491.290 182.880 ;
        RECT 2199.330 182.680 2491.290 182.820 ;
        RECT 2199.330 182.620 2199.650 182.680 ;
        RECT 2490.970 182.620 2491.290 182.680 ;
      LAYER via ;
        RECT 2199.360 400.220 2199.620 400.480 ;
        RECT 2199.820 399.540 2200.080 399.800 ;
        RECT 2199.820 385.940 2200.080 386.200 ;
        RECT 2200.280 338.000 2200.540 338.260 ;
        RECT 2199.360 289.720 2199.620 289.980 ;
        RECT 2199.820 289.720 2200.080 289.980 ;
        RECT 2199.360 289.040 2199.620 289.300 ;
        RECT 2199.820 241.440 2200.080 241.700 ;
        RECT 2199.820 207.100 2200.080 207.360 ;
        RECT 2199.360 193.160 2199.620 193.420 ;
        RECT 2199.360 182.620 2199.620 182.880 ;
        RECT 2491.000 182.620 2491.260 182.880 ;
      LAYER met2 ;
        RECT 2199.950 510.410 2200.230 514.000 ;
        RECT 2199.420 510.270 2200.230 510.410 ;
        RECT 2199.420 483.325 2199.560 510.270 ;
        RECT 2199.950 510.000 2200.230 510.270 ;
        RECT 2199.350 482.955 2199.630 483.325 ;
        RECT 2200.270 482.955 2200.550 483.325 ;
        RECT 2200.340 448.530 2200.480 482.955 ;
        RECT 2199.420 448.390 2200.480 448.530 ;
        RECT 2199.420 400.510 2199.560 448.390 ;
        RECT 2199.360 400.190 2199.620 400.510 ;
        RECT 2199.820 399.510 2200.080 399.830 ;
        RECT 2199.880 386.230 2200.020 399.510 ;
        RECT 2199.820 385.910 2200.080 386.230 ;
        RECT 2200.280 337.970 2200.540 338.290 ;
        RECT 2200.340 337.690 2200.480 337.970 ;
        RECT 2199.880 337.550 2200.480 337.690 ;
        RECT 2199.880 290.010 2200.020 337.550 ;
        RECT 2199.360 289.690 2199.620 290.010 ;
        RECT 2199.820 289.690 2200.080 290.010 ;
        RECT 2199.420 289.330 2199.560 289.690 ;
        RECT 2199.360 289.010 2199.620 289.330 ;
        RECT 2199.820 241.410 2200.080 241.730 ;
        RECT 2199.880 207.390 2200.020 241.410 ;
        RECT 2199.820 207.070 2200.080 207.390 ;
        RECT 2199.360 193.130 2199.620 193.450 ;
        RECT 2199.420 182.910 2199.560 193.130 ;
        RECT 2199.360 182.590 2199.620 182.910 ;
        RECT 2491.000 182.590 2491.260 182.910 ;
        RECT 2491.060 17.410 2491.200 182.590 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 2199.350 483.000 2199.630 483.280 ;
        RECT 2200.270 483.000 2200.550 483.280 ;
      LAYER met3 ;
        RECT 2199.325 483.290 2199.655 483.305 ;
        RECT 2200.245 483.290 2200.575 483.305 ;
        RECT 2199.325 482.990 2200.575 483.290 ;
        RECT 2199.325 482.975 2199.655 482.990 ;
        RECT 2200.245 482.975 2200.575 482.990 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2214.050 189.620 2214.370 189.680 ;
        RECT 2511.670 189.620 2511.990 189.680 ;
        RECT 2214.050 189.480 2511.990 189.620 ;
        RECT 2214.050 189.420 2214.370 189.480 ;
        RECT 2511.670 189.420 2511.990 189.480 ;
      LAYER via ;
        RECT 2214.080 189.420 2214.340 189.680 ;
        RECT 2511.700 189.420 2511.960 189.680 ;
      LAYER met2 ;
        RECT 2212.830 510.410 2213.110 514.000 ;
        RECT 2212.830 510.270 2214.280 510.410 ;
        RECT 2212.830 510.000 2213.110 510.270 ;
        RECT 2214.140 189.710 2214.280 510.270 ;
        RECT 2214.080 189.390 2214.340 189.710 ;
        RECT 2511.700 189.390 2511.960 189.710 ;
        RECT 2511.760 17.410 2511.900 189.390 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 196.760 2228.630 196.820 ;
        RECT 2525.470 196.760 2525.790 196.820 ;
        RECT 2228.310 196.620 2525.790 196.760 ;
        RECT 2228.310 196.560 2228.630 196.620 ;
        RECT 2525.470 196.560 2525.790 196.620 ;
      LAYER via ;
        RECT 2228.340 196.560 2228.600 196.820 ;
        RECT 2525.500 196.560 2525.760 196.820 ;
      LAYER met2 ;
        RECT 2225.710 510.410 2225.990 514.000 ;
        RECT 2225.710 510.270 2228.540 510.410 ;
        RECT 2225.710 510.000 2225.990 510.270 ;
        RECT 2228.400 196.850 2228.540 510.270 ;
        RECT 2228.340 196.530 2228.600 196.850 ;
        RECT 2525.500 196.530 2525.760 196.850 ;
        RECT 2525.560 16.730 2525.700 196.530 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.400 2530.300 16.590 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2238.430 500.720 2238.750 500.780 ;
        RECT 2242.110 500.720 2242.430 500.780 ;
        RECT 2238.430 500.580 2242.430 500.720 ;
        RECT 2238.430 500.520 2238.750 500.580 ;
        RECT 2242.110 500.520 2242.430 500.580 ;
        RECT 2242.110 210.360 2242.430 210.420 ;
        RECT 2546.170 210.360 2546.490 210.420 ;
        RECT 2242.110 210.220 2546.490 210.360 ;
        RECT 2242.110 210.160 2242.430 210.220 ;
        RECT 2546.170 210.160 2546.490 210.220 ;
      LAYER via ;
        RECT 2238.460 500.520 2238.720 500.780 ;
        RECT 2242.140 500.520 2242.400 500.780 ;
        RECT 2242.140 210.160 2242.400 210.420 ;
        RECT 2546.200 210.160 2546.460 210.420 ;
      LAYER met2 ;
        RECT 2238.590 510.340 2238.870 514.000 ;
        RECT 2238.520 510.000 2238.870 510.340 ;
        RECT 2238.520 500.810 2238.660 510.000 ;
        RECT 2238.460 500.490 2238.720 500.810 ;
        RECT 2242.140 500.490 2242.400 500.810 ;
        RECT 2242.200 210.450 2242.340 500.490 ;
        RECT 2242.140 210.130 2242.400 210.450 ;
        RECT 2546.200 210.130 2546.460 210.450 ;
        RECT 2546.260 17.410 2546.400 210.130 ;
        RECT 2546.260 17.270 2548.240 17.410 ;
        RECT 2548.100 2.400 2548.240 17.270 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2251.310 499.020 2251.630 499.080 ;
        RECT 2259.590 499.020 2259.910 499.080 ;
        RECT 2251.310 498.880 2259.910 499.020 ;
        RECT 2251.310 498.820 2251.630 498.880 ;
        RECT 2259.590 498.820 2259.910 498.880 ;
        RECT 2259.590 224.300 2259.910 224.360 ;
        RECT 2559.970 224.300 2560.290 224.360 ;
        RECT 2259.590 224.160 2560.290 224.300 ;
        RECT 2259.590 224.100 2259.910 224.160 ;
        RECT 2559.970 224.100 2560.290 224.160 ;
        RECT 2559.970 16.900 2560.290 16.960 ;
        RECT 2565.950 16.900 2566.270 16.960 ;
        RECT 2559.970 16.760 2566.270 16.900 ;
        RECT 2559.970 16.700 2560.290 16.760 ;
        RECT 2565.950 16.700 2566.270 16.760 ;
      LAYER via ;
        RECT 2251.340 498.820 2251.600 499.080 ;
        RECT 2259.620 498.820 2259.880 499.080 ;
        RECT 2259.620 224.100 2259.880 224.360 ;
        RECT 2560.000 224.100 2560.260 224.360 ;
        RECT 2560.000 16.700 2560.260 16.960 ;
        RECT 2565.980 16.700 2566.240 16.960 ;
      LAYER met2 ;
        RECT 2251.470 510.340 2251.750 514.000 ;
        RECT 2251.400 510.000 2251.750 510.340 ;
        RECT 2251.400 499.110 2251.540 510.000 ;
        RECT 2251.340 498.790 2251.600 499.110 ;
        RECT 2259.620 498.790 2259.880 499.110 ;
        RECT 2259.680 224.390 2259.820 498.790 ;
        RECT 2259.620 224.070 2259.880 224.390 ;
        RECT 2560.000 224.070 2560.260 224.390 ;
        RECT 2560.060 16.990 2560.200 224.070 ;
        RECT 2560.000 16.670 2560.260 16.990 ;
        RECT 2565.980 16.670 2566.240 16.990 ;
        RECT 2566.040 2.400 2566.180 16.670 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2263.730 503.440 2264.050 503.500 ;
        RECT 2269.250 503.440 2269.570 503.500 ;
        RECT 2263.730 503.300 2269.570 503.440 ;
        RECT 2263.730 503.240 2264.050 503.300 ;
        RECT 2269.250 503.240 2269.570 503.300 ;
        RECT 2269.250 410.620 2269.570 410.680 ;
        RECT 2580.670 410.620 2580.990 410.680 ;
        RECT 2269.250 410.480 2580.990 410.620 ;
        RECT 2269.250 410.420 2269.570 410.480 ;
        RECT 2580.670 410.420 2580.990 410.480 ;
      LAYER via ;
        RECT 2263.760 503.240 2264.020 503.500 ;
        RECT 2269.280 503.240 2269.540 503.500 ;
        RECT 2269.280 410.420 2269.540 410.680 ;
        RECT 2580.700 410.420 2580.960 410.680 ;
      LAYER met2 ;
        RECT 2263.890 510.340 2264.170 514.000 ;
        RECT 2263.820 510.000 2264.170 510.340 ;
        RECT 2263.820 503.530 2263.960 510.000 ;
        RECT 2263.760 503.210 2264.020 503.530 ;
        RECT 2269.280 503.210 2269.540 503.530 ;
        RECT 2269.340 410.710 2269.480 503.210 ;
        RECT 2269.280 410.390 2269.540 410.710 ;
        RECT 2580.700 410.390 2580.960 410.710 ;
        RECT 2580.760 17.410 2580.900 410.390 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 820.710 113.800 821.030 113.860 ;
        RECT 993.670 113.800 993.990 113.860 ;
        RECT 820.710 113.660 993.990 113.800 ;
        RECT 820.710 113.600 821.030 113.660 ;
        RECT 993.670 113.600 993.990 113.660 ;
        RECT 817.490 20.640 817.810 20.700 ;
        RECT 820.710 20.640 821.030 20.700 ;
        RECT 817.490 20.500 821.030 20.640 ;
        RECT 817.490 20.440 817.810 20.500 ;
        RECT 820.710 20.440 821.030 20.500 ;
      LAYER via ;
        RECT 820.740 113.600 821.000 113.860 ;
        RECT 993.700 113.600 993.960 113.860 ;
        RECT 817.520 20.440 817.780 20.700 ;
        RECT 820.740 20.440 821.000 20.700 ;
      LAYER met2 ;
        RECT 996.590 510.410 996.870 514.000 ;
        RECT 993.760 510.270 996.870 510.410 ;
        RECT 993.760 113.890 993.900 510.270 ;
        RECT 996.590 510.000 996.870 510.270 ;
        RECT 820.740 113.570 821.000 113.890 ;
        RECT 993.700 113.570 993.960 113.890 ;
        RECT 820.800 20.730 820.940 113.570 ;
        RECT 817.520 20.410 817.780 20.730 ;
        RECT 820.740 20.410 821.000 20.730 ;
        RECT 817.580 2.400 817.720 20.410 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2276.610 403.480 2276.930 403.540 ;
        RECT 2601.370 403.480 2601.690 403.540 ;
        RECT 2276.610 403.340 2601.690 403.480 ;
        RECT 2276.610 403.280 2276.930 403.340 ;
        RECT 2601.370 403.280 2601.690 403.340 ;
      LAYER via ;
        RECT 2276.640 403.280 2276.900 403.540 ;
        RECT 2601.400 403.280 2601.660 403.540 ;
      LAYER met2 ;
        RECT 2276.770 510.340 2277.050 514.000 ;
        RECT 2276.700 510.000 2277.050 510.340 ;
        RECT 2276.700 403.570 2276.840 510.000 ;
        RECT 2276.640 403.250 2276.900 403.570 ;
        RECT 2601.400 403.250 2601.660 403.570 ;
        RECT 2601.460 2.400 2601.600 403.250 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2290.410 99.860 2290.730 99.920 ;
        RECT 2615.170 99.860 2615.490 99.920 ;
        RECT 2290.410 99.720 2615.490 99.860 ;
        RECT 2290.410 99.660 2290.730 99.720 ;
        RECT 2615.170 99.660 2615.490 99.720 ;
      LAYER via ;
        RECT 2290.440 99.660 2290.700 99.920 ;
        RECT 2615.200 99.660 2615.460 99.920 ;
      LAYER met2 ;
        RECT 2289.650 510.410 2289.930 514.000 ;
        RECT 2289.650 510.270 2290.640 510.410 ;
        RECT 2289.650 510.000 2289.930 510.270 ;
        RECT 2290.500 99.950 2290.640 510.270 ;
        RECT 2290.440 99.630 2290.700 99.950 ;
        RECT 2615.200 99.630 2615.460 99.950 ;
        RECT 2615.260 17.410 2615.400 99.630 ;
        RECT 2615.260 17.270 2619.540 17.410 ;
        RECT 2619.400 2.400 2619.540 17.270 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2303.750 396.680 2304.070 396.740 ;
        RECT 2635.870 396.680 2636.190 396.740 ;
        RECT 2303.750 396.540 2636.190 396.680 ;
        RECT 2303.750 396.480 2304.070 396.540 ;
        RECT 2635.870 396.480 2636.190 396.540 ;
      LAYER via ;
        RECT 2303.780 396.480 2304.040 396.740 ;
        RECT 2635.900 396.480 2636.160 396.740 ;
      LAYER met2 ;
        RECT 2302.530 510.410 2302.810 514.000 ;
        RECT 2302.530 510.270 2303.980 510.410 ;
        RECT 2302.530 510.000 2302.810 510.270 ;
        RECT 2303.840 396.770 2303.980 510.270 ;
        RECT 2303.780 396.450 2304.040 396.770 ;
        RECT 2635.900 396.450 2636.160 396.770 ;
        RECT 2635.960 17.410 2636.100 396.450 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 107.000 2318.330 107.060 ;
        RECT 2649.670 107.000 2649.990 107.060 ;
        RECT 2318.010 106.860 2649.990 107.000 ;
        RECT 2318.010 106.800 2318.330 106.860 ;
        RECT 2649.670 106.800 2649.990 106.860 ;
      LAYER via ;
        RECT 2318.040 106.800 2318.300 107.060 ;
        RECT 2649.700 106.800 2649.960 107.060 ;
      LAYER met2 ;
        RECT 2315.410 510.410 2315.690 514.000 ;
        RECT 2315.410 510.270 2318.240 510.410 ;
        RECT 2315.410 510.000 2315.690 510.270 ;
        RECT 2318.100 107.090 2318.240 510.270 ;
        RECT 2318.040 106.770 2318.300 107.090 ;
        RECT 2649.700 106.770 2649.960 107.090 ;
        RECT 2649.760 17.410 2649.900 106.770 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2331.810 217.160 2332.130 217.220 ;
        RECT 2670.370 217.160 2670.690 217.220 ;
        RECT 2331.810 217.020 2670.690 217.160 ;
        RECT 2331.810 216.960 2332.130 217.020 ;
        RECT 2670.370 216.960 2670.690 217.020 ;
      LAYER via ;
        RECT 2331.840 216.960 2332.100 217.220 ;
        RECT 2670.400 216.960 2670.660 217.220 ;
      LAYER met2 ;
        RECT 2328.290 510.410 2328.570 514.000 ;
        RECT 2328.290 510.270 2332.040 510.410 ;
        RECT 2328.290 510.000 2328.570 510.270 ;
        RECT 2331.900 217.250 2332.040 510.270 ;
        RECT 2331.840 216.930 2332.100 217.250 ;
        RECT 2670.400 216.930 2670.660 217.250 ;
        RECT 2670.460 17.410 2670.600 216.930 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2340.550 503.440 2340.870 503.500 ;
        RECT 2349.290 503.440 2349.610 503.500 ;
        RECT 2340.550 503.300 2349.610 503.440 ;
        RECT 2340.550 503.240 2340.870 503.300 ;
        RECT 2349.290 503.240 2349.610 503.300 ;
        RECT 2349.290 113.800 2349.610 113.860 ;
        RECT 2684.630 113.800 2684.950 113.860 ;
        RECT 2349.290 113.660 2684.950 113.800 ;
        RECT 2349.290 113.600 2349.610 113.660 ;
        RECT 2684.630 113.600 2684.950 113.660 ;
        RECT 2684.630 20.980 2684.950 21.040 ;
        RECT 2690.610 20.980 2690.930 21.040 ;
        RECT 2684.630 20.840 2690.930 20.980 ;
        RECT 2684.630 20.780 2684.950 20.840 ;
        RECT 2690.610 20.780 2690.930 20.840 ;
      LAYER via ;
        RECT 2340.580 503.240 2340.840 503.500 ;
        RECT 2349.320 503.240 2349.580 503.500 ;
        RECT 2349.320 113.600 2349.580 113.860 ;
        RECT 2684.660 113.600 2684.920 113.860 ;
        RECT 2684.660 20.780 2684.920 21.040 ;
        RECT 2690.640 20.780 2690.900 21.040 ;
      LAYER met2 ;
        RECT 2340.710 510.340 2340.990 514.000 ;
        RECT 2340.640 510.000 2340.990 510.340 ;
        RECT 2340.640 503.530 2340.780 510.000 ;
        RECT 2340.580 503.210 2340.840 503.530 ;
        RECT 2349.320 503.210 2349.580 503.530 ;
        RECT 2349.380 113.890 2349.520 503.210 ;
        RECT 2349.320 113.570 2349.580 113.890 ;
        RECT 2684.660 113.570 2684.920 113.890 ;
        RECT 2684.720 21.070 2684.860 113.570 ;
        RECT 2684.660 20.750 2684.920 21.070 ;
        RECT 2690.640 20.750 2690.900 21.070 ;
        RECT 2690.700 2.400 2690.840 20.750 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2353.430 503.100 2353.750 503.160 ;
        RECT 2359.410 503.100 2359.730 503.160 ;
        RECT 2353.430 502.960 2359.730 503.100 ;
        RECT 2353.430 502.900 2353.750 502.960 ;
        RECT 2359.410 502.900 2359.730 502.960 ;
        RECT 2359.410 127.740 2359.730 127.800 ;
        RECT 2704.870 127.740 2705.190 127.800 ;
        RECT 2359.410 127.600 2705.190 127.740 ;
        RECT 2359.410 127.540 2359.730 127.600 ;
        RECT 2704.870 127.540 2705.190 127.600 ;
      LAYER via ;
        RECT 2353.460 502.900 2353.720 503.160 ;
        RECT 2359.440 502.900 2359.700 503.160 ;
        RECT 2359.440 127.540 2359.700 127.800 ;
        RECT 2704.900 127.540 2705.160 127.800 ;
      LAYER met2 ;
        RECT 2353.590 510.340 2353.870 514.000 ;
        RECT 2353.520 510.000 2353.870 510.340 ;
        RECT 2353.520 503.190 2353.660 510.000 ;
        RECT 2353.460 502.870 2353.720 503.190 ;
        RECT 2359.440 502.870 2359.700 503.190 ;
        RECT 2359.500 127.830 2359.640 502.870 ;
        RECT 2359.440 127.510 2359.700 127.830 ;
        RECT 2704.900 127.510 2705.160 127.830 ;
        RECT 2704.960 16.730 2705.100 127.510 ;
        RECT 2704.960 16.590 2708.780 16.730 ;
        RECT 2708.640 2.400 2708.780 16.590 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2366.310 231.100 2366.630 231.160 ;
        RECT 2725.570 231.100 2725.890 231.160 ;
        RECT 2366.310 230.960 2725.890 231.100 ;
        RECT 2366.310 230.900 2366.630 230.960 ;
        RECT 2725.570 230.900 2725.890 230.960 ;
      LAYER via ;
        RECT 2366.340 230.900 2366.600 231.160 ;
        RECT 2725.600 230.900 2725.860 231.160 ;
      LAYER met2 ;
        RECT 2366.470 510.340 2366.750 514.000 ;
        RECT 2366.400 510.000 2366.750 510.340 ;
        RECT 2366.400 231.190 2366.540 510.000 ;
        RECT 2366.340 230.870 2366.600 231.190 ;
        RECT 2725.600 230.870 2725.860 231.190 ;
        RECT 2725.660 16.730 2725.800 230.870 ;
        RECT 2725.660 16.590 2726.720 16.730 ;
        RECT 2726.580 2.400 2726.720 16.590 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2380.110 141.340 2380.430 141.400 ;
        RECT 2739.370 141.340 2739.690 141.400 ;
        RECT 2380.110 141.200 2739.690 141.340 ;
        RECT 2380.110 141.140 2380.430 141.200 ;
        RECT 2739.370 141.140 2739.690 141.200 ;
      LAYER via ;
        RECT 2380.140 141.140 2380.400 141.400 ;
        RECT 2739.400 141.140 2739.660 141.400 ;
      LAYER met2 ;
        RECT 2379.350 510.410 2379.630 514.000 ;
        RECT 2379.350 510.270 2380.340 510.410 ;
        RECT 2379.350 510.000 2379.630 510.270 ;
        RECT 2380.200 141.430 2380.340 510.270 ;
        RECT 2380.140 141.110 2380.400 141.430 ;
        RECT 2739.400 141.110 2739.660 141.430 ;
        RECT 2739.460 17.410 2739.600 141.110 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2393.450 389.880 2393.770 389.940 ;
        RECT 2760.070 389.880 2760.390 389.940 ;
        RECT 2393.450 389.740 2760.390 389.880 ;
        RECT 2393.450 389.680 2393.770 389.740 ;
        RECT 2760.070 389.680 2760.390 389.740 ;
      LAYER via ;
        RECT 2393.480 389.680 2393.740 389.940 ;
        RECT 2760.100 389.680 2760.360 389.940 ;
      LAYER met2 ;
        RECT 2392.230 510.410 2392.510 514.000 ;
        RECT 2392.230 510.270 2393.680 510.410 ;
        RECT 2392.230 510.000 2392.510 510.270 ;
        RECT 2393.540 389.970 2393.680 510.270 ;
        RECT 2393.480 389.650 2393.740 389.970 ;
        RECT 2760.100 389.650 2760.360 389.970 ;
        RECT 2760.160 17.410 2760.300 389.650 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1003.790 502.080 1004.110 502.140 ;
        RECT 1008.850 502.080 1009.170 502.140 ;
        RECT 1003.790 501.940 1009.170 502.080 ;
        RECT 1003.790 501.880 1004.110 501.940 ;
        RECT 1008.850 501.880 1009.170 501.940 ;
        RECT 840.950 120.600 841.270 120.660 ;
        RECT 1003.790 120.600 1004.110 120.660 ;
        RECT 840.950 120.460 1004.110 120.600 ;
        RECT 840.950 120.400 841.270 120.460 ;
        RECT 1003.790 120.400 1004.110 120.460 ;
        RECT 835.430 20.640 835.750 20.700 ;
        RECT 840.950 20.640 841.270 20.700 ;
        RECT 835.430 20.500 841.270 20.640 ;
        RECT 835.430 20.440 835.750 20.500 ;
        RECT 840.950 20.440 841.270 20.500 ;
      LAYER via ;
        RECT 1003.820 501.880 1004.080 502.140 ;
        RECT 1008.880 501.880 1009.140 502.140 ;
        RECT 840.980 120.400 841.240 120.660 ;
        RECT 1003.820 120.400 1004.080 120.660 ;
        RECT 835.460 20.440 835.720 20.700 ;
        RECT 840.980 20.440 841.240 20.700 ;
      LAYER met2 ;
        RECT 1009.010 510.340 1009.290 514.000 ;
        RECT 1008.940 510.000 1009.290 510.340 ;
        RECT 1008.940 502.170 1009.080 510.000 ;
        RECT 1003.820 501.850 1004.080 502.170 ;
        RECT 1008.880 501.850 1009.140 502.170 ;
        RECT 1003.880 120.690 1004.020 501.850 ;
        RECT 840.980 120.370 841.240 120.690 ;
        RECT 1003.820 120.370 1004.080 120.690 ;
        RECT 841.040 20.730 841.180 120.370 ;
        RECT 835.460 20.410 835.720 20.730 ;
        RECT 840.980 20.410 841.240 20.730 ;
        RECT 835.520 2.400 835.660 20.410 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2407.710 155.280 2408.030 155.340 ;
        RECT 2774.330 155.280 2774.650 155.340 ;
        RECT 2407.710 155.140 2774.650 155.280 ;
        RECT 2407.710 155.080 2408.030 155.140 ;
        RECT 2774.330 155.080 2774.650 155.140 ;
      LAYER via ;
        RECT 2407.740 155.080 2408.000 155.340 ;
        RECT 2774.360 155.080 2774.620 155.340 ;
      LAYER met2 ;
        RECT 2405.110 510.410 2405.390 514.000 ;
        RECT 2405.110 510.270 2407.940 510.410 ;
        RECT 2405.110 510.000 2405.390 510.270 ;
        RECT 2407.800 155.370 2407.940 510.270 ;
        RECT 2407.740 155.050 2408.000 155.370 ;
        RECT 2774.360 155.050 2774.620 155.370 ;
        RECT 2774.420 17.410 2774.560 155.050 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2417.370 496.980 2417.690 497.040 ;
        RECT 2421.510 496.980 2421.830 497.040 ;
        RECT 2417.370 496.840 2421.830 496.980 ;
        RECT 2417.370 496.780 2417.690 496.840 ;
        RECT 2421.510 496.780 2421.830 496.840 ;
        RECT 2421.510 245.040 2421.830 245.100 ;
        RECT 2794.570 245.040 2794.890 245.100 ;
        RECT 2421.510 244.900 2794.890 245.040 ;
        RECT 2421.510 244.840 2421.830 244.900 ;
        RECT 2794.570 244.840 2794.890 244.900 ;
      LAYER via ;
        RECT 2417.400 496.780 2417.660 497.040 ;
        RECT 2421.540 496.780 2421.800 497.040 ;
        RECT 2421.540 244.840 2421.800 245.100 ;
        RECT 2794.600 244.840 2794.860 245.100 ;
      LAYER met2 ;
        RECT 2417.530 510.340 2417.810 514.000 ;
        RECT 2417.460 510.000 2417.810 510.340 ;
        RECT 2417.460 497.070 2417.600 510.000 ;
        RECT 2417.400 496.750 2417.660 497.070 ;
        RECT 2421.540 496.750 2421.800 497.070 ;
        RECT 2421.600 245.130 2421.740 496.750 ;
        RECT 2421.540 244.810 2421.800 245.130 ;
        RECT 2794.600 244.810 2794.860 245.130 ;
        RECT 2794.660 17.410 2794.800 244.810 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2430.250 496.980 2430.570 497.040 ;
        RECT 2434.850 496.980 2435.170 497.040 ;
        RECT 2430.250 496.840 2435.170 496.980 ;
        RECT 2430.250 496.780 2430.570 496.840 ;
        RECT 2434.850 496.780 2435.170 496.840 ;
        RECT 2434.850 375.940 2435.170 376.000 ;
        RECT 2815.730 375.940 2816.050 376.000 ;
        RECT 2434.850 375.800 2816.050 375.940 ;
        RECT 2434.850 375.740 2435.170 375.800 ;
        RECT 2815.730 375.740 2816.050 375.800 ;
      LAYER via ;
        RECT 2430.280 496.780 2430.540 497.040 ;
        RECT 2434.880 496.780 2435.140 497.040 ;
        RECT 2434.880 375.740 2435.140 376.000 ;
        RECT 2815.760 375.740 2816.020 376.000 ;
      LAYER met2 ;
        RECT 2430.410 510.340 2430.690 514.000 ;
        RECT 2430.340 510.000 2430.690 510.340 ;
        RECT 2430.340 497.070 2430.480 510.000 ;
        RECT 2430.280 496.750 2430.540 497.070 ;
        RECT 2434.880 496.750 2435.140 497.070 ;
        RECT 2434.940 376.030 2435.080 496.750 ;
        RECT 2434.880 375.710 2435.140 376.030 ;
        RECT 2815.760 375.710 2816.020 376.030 ;
        RECT 2815.820 2.400 2815.960 375.710 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2443.130 496.980 2443.450 497.040 ;
        RECT 2448.650 496.980 2448.970 497.040 ;
        RECT 2443.130 496.840 2448.970 496.980 ;
        RECT 2443.130 496.780 2443.450 496.840 ;
        RECT 2448.650 496.780 2448.970 496.840 ;
        RECT 2448.650 162.080 2448.970 162.140 ;
        RECT 2829.070 162.080 2829.390 162.140 ;
        RECT 2448.650 161.940 2829.390 162.080 ;
        RECT 2448.650 161.880 2448.970 161.940 ;
        RECT 2829.070 161.880 2829.390 161.940 ;
      LAYER via ;
        RECT 2443.160 496.780 2443.420 497.040 ;
        RECT 2448.680 496.780 2448.940 497.040 ;
        RECT 2448.680 161.880 2448.940 162.140 ;
        RECT 2829.100 161.880 2829.360 162.140 ;
      LAYER met2 ;
        RECT 2443.290 510.340 2443.570 514.000 ;
        RECT 2443.220 510.000 2443.570 510.340 ;
        RECT 2443.220 497.070 2443.360 510.000 ;
        RECT 2443.160 496.750 2443.420 497.070 ;
        RECT 2448.680 496.750 2448.940 497.070 ;
        RECT 2448.740 162.170 2448.880 496.750 ;
        RECT 2448.680 161.850 2448.940 162.170 ;
        RECT 2829.100 161.850 2829.360 162.170 ;
        RECT 2829.160 17.410 2829.300 161.850 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2456.010 369.140 2456.330 369.200 ;
        RECT 2849.770 369.140 2850.090 369.200 ;
        RECT 2456.010 369.000 2850.090 369.140 ;
        RECT 2456.010 368.940 2456.330 369.000 ;
        RECT 2849.770 368.940 2850.090 369.000 ;
      LAYER via ;
        RECT 2456.040 368.940 2456.300 369.200 ;
        RECT 2849.800 368.940 2850.060 369.200 ;
      LAYER met2 ;
        RECT 2456.170 510.340 2456.450 514.000 ;
        RECT 2456.100 510.000 2456.450 510.340 ;
        RECT 2456.100 369.230 2456.240 510.000 ;
        RECT 2456.040 368.910 2456.300 369.230 ;
        RECT 2849.800 368.910 2850.060 369.230 ;
        RECT 2849.860 17.410 2850.000 368.910 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2469.810 168.880 2470.130 168.940 ;
        RECT 2863.570 168.880 2863.890 168.940 ;
        RECT 2469.810 168.740 2863.890 168.880 ;
        RECT 2469.810 168.680 2470.130 168.740 ;
        RECT 2863.570 168.680 2863.890 168.740 ;
      LAYER via ;
        RECT 2469.840 168.680 2470.100 168.940 ;
        RECT 2863.600 168.680 2863.860 168.940 ;
      LAYER met2 ;
        RECT 2469.050 510.410 2469.330 514.000 ;
        RECT 2469.050 510.270 2470.040 510.410 ;
        RECT 2469.050 510.000 2469.330 510.270 ;
        RECT 2469.900 168.970 2470.040 510.270 ;
        RECT 2469.840 168.650 2470.100 168.970 ;
        RECT 2863.600 168.650 2863.860 168.970 ;
        RECT 2863.660 17.410 2863.800 168.650 ;
        RECT 2863.660 17.270 2869.320 17.410 ;
        RECT 2869.180 2.400 2869.320 17.270 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2483.610 37.980 2483.930 38.040 ;
        RECT 2887.030 37.980 2887.350 38.040 ;
        RECT 2483.610 37.840 2887.350 37.980 ;
        RECT 2483.610 37.780 2483.930 37.840 ;
        RECT 2887.030 37.780 2887.350 37.840 ;
      LAYER via ;
        RECT 2483.640 37.780 2483.900 38.040 ;
        RECT 2887.060 37.780 2887.320 38.040 ;
      LAYER met2 ;
        RECT 2481.930 510.410 2482.210 514.000 ;
        RECT 2481.930 510.270 2483.840 510.410 ;
        RECT 2481.930 510.000 2482.210 510.270 ;
        RECT 2483.700 38.070 2483.840 510.270 ;
        RECT 2483.640 37.750 2483.900 38.070 ;
        RECT 2887.060 37.750 2887.320 38.070 ;
        RECT 2887.120 2.400 2887.260 37.750 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2497.410 44.780 2497.730 44.840 ;
        RECT 2904.970 44.780 2905.290 44.840 ;
        RECT 2497.410 44.640 2905.290 44.780 ;
        RECT 2497.410 44.580 2497.730 44.640 ;
        RECT 2904.970 44.580 2905.290 44.640 ;
      LAYER via ;
        RECT 2497.440 44.580 2497.700 44.840 ;
        RECT 2905.000 44.580 2905.260 44.840 ;
      LAYER met2 ;
        RECT 2494.350 510.410 2494.630 514.000 ;
        RECT 2494.350 510.270 2497.640 510.410 ;
        RECT 2494.350 510.000 2494.630 510.270 ;
        RECT 2497.500 44.870 2497.640 510.270 ;
        RECT 2497.440 44.550 2497.700 44.870 ;
        RECT 2905.000 44.550 2905.260 44.870 ;
        RECT 2905.060 2.400 2905.200 44.550 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 107.000 855.530 107.060 ;
        RECT 1021.730 107.000 1022.050 107.060 ;
        RECT 855.210 106.860 1022.050 107.000 ;
        RECT 855.210 106.800 855.530 106.860 ;
        RECT 1021.730 106.800 1022.050 106.860 ;
        RECT 852.910 20.640 853.230 20.700 ;
        RECT 855.210 20.640 855.530 20.700 ;
        RECT 852.910 20.500 855.530 20.640 ;
        RECT 852.910 20.440 853.230 20.500 ;
        RECT 855.210 20.440 855.530 20.500 ;
      LAYER via ;
        RECT 855.240 106.800 855.500 107.060 ;
        RECT 1021.760 106.800 1022.020 107.060 ;
        RECT 852.940 20.440 853.200 20.700 ;
        RECT 855.240 20.440 855.500 20.700 ;
      LAYER met2 ;
        RECT 1021.890 510.340 1022.170 514.000 ;
        RECT 1021.820 510.000 1022.170 510.340 ;
        RECT 1021.820 107.090 1021.960 510.000 ;
        RECT 855.240 106.770 855.500 107.090 ;
        RECT 1021.760 106.770 1022.020 107.090 ;
        RECT 855.300 20.730 855.440 106.770 ;
        RECT 852.940 20.410 853.200 20.730 ;
        RECT 855.240 20.410 855.500 20.730 ;
        RECT 853.000 2.400 853.140 20.410 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1028.630 401.100 1028.950 401.160 ;
        RECT 1032.310 401.100 1032.630 401.160 ;
        RECT 1028.630 400.960 1032.630 401.100 ;
        RECT 1028.630 400.900 1028.950 400.960 ;
        RECT 1032.310 400.900 1032.630 400.960 ;
        RECT 1028.630 241.300 1028.950 241.360 ;
        RECT 1029.090 241.300 1029.410 241.360 ;
        RECT 1028.630 241.160 1029.410 241.300 ;
        RECT 1028.630 241.100 1028.950 241.160 ;
        RECT 1029.090 241.100 1029.410 241.160 ;
        RECT 875.910 127.740 876.230 127.800 ;
        RECT 1028.630 127.740 1028.950 127.800 ;
        RECT 875.910 127.600 1028.950 127.740 ;
        RECT 875.910 127.540 876.230 127.600 ;
        RECT 1028.630 127.540 1028.950 127.600 ;
        RECT 870.850 20.640 871.170 20.700 ;
        RECT 875.910 20.640 876.230 20.700 ;
        RECT 870.850 20.500 876.230 20.640 ;
        RECT 870.850 20.440 871.170 20.500 ;
        RECT 875.910 20.440 876.230 20.500 ;
      LAYER via ;
        RECT 1028.660 400.900 1028.920 401.160 ;
        RECT 1032.340 400.900 1032.600 401.160 ;
        RECT 1028.660 241.100 1028.920 241.360 ;
        RECT 1029.120 241.100 1029.380 241.360 ;
        RECT 875.940 127.540 876.200 127.800 ;
        RECT 1028.660 127.540 1028.920 127.800 ;
        RECT 870.880 20.440 871.140 20.700 ;
        RECT 875.940 20.440 876.200 20.700 ;
      LAYER met2 ;
        RECT 1034.770 510.340 1035.050 514.000 ;
        RECT 1034.700 510.000 1035.050 510.340 ;
        RECT 1034.700 483.325 1034.840 510.000 ;
        RECT 1032.790 482.955 1033.070 483.325 ;
        RECT 1034.630 482.955 1034.910 483.325 ;
        RECT 1032.860 434.930 1033.000 482.955 ;
        RECT 1032.400 434.790 1033.000 434.930 ;
        RECT 1032.400 401.190 1032.540 434.790 ;
        RECT 1028.660 400.870 1028.920 401.190 ;
        RECT 1032.340 400.870 1032.600 401.190 ;
        RECT 1028.720 364.890 1028.860 400.870 ;
        RECT 1028.720 364.750 1029.780 364.890 ;
        RECT 1029.640 265.610 1029.780 364.750 ;
        RECT 1029.180 265.470 1029.780 265.610 ;
        RECT 1029.180 241.390 1029.320 265.470 ;
        RECT 1028.660 241.070 1028.920 241.390 ;
        RECT 1029.120 241.070 1029.380 241.390 ;
        RECT 1028.720 127.830 1028.860 241.070 ;
        RECT 875.940 127.510 876.200 127.830 ;
        RECT 1028.660 127.510 1028.920 127.830 ;
        RECT 876.000 20.730 876.140 127.510 ;
        RECT 870.880 20.410 871.140 20.730 ;
        RECT 875.940 20.410 876.200 20.730 ;
        RECT 870.940 2.400 871.080 20.410 ;
        RECT 870.730 -4.800 871.290 2.400 ;
      LAYER via2 ;
        RECT 1032.790 483.000 1033.070 483.280 ;
        RECT 1034.630 483.000 1034.910 483.280 ;
      LAYER met3 ;
        RECT 1032.765 483.290 1033.095 483.305 ;
        RECT 1034.605 483.290 1034.935 483.305 ;
        RECT 1032.765 482.990 1034.935 483.290 ;
        RECT 1032.765 482.975 1033.095 482.990 ;
        RECT 1034.605 482.975 1034.935 482.990 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1042.505 193.205 1042.675 241.315 ;
        RECT 888.865 2.805 889.035 14.195 ;
      LAYER mcon ;
        RECT 1042.505 241.145 1042.675 241.315 ;
        RECT 888.865 14.025 889.035 14.195 ;
      LAYER met1 ;
        RECT 1043.350 483.040 1043.670 483.100 ;
        RECT 1044.270 483.040 1044.590 483.100 ;
        RECT 1043.350 482.900 1044.590 483.040 ;
        RECT 1043.350 482.840 1043.670 482.900 ;
        RECT 1044.270 482.840 1044.590 482.900 ;
        RECT 1042.430 351.940 1042.750 352.200 ;
        RECT 1042.520 351.460 1042.660 351.940 ;
        RECT 1042.890 351.460 1043.210 351.520 ;
        RECT 1042.520 351.320 1043.210 351.460 ;
        RECT 1042.890 351.260 1043.210 351.320 ;
        RECT 1042.430 283.120 1042.750 283.180 ;
        RECT 1043.350 283.120 1043.670 283.180 ;
        RECT 1042.430 282.980 1043.670 283.120 ;
        RECT 1042.430 282.920 1042.750 282.980 ;
        RECT 1043.350 282.920 1043.670 282.980 ;
        RECT 1042.445 241.300 1042.735 241.345 ;
        RECT 1042.890 241.300 1043.210 241.360 ;
        RECT 1042.445 241.160 1043.210 241.300 ;
        RECT 1042.445 241.115 1042.735 241.160 ;
        RECT 1042.890 241.100 1043.210 241.160 ;
        RECT 1042.430 193.360 1042.750 193.420 ;
        RECT 1042.235 193.220 1042.750 193.360 ;
        RECT 1042.430 193.160 1042.750 193.220 ;
        RECT 889.710 134.540 890.030 134.600 ;
        RECT 1042.430 134.540 1042.750 134.600 ;
        RECT 889.710 134.400 1042.750 134.540 ;
        RECT 889.710 134.340 890.030 134.400 ;
        RECT 1042.430 134.340 1042.750 134.400 ;
        RECT 888.805 14.180 889.095 14.225 ;
        RECT 889.710 14.180 890.030 14.240 ;
        RECT 888.805 14.040 890.030 14.180 ;
        RECT 888.805 13.995 889.095 14.040 ;
        RECT 889.710 13.980 890.030 14.040 ;
        RECT 888.790 2.960 889.110 3.020 ;
        RECT 888.595 2.820 889.110 2.960 ;
        RECT 888.790 2.760 889.110 2.820 ;
      LAYER via ;
        RECT 1043.380 482.840 1043.640 483.100 ;
        RECT 1044.300 482.840 1044.560 483.100 ;
        RECT 1042.460 351.940 1042.720 352.200 ;
        RECT 1042.920 351.260 1043.180 351.520 ;
        RECT 1042.460 282.920 1042.720 283.180 ;
        RECT 1043.380 282.920 1043.640 283.180 ;
        RECT 1042.920 241.100 1043.180 241.360 ;
        RECT 1042.460 193.160 1042.720 193.420 ;
        RECT 889.740 134.340 890.000 134.600 ;
        RECT 1042.460 134.340 1042.720 134.600 ;
        RECT 889.740 13.980 890.000 14.240 ;
        RECT 888.820 2.760 889.080 3.020 ;
      LAYER met2 ;
        RECT 1047.650 510.340 1047.930 514.000 ;
        RECT 1047.580 510.000 1047.930 510.340 ;
        RECT 1047.580 483.325 1047.720 510.000 ;
        RECT 1043.380 482.810 1043.640 483.130 ;
        RECT 1044.290 482.955 1044.570 483.325 ;
        RECT 1047.510 482.955 1047.790 483.325 ;
        RECT 1044.300 482.810 1044.560 482.955 ;
        RECT 1043.440 434.930 1043.580 482.810 ;
        RECT 1042.520 434.790 1043.580 434.930 ;
        RECT 1042.520 352.230 1042.660 434.790 ;
        RECT 1042.460 351.910 1042.720 352.230 ;
        RECT 1042.920 351.230 1043.180 351.550 ;
        RECT 1042.980 304.370 1043.120 351.230 ;
        RECT 1042.980 304.230 1043.580 304.370 ;
        RECT 1043.440 283.210 1043.580 304.230 ;
        RECT 1042.460 282.890 1042.720 283.210 ;
        RECT 1043.380 282.890 1043.640 283.210 ;
        RECT 1042.520 265.610 1042.660 282.890 ;
        RECT 1042.520 265.470 1043.580 265.610 ;
        RECT 1043.440 254.730 1043.580 265.470 ;
        RECT 1042.980 254.590 1043.580 254.730 ;
        RECT 1042.980 241.390 1043.120 254.590 ;
        RECT 1042.920 241.070 1043.180 241.390 ;
        RECT 1042.460 193.130 1042.720 193.450 ;
        RECT 1042.520 134.630 1042.660 193.130 ;
        RECT 889.740 134.310 890.000 134.630 ;
        RECT 1042.460 134.310 1042.720 134.630 ;
        RECT 889.800 14.270 889.940 134.310 ;
        RECT 889.740 13.950 890.000 14.270 ;
        RECT 888.820 2.730 889.080 3.050 ;
        RECT 888.880 2.400 889.020 2.730 ;
        RECT 888.670 -4.800 889.230 2.400 ;
      LAYER via2 ;
        RECT 1044.290 483.000 1044.570 483.280 ;
        RECT 1047.510 483.000 1047.790 483.280 ;
      LAYER met3 ;
        RECT 1044.265 483.290 1044.595 483.305 ;
        RECT 1047.485 483.290 1047.815 483.305 ;
        RECT 1044.265 482.990 1047.815 483.290 ;
        RECT 1044.265 482.975 1044.595 482.990 ;
        RECT 1047.485 482.975 1047.815 482.990 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1057.150 483.720 1057.470 483.780 ;
        RECT 1060.370 483.720 1060.690 483.780 ;
        RECT 1057.150 483.580 1060.690 483.720 ;
        RECT 1057.150 483.520 1057.470 483.580 ;
        RECT 1060.370 483.520 1060.690 483.580 ;
        RECT 1056.690 193.360 1057.010 193.420 ;
        RECT 1057.610 193.360 1057.930 193.420 ;
        RECT 1056.690 193.220 1057.930 193.360 ;
        RECT 1056.690 193.160 1057.010 193.220 ;
        RECT 1057.610 193.160 1057.930 193.220 ;
        RECT 910.410 141.340 910.730 141.400 ;
        RECT 1056.690 141.340 1057.010 141.400 ;
        RECT 910.410 141.200 1057.010 141.340 ;
        RECT 910.410 141.140 910.730 141.200 ;
        RECT 1056.690 141.140 1057.010 141.200 ;
        RECT 906.730 16.220 907.050 16.280 ;
        RECT 910.410 16.220 910.730 16.280 ;
        RECT 906.730 16.080 910.730 16.220 ;
        RECT 906.730 16.020 907.050 16.080 ;
        RECT 910.410 16.020 910.730 16.080 ;
      LAYER via ;
        RECT 1057.180 483.520 1057.440 483.780 ;
        RECT 1060.400 483.520 1060.660 483.780 ;
        RECT 1056.720 193.160 1056.980 193.420 ;
        RECT 1057.640 193.160 1057.900 193.420 ;
        RECT 910.440 141.140 910.700 141.400 ;
        RECT 1056.720 141.140 1056.980 141.400 ;
        RECT 906.760 16.020 907.020 16.280 ;
        RECT 910.440 16.020 910.700 16.280 ;
      LAYER met2 ;
        RECT 1060.530 510.340 1060.810 514.000 ;
        RECT 1060.460 510.000 1060.810 510.340 ;
        RECT 1060.460 483.810 1060.600 510.000 ;
        RECT 1057.180 483.490 1057.440 483.810 ;
        RECT 1060.400 483.490 1060.660 483.810 ;
        RECT 1057.240 400.930 1057.380 483.490 ;
        RECT 1057.240 400.790 1057.840 400.930 ;
        RECT 1057.700 400.250 1057.840 400.790 ;
        RECT 1056.780 400.110 1057.840 400.250 ;
        RECT 1056.780 265.610 1056.920 400.110 ;
        RECT 1056.780 265.470 1057.380 265.610 ;
        RECT 1057.240 207.130 1057.380 265.470 ;
        RECT 1057.240 206.990 1057.840 207.130 ;
        RECT 1057.700 193.450 1057.840 206.990 ;
        RECT 1056.720 193.130 1056.980 193.450 ;
        RECT 1057.640 193.130 1057.900 193.450 ;
        RECT 1056.780 141.430 1056.920 193.130 ;
        RECT 910.440 141.110 910.700 141.430 ;
        RECT 1056.720 141.110 1056.980 141.430 ;
        RECT 910.500 16.310 910.640 141.110 ;
        RECT 906.760 15.990 907.020 16.310 ;
        RECT 910.440 15.990 910.700 16.310 ;
        RECT 906.820 2.400 906.960 15.990 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 86.600 924.530 86.660 ;
        RECT 1069.570 86.600 1069.890 86.660 ;
        RECT 924.210 86.460 1069.890 86.600 ;
        RECT 924.210 86.400 924.530 86.460 ;
        RECT 1069.570 86.400 1069.890 86.460 ;
      LAYER via ;
        RECT 924.240 86.400 924.500 86.660 ;
        RECT 1069.600 86.400 1069.860 86.660 ;
      LAYER met2 ;
        RECT 1073.410 510.410 1073.690 514.000 ;
        RECT 1069.660 510.270 1073.690 510.410 ;
        RECT 1069.660 86.690 1069.800 510.270 ;
        RECT 1073.410 510.000 1073.690 510.270 ;
        RECT 924.240 86.370 924.500 86.690 ;
        RECT 1069.600 86.370 1069.860 86.690 ;
        RECT 924.300 2.400 924.440 86.370 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.910 148.140 945.230 148.200 ;
        RECT 1083.370 148.140 1083.690 148.200 ;
        RECT 944.910 148.000 1083.690 148.140 ;
        RECT 944.910 147.940 945.230 148.000 ;
        RECT 1083.370 147.940 1083.690 148.000 ;
        RECT 942.150 16.900 942.470 16.960 ;
        RECT 944.910 16.900 945.230 16.960 ;
        RECT 942.150 16.760 945.230 16.900 ;
        RECT 942.150 16.700 942.470 16.760 ;
        RECT 944.910 16.700 945.230 16.760 ;
      LAYER via ;
        RECT 944.940 147.940 945.200 148.200 ;
        RECT 1083.400 147.940 1083.660 148.200 ;
        RECT 942.180 16.700 942.440 16.960 ;
        RECT 944.940 16.700 945.200 16.960 ;
      LAYER met2 ;
        RECT 1085.830 510.410 1086.110 514.000 ;
        RECT 1083.460 510.270 1086.110 510.410 ;
        RECT 1083.460 148.230 1083.600 510.270 ;
        RECT 1085.830 510.000 1086.110 510.270 ;
        RECT 944.940 147.910 945.200 148.230 ;
        RECT 1083.400 147.910 1083.660 148.230 ;
        RECT 945.000 16.990 945.140 147.910 ;
        RECT 942.180 16.670 942.440 16.990 ;
        RECT 944.940 16.670 945.200 16.990 ;
        RECT 942.240 2.400 942.380 16.670 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1072.790 496.980 1073.110 497.040 ;
        RECT 1098.550 496.980 1098.870 497.040 ;
        RECT 1072.790 496.840 1098.870 496.980 ;
        RECT 1072.790 496.780 1073.110 496.840 ;
        RECT 1098.550 496.780 1098.870 496.840 ;
        RECT 965.610 93.400 965.930 93.460 ;
        RECT 1072.790 93.400 1073.110 93.460 ;
        RECT 965.610 93.260 1073.110 93.400 ;
        RECT 965.610 93.200 965.930 93.260 ;
        RECT 1072.790 93.200 1073.110 93.260 ;
        RECT 960.090 16.900 960.410 16.960 ;
        RECT 965.610 16.900 965.930 16.960 ;
        RECT 960.090 16.760 965.930 16.900 ;
        RECT 960.090 16.700 960.410 16.760 ;
        RECT 965.610 16.700 965.930 16.760 ;
      LAYER via ;
        RECT 1072.820 496.780 1073.080 497.040 ;
        RECT 1098.580 496.780 1098.840 497.040 ;
        RECT 965.640 93.200 965.900 93.460 ;
        RECT 1072.820 93.200 1073.080 93.460 ;
        RECT 960.120 16.700 960.380 16.960 ;
        RECT 965.640 16.700 965.900 16.960 ;
      LAYER met2 ;
        RECT 1098.710 510.340 1098.990 514.000 ;
        RECT 1098.640 510.000 1098.990 510.340 ;
        RECT 1098.640 497.070 1098.780 510.000 ;
        RECT 1072.820 496.750 1073.080 497.070 ;
        RECT 1098.580 496.750 1098.840 497.070 ;
        RECT 1072.880 93.490 1073.020 496.750 ;
        RECT 965.640 93.170 965.900 93.490 ;
        RECT 1072.820 93.170 1073.080 93.490 ;
        RECT 965.700 16.990 965.840 93.170 ;
        RECT 960.120 16.670 960.380 16.990 ;
        RECT 965.640 16.670 965.900 16.990 ;
        RECT 960.180 2.400 960.320 16.670 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 979.410 99.860 979.730 99.920 ;
        RECT 1111.430 99.860 1111.750 99.920 ;
        RECT 979.410 99.720 1111.750 99.860 ;
        RECT 979.410 99.660 979.730 99.720 ;
        RECT 1111.430 99.660 1111.750 99.720 ;
      LAYER via ;
        RECT 979.440 99.660 979.700 99.920 ;
        RECT 1111.460 99.660 1111.720 99.920 ;
      LAYER met2 ;
        RECT 1111.590 510.340 1111.870 514.000 ;
        RECT 1111.520 510.000 1111.870 510.340 ;
        RECT 1111.520 99.950 1111.660 510.000 ;
        RECT 979.440 99.630 979.700 99.950 ;
        RECT 1111.460 99.630 1111.720 99.950 ;
        RECT 979.500 17.410 979.640 99.630 ;
        RECT 978.120 17.270 979.640 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 877.750 449.040 878.070 449.100 ;
        RECT 877.380 448.900 878.070 449.040 ;
        RECT 877.380 448.760 877.520 448.900 ;
        RECT 877.750 448.840 878.070 448.900 ;
        RECT 877.290 448.500 877.610 448.760 ;
        RECT 877.290 351.940 877.610 352.200 ;
        RECT 877.380 351.460 877.520 351.940 ;
        RECT 877.750 351.460 878.070 351.520 ;
        RECT 877.380 351.320 878.070 351.460 ;
        RECT 877.750 351.260 878.070 351.320 ;
        RECT 876.830 303.520 877.150 303.580 ;
        RECT 877.750 303.520 878.070 303.580 ;
        RECT 876.830 303.380 878.070 303.520 ;
        RECT 876.830 303.320 877.150 303.380 ;
        RECT 877.750 303.320 878.070 303.380 ;
        RECT 877.750 255.580 878.070 255.640 ;
        RECT 876.920 255.440 878.070 255.580 ;
        RECT 876.920 255.300 877.060 255.440 ;
        RECT 877.750 255.380 878.070 255.440 ;
        RECT 876.830 255.040 877.150 255.300 ;
        RECT 662.010 134.540 662.330 134.600 ;
        RECT 877.290 134.540 877.610 134.600 ;
        RECT 662.010 134.400 877.610 134.540 ;
        RECT 662.010 134.340 662.330 134.400 ;
        RECT 877.290 134.340 877.610 134.400 ;
        RECT 656.950 16.900 657.270 16.960 ;
        RECT 662.010 16.900 662.330 16.960 ;
        RECT 656.950 16.760 662.330 16.900 ;
        RECT 656.950 16.700 657.270 16.760 ;
        RECT 662.010 16.700 662.330 16.760 ;
      LAYER via ;
        RECT 877.780 448.840 878.040 449.100 ;
        RECT 877.320 448.500 877.580 448.760 ;
        RECT 877.320 351.940 877.580 352.200 ;
        RECT 877.780 351.260 878.040 351.520 ;
        RECT 876.860 303.320 877.120 303.580 ;
        RECT 877.780 303.320 878.040 303.580 ;
        RECT 877.780 255.380 878.040 255.640 ;
        RECT 876.860 255.040 877.120 255.300 ;
        RECT 662.040 134.340 662.300 134.600 ;
        RECT 877.320 134.340 877.580 134.600 ;
        RECT 656.980 16.700 657.240 16.960 ;
        RECT 662.040 16.700 662.300 16.960 ;
      LAYER met2 ;
        RECT 881.130 511.090 881.410 514.000 ;
        RECT 877.840 510.950 881.410 511.090 ;
        RECT 877.840 449.130 877.980 510.950 ;
        RECT 881.130 510.000 881.410 510.950 ;
        RECT 877.780 448.810 878.040 449.130 ;
        RECT 877.320 448.470 877.580 448.790 ;
        RECT 877.380 352.230 877.520 448.470 ;
        RECT 877.320 351.910 877.580 352.230 ;
        RECT 877.780 351.230 878.040 351.550 ;
        RECT 877.840 303.690 877.980 351.230 ;
        RECT 876.920 303.610 877.980 303.690 ;
        RECT 876.860 303.550 878.040 303.610 ;
        RECT 876.860 303.290 877.120 303.550 ;
        RECT 877.780 303.290 878.040 303.550 ;
        RECT 877.840 255.670 877.980 303.290 ;
        RECT 877.780 255.350 878.040 255.670 ;
        RECT 876.860 255.010 877.120 255.330 ;
        RECT 876.920 241.245 877.060 255.010 ;
        RECT 876.850 240.875 877.130 241.245 ;
        RECT 877.310 240.195 877.590 240.565 ;
        RECT 877.380 134.630 877.520 240.195 ;
        RECT 662.040 134.310 662.300 134.630 ;
        RECT 877.320 134.310 877.580 134.630 ;
        RECT 662.100 16.990 662.240 134.310 ;
        RECT 656.980 16.670 657.240 16.990 ;
        RECT 662.040 16.670 662.300 16.990 ;
        RECT 657.040 2.400 657.180 16.670 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 876.850 240.920 877.130 241.200 ;
        RECT 877.310 240.240 877.590 240.520 ;
      LAYER met3 ;
        RECT 876.825 241.210 877.155 241.225 ;
        RECT 876.150 240.910 877.155 241.210 ;
        RECT 876.150 240.530 876.450 240.910 ;
        RECT 876.825 240.895 877.155 240.910 ;
        RECT 877.285 240.530 877.615 240.545 ;
        RECT 876.150 240.230 877.615 240.530 ;
        RECT 877.285 240.215 877.615 240.230 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1117.945 186.405 1118.115 193.715 ;
      LAYER mcon ;
        RECT 1117.945 193.545 1118.115 193.715 ;
      LAYER met1 ;
        RECT 1118.330 392.940 1118.650 393.000 ;
        RECT 1120.630 392.940 1120.950 393.000 ;
        RECT 1118.330 392.800 1120.950 392.940 ;
        RECT 1118.330 392.740 1118.650 392.800 ;
        RECT 1120.630 392.740 1120.950 392.800 ;
        RECT 1118.330 255.720 1118.650 255.980 ;
        RECT 1118.420 255.300 1118.560 255.720 ;
        RECT 1118.330 255.040 1118.650 255.300 ;
        RECT 1117.885 193.700 1118.175 193.745 ;
        RECT 1118.330 193.700 1118.650 193.760 ;
        RECT 1117.885 193.560 1118.650 193.700 ;
        RECT 1117.885 193.515 1118.175 193.560 ;
        RECT 1118.330 193.500 1118.650 193.560 ;
        RECT 1117.870 186.560 1118.190 186.620 ;
        RECT 1117.675 186.420 1118.190 186.560 ;
        RECT 1117.870 186.360 1118.190 186.420 ;
        RECT 1000.110 113.800 1000.430 113.860 ;
        RECT 1117.870 113.800 1118.190 113.860 ;
        RECT 1000.110 113.660 1118.190 113.800 ;
        RECT 1000.110 113.600 1000.430 113.660 ;
        RECT 1117.870 113.600 1118.190 113.660 ;
        RECT 995.970 16.900 996.290 16.960 ;
        RECT 1000.110 16.900 1000.430 16.960 ;
        RECT 995.970 16.760 1000.430 16.900 ;
        RECT 995.970 16.700 996.290 16.760 ;
        RECT 1000.110 16.700 1000.430 16.760 ;
      LAYER via ;
        RECT 1118.360 392.740 1118.620 393.000 ;
        RECT 1120.660 392.740 1120.920 393.000 ;
        RECT 1118.360 255.720 1118.620 255.980 ;
        RECT 1118.360 255.040 1118.620 255.300 ;
        RECT 1118.360 193.500 1118.620 193.760 ;
        RECT 1117.900 186.360 1118.160 186.620 ;
        RECT 1000.140 113.600 1000.400 113.860 ;
        RECT 1117.900 113.600 1118.160 113.860 ;
        RECT 996.000 16.700 996.260 16.960 ;
        RECT 1000.140 16.700 1000.400 16.960 ;
      LAYER met2 ;
        RECT 1124.470 510.410 1124.750 514.000 ;
        RECT 1121.180 510.270 1124.750 510.410 ;
        RECT 1121.180 449.210 1121.320 510.270 ;
        RECT 1124.470 510.000 1124.750 510.270 ;
        RECT 1120.720 449.070 1121.320 449.210 ;
        RECT 1120.720 393.030 1120.860 449.070 ;
        RECT 1118.360 392.710 1118.620 393.030 ;
        RECT 1120.660 392.710 1120.920 393.030 ;
        RECT 1118.420 256.010 1118.560 392.710 ;
        RECT 1118.360 255.690 1118.620 256.010 ;
        RECT 1118.360 255.010 1118.620 255.330 ;
        RECT 1118.420 193.790 1118.560 255.010 ;
        RECT 1118.360 193.470 1118.620 193.790 ;
        RECT 1117.900 186.330 1118.160 186.650 ;
        RECT 1117.960 113.890 1118.100 186.330 ;
        RECT 1000.140 113.570 1000.400 113.890 ;
        RECT 1117.900 113.570 1118.160 113.890 ;
        RECT 1000.200 16.990 1000.340 113.570 ;
        RECT 996.000 16.670 996.260 16.990 ;
        RECT 1000.140 16.670 1000.400 16.990 ;
        RECT 996.060 2.400 996.200 16.670 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1132.665 379.525 1132.835 427.635 ;
        RECT 1133.125 241.485 1133.295 319.855 ;
        RECT 1133.125 144.925 1133.295 193.035 ;
      LAYER mcon ;
        RECT 1132.665 427.465 1132.835 427.635 ;
        RECT 1133.125 319.685 1133.295 319.855 ;
        RECT 1133.125 192.865 1133.295 193.035 ;
      LAYER met1 ;
        RECT 1132.590 427.620 1132.910 427.680 ;
        RECT 1132.395 427.480 1132.910 427.620 ;
        RECT 1132.590 427.420 1132.910 427.480 ;
        RECT 1132.605 379.680 1132.895 379.725 ;
        RECT 1133.050 379.680 1133.370 379.740 ;
        RECT 1132.605 379.540 1133.370 379.680 ;
        RECT 1132.605 379.495 1132.895 379.540 ;
        RECT 1133.050 379.480 1133.370 379.540 ;
        RECT 1133.050 338.540 1133.370 338.600 ;
        RECT 1132.680 338.400 1133.370 338.540 ;
        RECT 1132.680 337.920 1132.820 338.400 ;
        RECT 1133.050 338.340 1133.370 338.400 ;
        RECT 1132.590 337.660 1132.910 337.920 ;
        RECT 1132.590 319.840 1132.910 319.900 ;
        RECT 1133.065 319.840 1133.355 319.885 ;
        RECT 1132.590 319.700 1133.355 319.840 ;
        RECT 1132.590 319.640 1132.910 319.700 ;
        RECT 1133.065 319.655 1133.355 319.700 ;
        RECT 1133.050 241.640 1133.370 241.700 ;
        RECT 1132.855 241.500 1133.370 241.640 ;
        RECT 1133.050 241.440 1133.370 241.500 ;
        RECT 1133.050 193.020 1133.370 193.080 ;
        RECT 1132.855 192.880 1133.370 193.020 ;
        RECT 1133.050 192.820 1133.370 192.880 ;
        RECT 1133.050 145.080 1133.370 145.140 ;
        RECT 1132.855 144.940 1133.370 145.080 ;
        RECT 1133.050 144.880 1133.370 144.940 ;
        RECT 1013.450 120.600 1013.770 120.660 ;
        RECT 1133.050 120.600 1133.370 120.660 ;
        RECT 1013.450 120.460 1133.370 120.600 ;
        RECT 1013.450 120.400 1013.770 120.460 ;
        RECT 1133.050 120.400 1133.370 120.460 ;
      LAYER via ;
        RECT 1132.620 427.420 1132.880 427.680 ;
        RECT 1133.080 379.480 1133.340 379.740 ;
        RECT 1133.080 338.340 1133.340 338.600 ;
        RECT 1132.620 337.660 1132.880 337.920 ;
        RECT 1132.620 319.640 1132.880 319.900 ;
        RECT 1133.080 241.440 1133.340 241.700 ;
        RECT 1133.080 192.820 1133.340 193.080 ;
        RECT 1133.080 144.880 1133.340 145.140 ;
        RECT 1013.480 120.400 1013.740 120.660 ;
        RECT 1133.080 120.400 1133.340 120.660 ;
      LAYER met2 ;
        RECT 1137.350 510.410 1137.630 514.000 ;
        RECT 1134.980 510.270 1137.630 510.410 ;
        RECT 1134.980 435.045 1135.120 510.270 ;
        RECT 1137.350 510.000 1137.630 510.270 ;
        RECT 1132.610 434.675 1132.890 435.045 ;
        RECT 1134.910 434.675 1135.190 435.045 ;
        RECT 1132.680 427.710 1132.820 434.675 ;
        RECT 1132.620 427.390 1132.880 427.710 ;
        RECT 1133.080 379.450 1133.340 379.770 ;
        RECT 1133.140 338.630 1133.280 379.450 ;
        RECT 1133.080 338.310 1133.340 338.630 ;
        RECT 1132.620 337.630 1132.880 337.950 ;
        RECT 1132.680 319.930 1132.820 337.630 ;
        RECT 1132.620 319.610 1132.880 319.930 ;
        RECT 1133.080 241.410 1133.340 241.730 ;
        RECT 1133.140 193.110 1133.280 241.410 ;
        RECT 1133.080 192.790 1133.340 193.110 ;
        RECT 1133.080 144.850 1133.340 145.170 ;
        RECT 1133.140 120.690 1133.280 144.850 ;
        RECT 1013.480 120.370 1013.740 120.690 ;
        RECT 1133.080 120.370 1133.340 120.690 ;
        RECT 1013.540 2.400 1013.680 120.370 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 1132.610 434.720 1132.890 435.000 ;
        RECT 1134.910 434.720 1135.190 435.000 ;
      LAYER met3 ;
        RECT 1132.585 435.010 1132.915 435.025 ;
        RECT 1134.885 435.010 1135.215 435.025 ;
        RECT 1132.585 434.710 1135.215 435.010 ;
        RECT 1132.585 434.695 1132.915 434.710 ;
        RECT 1134.885 434.695 1135.215 434.710 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1146.925 241.485 1147.095 331.075 ;
        RECT 1146.925 144.925 1147.095 193.035 ;
        RECT 1146.925 106.845 1147.095 111.095 ;
      LAYER mcon ;
        RECT 1146.925 330.905 1147.095 331.075 ;
        RECT 1146.925 192.865 1147.095 193.035 ;
        RECT 1146.925 110.925 1147.095 111.095 ;
      LAYER met1 ;
        RECT 1146.390 427.960 1146.710 428.020 ;
        RECT 1148.230 427.960 1148.550 428.020 ;
        RECT 1146.390 427.820 1148.550 427.960 ;
        RECT 1146.390 427.760 1146.710 427.820 ;
        RECT 1148.230 427.760 1148.550 427.820 ;
        RECT 1146.390 331.060 1146.710 331.120 ;
        RECT 1146.865 331.060 1147.155 331.105 ;
        RECT 1146.390 330.920 1147.155 331.060 ;
        RECT 1146.390 330.860 1146.710 330.920 ;
        RECT 1146.865 330.875 1147.155 330.920 ;
        RECT 1146.850 241.640 1147.170 241.700 ;
        RECT 1146.655 241.500 1147.170 241.640 ;
        RECT 1146.850 241.440 1147.170 241.500 ;
        RECT 1146.850 193.020 1147.170 193.080 ;
        RECT 1146.655 192.880 1147.170 193.020 ;
        RECT 1146.850 192.820 1147.170 192.880 ;
        RECT 1146.850 145.080 1147.170 145.140 ;
        RECT 1146.655 144.940 1147.170 145.080 ;
        RECT 1146.850 144.880 1147.170 144.940 ;
        RECT 1146.850 111.080 1147.170 111.140 ;
        RECT 1146.655 110.940 1147.170 111.080 ;
        RECT 1146.850 110.880 1147.170 110.940 ;
        RECT 1034.610 107.000 1034.930 107.060 ;
        RECT 1146.865 107.000 1147.155 107.045 ;
        RECT 1034.610 106.860 1147.155 107.000 ;
        RECT 1034.610 106.800 1034.930 106.860 ;
        RECT 1146.865 106.815 1147.155 106.860 ;
        RECT 1031.390 5.680 1031.710 5.740 ;
        RECT 1034.610 5.680 1034.930 5.740 ;
        RECT 1031.390 5.540 1034.930 5.680 ;
        RECT 1031.390 5.480 1031.710 5.540 ;
        RECT 1034.610 5.480 1034.930 5.540 ;
      LAYER via ;
        RECT 1146.420 427.760 1146.680 428.020 ;
        RECT 1148.260 427.760 1148.520 428.020 ;
        RECT 1146.420 330.860 1146.680 331.120 ;
        RECT 1146.880 241.440 1147.140 241.700 ;
        RECT 1146.880 192.820 1147.140 193.080 ;
        RECT 1146.880 144.880 1147.140 145.140 ;
        RECT 1146.880 110.880 1147.140 111.140 ;
        RECT 1034.640 106.800 1034.900 107.060 ;
        RECT 1031.420 5.480 1031.680 5.740 ;
        RECT 1034.640 5.480 1034.900 5.740 ;
      LAYER met2 ;
        RECT 1150.230 510.410 1150.510 514.000 ;
        RECT 1148.320 510.270 1150.510 510.410 ;
        RECT 1148.320 428.050 1148.460 510.270 ;
        RECT 1150.230 510.000 1150.510 510.270 ;
        RECT 1146.420 427.730 1146.680 428.050 ;
        RECT 1148.260 427.730 1148.520 428.050 ;
        RECT 1146.480 379.285 1146.620 427.730 ;
        RECT 1145.030 378.915 1145.310 379.285 ;
        RECT 1146.410 378.915 1146.690 379.285 ;
        RECT 1145.100 331.685 1145.240 378.915 ;
        RECT 1145.030 331.315 1145.310 331.685 ;
        RECT 1146.410 331.315 1146.690 331.685 ;
        RECT 1146.480 331.150 1146.620 331.315 ;
        RECT 1146.420 330.830 1146.680 331.150 ;
        RECT 1146.880 241.410 1147.140 241.730 ;
        RECT 1146.940 193.110 1147.080 241.410 ;
        RECT 1146.880 192.790 1147.140 193.110 ;
        RECT 1146.880 144.850 1147.140 145.170 ;
        RECT 1146.940 111.170 1147.080 144.850 ;
        RECT 1146.880 110.850 1147.140 111.170 ;
        RECT 1034.640 106.770 1034.900 107.090 ;
        RECT 1034.700 5.770 1034.840 106.770 ;
        RECT 1031.420 5.450 1031.680 5.770 ;
        RECT 1034.640 5.450 1034.900 5.770 ;
        RECT 1031.480 2.400 1031.620 5.450 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 1145.030 378.960 1145.310 379.240 ;
        RECT 1146.410 378.960 1146.690 379.240 ;
        RECT 1145.030 331.360 1145.310 331.640 ;
        RECT 1146.410 331.360 1146.690 331.640 ;
      LAYER met3 ;
        RECT 1145.005 379.250 1145.335 379.265 ;
        RECT 1146.385 379.250 1146.715 379.265 ;
        RECT 1145.005 378.950 1146.715 379.250 ;
        RECT 1145.005 378.935 1145.335 378.950 ;
        RECT 1146.385 378.935 1146.715 378.950 ;
        RECT 1145.005 331.650 1145.335 331.665 ;
        RECT 1146.385 331.650 1146.715 331.665 ;
        RECT 1145.005 331.350 1146.715 331.650 ;
        RECT 1145.005 331.335 1145.335 331.350 ;
        RECT 1146.385 331.335 1146.715 331.350 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1055.310 79.460 1055.630 79.520 ;
        RECT 1159.270 79.460 1159.590 79.520 ;
        RECT 1055.310 79.320 1159.590 79.460 ;
        RECT 1055.310 79.260 1055.630 79.320 ;
        RECT 1159.270 79.260 1159.590 79.320 ;
        RECT 1049.330 17.240 1049.650 17.300 ;
        RECT 1055.310 17.240 1055.630 17.300 ;
        RECT 1049.330 17.100 1055.630 17.240 ;
        RECT 1049.330 17.040 1049.650 17.100 ;
        RECT 1055.310 17.040 1055.630 17.100 ;
      LAYER via ;
        RECT 1055.340 79.260 1055.600 79.520 ;
        RECT 1159.300 79.260 1159.560 79.520 ;
        RECT 1049.360 17.040 1049.620 17.300 ;
        RECT 1055.340 17.040 1055.600 17.300 ;
      LAYER met2 ;
        RECT 1163.110 510.410 1163.390 514.000 ;
        RECT 1159.360 510.270 1163.390 510.410 ;
        RECT 1159.360 79.550 1159.500 510.270 ;
        RECT 1163.110 510.000 1163.390 510.270 ;
        RECT 1055.340 79.230 1055.600 79.550 ;
        RECT 1159.300 79.230 1159.560 79.550 ;
        RECT 1055.400 17.330 1055.540 79.230 ;
        RECT 1049.360 17.010 1049.620 17.330 ;
        RECT 1055.340 17.010 1055.600 17.330 ;
        RECT 1049.420 2.400 1049.560 17.010 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1067.345 48.365 1067.515 86.275 ;
      LAYER mcon ;
        RECT 1067.345 86.105 1067.515 86.275 ;
      LAYER met1 ;
        RECT 1067.285 86.260 1067.575 86.305 ;
        RECT 1173.070 86.260 1173.390 86.320 ;
        RECT 1067.285 86.120 1173.390 86.260 ;
        RECT 1067.285 86.075 1067.575 86.120 ;
        RECT 1173.070 86.060 1173.390 86.120 ;
        RECT 1067.270 48.520 1067.590 48.580 ;
        RECT 1067.075 48.380 1067.590 48.520 ;
        RECT 1067.270 48.320 1067.590 48.380 ;
      LAYER via ;
        RECT 1173.100 86.060 1173.360 86.320 ;
        RECT 1067.300 48.320 1067.560 48.580 ;
      LAYER met2 ;
        RECT 1175.530 510.410 1175.810 514.000 ;
        RECT 1173.160 510.270 1175.810 510.410 ;
        RECT 1173.160 86.350 1173.300 510.270 ;
        RECT 1175.530 510.000 1175.810 510.270 ;
        RECT 1173.100 86.030 1173.360 86.350 ;
        RECT 1067.300 48.290 1067.560 48.610 ;
        RECT 1067.360 2.400 1067.500 48.290 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 93.060 1090.130 93.120 ;
        RECT 1187.330 93.060 1187.650 93.120 ;
        RECT 1089.810 92.920 1187.650 93.060 ;
        RECT 1089.810 92.860 1090.130 92.920 ;
        RECT 1187.330 92.860 1187.650 92.920 ;
        RECT 1085.210 16.900 1085.530 16.960 ;
        RECT 1089.810 16.900 1090.130 16.960 ;
        RECT 1085.210 16.760 1090.130 16.900 ;
        RECT 1085.210 16.700 1085.530 16.760 ;
        RECT 1089.810 16.700 1090.130 16.760 ;
      LAYER via ;
        RECT 1089.840 92.860 1090.100 93.120 ;
        RECT 1187.360 92.860 1187.620 93.120 ;
        RECT 1085.240 16.700 1085.500 16.960 ;
        RECT 1089.840 16.700 1090.100 16.960 ;
      LAYER met2 ;
        RECT 1188.410 510.410 1188.690 514.000 ;
        RECT 1187.420 510.270 1188.690 510.410 ;
        RECT 1187.420 93.150 1187.560 510.270 ;
        RECT 1188.410 510.000 1188.690 510.270 ;
        RECT 1089.840 92.830 1090.100 93.150 ;
        RECT 1187.360 92.830 1187.620 93.150 ;
        RECT 1089.900 16.990 1090.040 92.830 ;
        RECT 1085.240 16.670 1085.500 16.990 ;
        RECT 1089.840 16.670 1090.100 16.990 ;
        RECT 1085.300 2.400 1085.440 16.670 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1102.765 48.365 1102.935 72.335 ;
      LAYER mcon ;
        RECT 1102.765 72.165 1102.935 72.335 ;
      LAYER met1 ;
        RECT 1102.705 72.320 1102.995 72.365 ;
        RECT 1201.130 72.320 1201.450 72.380 ;
        RECT 1102.705 72.180 1201.450 72.320 ;
        RECT 1102.705 72.135 1102.995 72.180 ;
        RECT 1201.130 72.120 1201.450 72.180 ;
        RECT 1102.690 48.520 1103.010 48.580 ;
        RECT 1102.495 48.380 1103.010 48.520 ;
        RECT 1102.690 48.320 1103.010 48.380 ;
      LAYER via ;
        RECT 1201.160 72.120 1201.420 72.380 ;
        RECT 1102.720 48.320 1102.980 48.580 ;
      LAYER met2 ;
        RECT 1201.290 510.340 1201.570 514.000 ;
        RECT 1201.220 510.000 1201.570 510.340 ;
        RECT 1201.220 72.410 1201.360 510.000 ;
        RECT 1201.160 72.090 1201.420 72.410 ;
        RECT 1102.720 48.290 1102.980 48.610 ;
        RECT 1102.780 2.400 1102.920 48.290 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1208.030 421.160 1208.350 421.220 ;
        RECT 1208.950 421.160 1209.270 421.220 ;
        RECT 1208.030 421.020 1209.270 421.160 ;
        RECT 1208.030 420.960 1208.350 421.020 ;
        RECT 1208.950 420.960 1209.270 421.020 ;
        RECT 1208.490 241.640 1208.810 241.700 ;
        RECT 1208.950 241.640 1209.270 241.700 ;
        RECT 1208.490 241.500 1209.270 241.640 ;
        RECT 1208.490 241.440 1208.810 241.500 ;
        RECT 1208.950 241.440 1209.270 241.500 ;
        RECT 1120.630 16.900 1120.950 16.960 ;
        RECT 1208.030 16.900 1208.350 16.960 ;
        RECT 1120.630 16.760 1208.350 16.900 ;
        RECT 1120.630 16.700 1120.950 16.760 ;
        RECT 1208.030 16.700 1208.350 16.760 ;
      LAYER via ;
        RECT 1208.060 420.960 1208.320 421.220 ;
        RECT 1208.980 420.960 1209.240 421.220 ;
        RECT 1208.520 241.440 1208.780 241.700 ;
        RECT 1208.980 241.440 1209.240 241.700 ;
        RECT 1120.660 16.700 1120.920 16.960 ;
        RECT 1208.060 16.700 1208.320 16.960 ;
      LAYER met2 ;
        RECT 1214.170 510.410 1214.450 514.000 ;
        RECT 1212.260 510.270 1214.450 510.410 ;
        RECT 1212.260 472.330 1212.400 510.270 ;
        RECT 1214.170 510.000 1214.450 510.270 ;
        RECT 1209.040 472.190 1212.400 472.330 ;
        RECT 1209.040 421.250 1209.180 472.190 ;
        RECT 1208.060 420.930 1208.320 421.250 ;
        RECT 1208.980 420.930 1209.240 421.250 ;
        RECT 1208.120 400.250 1208.260 420.930 ;
        RECT 1208.120 400.110 1208.720 400.250 ;
        RECT 1208.580 351.970 1208.720 400.110 ;
        RECT 1208.580 351.830 1209.180 351.970 ;
        RECT 1209.040 241.730 1209.180 351.830 ;
        RECT 1208.520 241.410 1208.780 241.730 ;
        RECT 1208.980 241.410 1209.240 241.730 ;
        RECT 1208.580 207.130 1208.720 241.410 ;
        RECT 1208.580 206.990 1209.180 207.130 ;
        RECT 1209.040 158.850 1209.180 206.990 ;
        RECT 1208.120 158.710 1209.180 158.850 ;
        RECT 1208.120 158.170 1208.260 158.710 ;
        RECT 1208.120 158.030 1208.720 158.170 ;
        RECT 1208.580 62.290 1208.720 158.030 ;
        RECT 1208.120 62.150 1208.720 62.290 ;
        RECT 1208.120 16.990 1208.260 62.150 ;
        RECT 1120.660 16.670 1120.920 16.990 ;
        RECT 1208.060 16.670 1208.320 16.990 ;
        RECT 1120.720 2.400 1120.860 16.670 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1221.370 461.960 1221.690 462.020 ;
        RECT 1225.510 461.960 1225.830 462.020 ;
        RECT 1221.370 461.820 1225.830 461.960 ;
        RECT 1221.370 461.760 1221.690 461.820 ;
        RECT 1225.510 461.760 1225.830 461.820 ;
        RECT 1139.030 20.300 1139.350 20.360 ;
        RECT 1221.370 20.300 1221.690 20.360 ;
        RECT 1139.030 20.160 1221.690 20.300 ;
        RECT 1139.030 20.100 1139.350 20.160 ;
        RECT 1221.370 20.100 1221.690 20.160 ;
      LAYER via ;
        RECT 1221.400 461.760 1221.660 462.020 ;
        RECT 1225.540 461.760 1225.800 462.020 ;
        RECT 1139.060 20.100 1139.320 20.360 ;
        RECT 1221.400 20.100 1221.660 20.360 ;
      LAYER met2 ;
        RECT 1227.050 510.410 1227.330 514.000 ;
        RECT 1225.600 510.270 1227.330 510.410 ;
        RECT 1225.600 462.050 1225.740 510.270 ;
        RECT 1227.050 510.000 1227.330 510.270 ;
        RECT 1221.400 461.730 1221.660 462.050 ;
        RECT 1225.540 461.730 1225.800 462.050 ;
        RECT 1221.460 20.390 1221.600 461.730 ;
        RECT 1139.060 20.070 1139.320 20.390 ;
        RECT 1221.400 20.070 1221.660 20.390 ;
        RECT 1139.120 10.610 1139.260 20.070 ;
        RECT 1138.660 10.470 1139.260 10.610 ;
        RECT 1138.660 2.400 1138.800 10.470 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1235.170 472.840 1235.490 472.900 ;
        RECT 1238.390 472.840 1238.710 472.900 ;
        RECT 1235.170 472.700 1238.710 472.840 ;
        RECT 1235.170 472.640 1235.490 472.700 ;
        RECT 1238.390 472.640 1238.710 472.700 ;
        RECT 1156.510 19.960 1156.830 20.020 ;
        RECT 1235.170 19.960 1235.490 20.020 ;
        RECT 1156.510 19.820 1235.490 19.960 ;
        RECT 1156.510 19.760 1156.830 19.820 ;
        RECT 1235.170 19.760 1235.490 19.820 ;
      LAYER via ;
        RECT 1235.200 472.640 1235.460 472.900 ;
        RECT 1238.420 472.640 1238.680 472.900 ;
        RECT 1156.540 19.760 1156.800 20.020 ;
        RECT 1235.200 19.760 1235.460 20.020 ;
      LAYER met2 ;
        RECT 1239.930 510.410 1240.210 514.000 ;
        RECT 1238.480 510.270 1240.210 510.410 ;
        RECT 1238.480 472.930 1238.620 510.270 ;
        RECT 1239.930 510.000 1240.210 510.270 ;
        RECT 1235.200 472.610 1235.460 472.930 ;
        RECT 1238.420 472.610 1238.680 472.930 ;
        RECT 1235.260 20.050 1235.400 472.610 ;
        RECT 1156.540 19.730 1156.800 20.050 ;
        RECT 1235.200 19.730 1235.460 20.050 ;
        RECT 1156.600 2.400 1156.740 19.730 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 890.705 435.285 890.875 483.055 ;
        RECT 890.705 379.525 890.875 427.635 ;
        RECT 892.085 282.965 892.255 331.075 ;
      LAYER mcon ;
        RECT 890.705 482.885 890.875 483.055 ;
        RECT 890.705 427.465 890.875 427.635 ;
        RECT 892.085 330.905 892.255 331.075 ;
      LAYER met1 ;
        RECT 890.645 483.040 890.935 483.085 ;
        RECT 892.010 483.040 892.330 483.100 ;
        RECT 890.645 482.900 892.330 483.040 ;
        RECT 890.645 482.855 890.935 482.900 ;
        RECT 892.010 482.840 892.330 482.900 ;
        RECT 890.630 435.440 890.950 435.500 ;
        RECT 890.435 435.300 890.950 435.440 ;
        RECT 890.630 435.240 890.950 435.300 ;
        RECT 890.630 427.620 890.950 427.680 ;
        RECT 890.435 427.480 890.950 427.620 ;
        RECT 890.630 427.420 890.950 427.480 ;
        RECT 890.645 379.680 890.935 379.725 ;
        RECT 892.010 379.680 892.330 379.740 ;
        RECT 890.645 379.540 892.330 379.680 ;
        RECT 890.645 379.495 890.935 379.540 ;
        RECT 892.010 379.480 892.330 379.540 ;
        RECT 890.630 338.540 890.950 338.600 ;
        RECT 892.010 338.540 892.330 338.600 ;
        RECT 890.630 338.400 892.330 338.540 ;
        RECT 890.630 338.340 890.950 338.400 ;
        RECT 892.010 338.340 892.330 338.400 ;
        RECT 890.630 331.060 890.950 331.120 ;
        RECT 892.025 331.060 892.315 331.105 ;
        RECT 890.630 330.920 892.315 331.060 ;
        RECT 890.630 330.860 890.950 330.920 ;
        RECT 892.025 330.875 892.315 330.920 ;
        RECT 892.010 283.120 892.330 283.180 ;
        RECT 892.010 282.980 892.525 283.120 ;
        RECT 892.010 282.920 892.330 282.980 ;
        RECT 890.630 241.640 890.950 241.700 ;
        RECT 892.010 241.640 892.330 241.700 ;
        RECT 890.630 241.500 892.330 241.640 ;
        RECT 890.630 241.440 890.950 241.500 ;
        RECT 892.010 241.440 892.330 241.500 ;
        RECT 891.090 193.840 891.410 194.100 ;
        RECT 891.180 193.420 891.320 193.840 ;
        RECT 891.090 193.160 891.410 193.420 ;
        RECT 674.430 37.980 674.750 38.040 ;
        RECT 891.090 37.980 891.410 38.040 ;
        RECT 674.430 37.840 891.410 37.980 ;
        RECT 674.430 37.780 674.750 37.840 ;
        RECT 891.090 37.780 891.410 37.840 ;
      LAYER via ;
        RECT 892.040 482.840 892.300 483.100 ;
        RECT 890.660 435.240 890.920 435.500 ;
        RECT 890.660 427.420 890.920 427.680 ;
        RECT 892.040 379.480 892.300 379.740 ;
        RECT 890.660 338.340 890.920 338.600 ;
        RECT 892.040 338.340 892.300 338.600 ;
        RECT 890.660 330.860 890.920 331.120 ;
        RECT 892.040 282.920 892.300 283.180 ;
        RECT 890.660 241.440 890.920 241.700 ;
        RECT 892.040 241.440 892.300 241.700 ;
        RECT 891.120 193.840 891.380 194.100 ;
        RECT 891.120 193.160 891.380 193.420 ;
        RECT 674.460 37.780 674.720 38.040 ;
        RECT 891.120 37.780 891.380 38.040 ;
      LAYER met2 ;
        RECT 894.010 510.410 894.290 514.000 ;
        RECT 892.100 510.270 894.290 510.410 ;
        RECT 892.100 483.130 892.240 510.270 ;
        RECT 894.010 510.000 894.290 510.270 ;
        RECT 892.040 482.810 892.300 483.130 ;
        RECT 890.660 435.210 890.920 435.530 ;
        RECT 890.720 427.710 890.860 435.210 ;
        RECT 890.660 427.390 890.920 427.710 ;
        RECT 892.040 379.450 892.300 379.770 ;
        RECT 892.100 338.630 892.240 379.450 ;
        RECT 890.660 338.310 890.920 338.630 ;
        RECT 892.040 338.310 892.300 338.630 ;
        RECT 890.720 331.150 890.860 338.310 ;
        RECT 890.660 330.830 890.920 331.150 ;
        RECT 892.040 282.890 892.300 283.210 ;
        RECT 892.100 241.730 892.240 282.890 ;
        RECT 890.660 241.410 890.920 241.730 ;
        RECT 892.040 241.410 892.300 241.730 ;
        RECT 890.720 224.810 890.860 241.410 ;
        RECT 890.720 224.670 891.320 224.810 ;
        RECT 891.180 194.130 891.320 224.670 ;
        RECT 891.120 193.810 891.380 194.130 ;
        RECT 891.120 193.130 891.380 193.450 ;
        RECT 891.180 169.050 891.320 193.130 ;
        RECT 890.720 168.910 891.320 169.050 ;
        RECT 890.720 158.170 890.860 168.910 ;
        RECT 890.720 158.030 891.780 158.170 ;
        RECT 891.640 110.570 891.780 158.030 ;
        RECT 890.720 110.430 891.780 110.570 ;
        RECT 890.720 109.890 890.860 110.430 ;
        RECT 890.720 109.750 891.320 109.890 ;
        RECT 891.180 38.070 891.320 109.750 ;
        RECT 674.460 37.750 674.720 38.070 ;
        RECT 891.120 37.750 891.380 38.070 ;
        RECT 674.520 2.400 674.660 37.750 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 17.240 1174.310 17.300 ;
        RECT 1248.970 17.240 1249.290 17.300 ;
        RECT 1173.990 17.100 1249.290 17.240 ;
        RECT 1173.990 17.040 1174.310 17.100 ;
        RECT 1248.970 17.040 1249.290 17.100 ;
      LAYER via ;
        RECT 1174.020 17.040 1174.280 17.300 ;
        RECT 1249.000 17.040 1249.260 17.300 ;
      LAYER met2 ;
        RECT 1252.350 510.410 1252.630 514.000 ;
        RECT 1249.060 510.270 1252.630 510.410 ;
        RECT 1249.060 17.330 1249.200 510.270 ;
        RECT 1252.350 510.000 1252.630 510.270 ;
        RECT 1174.020 17.010 1174.280 17.330 ;
        RECT 1249.000 17.010 1249.260 17.330 ;
        RECT 1174.080 2.400 1174.220 17.010 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.770 241.780 1263.090 242.040 ;
        RECT 1262.860 241.020 1263.000 241.780 ;
        RECT 1262.770 240.760 1263.090 241.020 ;
        RECT 1191.930 17.580 1192.250 17.640 ;
        RECT 1262.770 17.580 1263.090 17.640 ;
        RECT 1191.930 17.440 1263.090 17.580 ;
        RECT 1191.930 17.380 1192.250 17.440 ;
        RECT 1262.770 17.380 1263.090 17.440 ;
      LAYER via ;
        RECT 1262.800 241.780 1263.060 242.040 ;
        RECT 1262.800 240.760 1263.060 241.020 ;
        RECT 1191.960 17.380 1192.220 17.640 ;
        RECT 1262.800 17.380 1263.060 17.640 ;
      LAYER met2 ;
        RECT 1265.230 510.410 1265.510 514.000 ;
        RECT 1262.860 510.270 1265.510 510.410 ;
        RECT 1262.860 242.070 1263.000 510.270 ;
        RECT 1265.230 510.000 1265.510 510.270 ;
        RECT 1262.800 241.750 1263.060 242.070 ;
        RECT 1262.800 240.730 1263.060 241.050 ;
        RECT 1262.860 17.670 1263.000 240.730 ;
        RECT 1191.960 17.350 1192.220 17.670 ;
        RECT 1262.800 17.350 1263.060 17.670 ;
        RECT 1192.020 2.400 1192.160 17.350 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1209.870 18.940 1210.190 19.000 ;
        RECT 1276.570 18.940 1276.890 19.000 ;
        RECT 1209.870 18.800 1276.890 18.940 ;
        RECT 1209.870 18.740 1210.190 18.800 ;
        RECT 1276.570 18.740 1276.890 18.800 ;
      LAYER via ;
        RECT 1209.900 18.740 1210.160 19.000 ;
        RECT 1276.600 18.740 1276.860 19.000 ;
      LAYER met2 ;
        RECT 1278.110 510.410 1278.390 514.000 ;
        RECT 1276.660 510.270 1278.390 510.410 ;
        RECT 1276.660 19.030 1276.800 510.270 ;
        RECT 1278.110 510.000 1278.390 510.270 ;
        RECT 1209.900 18.710 1210.160 19.030 ;
        RECT 1276.600 18.710 1276.860 19.030 ;
        RECT 1209.960 2.400 1210.100 18.710 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 18.260 1228.130 18.320 ;
        RECT 1290.370 18.260 1290.690 18.320 ;
        RECT 1227.810 18.120 1290.690 18.260 ;
        RECT 1227.810 18.060 1228.130 18.120 ;
        RECT 1290.370 18.060 1290.690 18.120 ;
      LAYER via ;
        RECT 1227.840 18.060 1228.100 18.320 ;
        RECT 1290.400 18.060 1290.660 18.320 ;
      LAYER met2 ;
        RECT 1290.990 510.410 1291.270 514.000 ;
        RECT 1290.460 510.270 1291.270 510.410 ;
        RECT 1290.460 18.350 1290.600 510.270 ;
        RECT 1290.990 510.000 1291.270 510.270 ;
        RECT 1227.840 18.030 1228.100 18.350 ;
        RECT 1290.400 18.030 1290.660 18.350 ;
        RECT 1227.900 2.400 1228.040 18.030 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1297.270 456.520 1297.590 456.580 ;
        RECT 1301.870 456.520 1302.190 456.580 ;
        RECT 1297.270 456.380 1302.190 456.520 ;
        RECT 1297.270 456.320 1297.590 456.380 ;
        RECT 1301.870 456.320 1302.190 456.380 ;
        RECT 1245.750 20.300 1246.070 20.360 ;
        RECT 1297.270 20.300 1297.590 20.360 ;
        RECT 1245.750 20.160 1297.590 20.300 ;
        RECT 1245.750 20.100 1246.070 20.160 ;
        RECT 1297.270 20.100 1297.590 20.160 ;
      LAYER via ;
        RECT 1297.300 456.320 1297.560 456.580 ;
        RECT 1301.900 456.320 1302.160 456.580 ;
        RECT 1245.780 20.100 1246.040 20.360 ;
        RECT 1297.300 20.100 1297.560 20.360 ;
      LAYER met2 ;
        RECT 1303.870 510.410 1304.150 514.000 ;
        RECT 1301.960 510.270 1304.150 510.410 ;
        RECT 1301.960 456.610 1302.100 510.270 ;
        RECT 1303.870 510.000 1304.150 510.270 ;
        RECT 1297.300 456.290 1297.560 456.610 ;
        RECT 1301.900 456.290 1302.160 456.610 ;
        RECT 1297.360 20.390 1297.500 456.290 ;
        RECT 1245.780 20.070 1246.040 20.390 ;
        RECT 1297.300 20.070 1297.560 20.390 ;
        RECT 1245.840 2.400 1245.980 20.070 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1311.070 461.960 1311.390 462.020 ;
        RECT 1314.750 461.960 1315.070 462.020 ;
        RECT 1311.070 461.820 1315.070 461.960 ;
        RECT 1311.070 461.760 1311.390 461.820 ;
        RECT 1314.750 461.760 1315.070 461.820 ;
        RECT 1263.690 20.640 1264.010 20.700 ;
        RECT 1311.070 20.640 1311.390 20.700 ;
        RECT 1263.690 20.500 1311.390 20.640 ;
        RECT 1263.690 20.440 1264.010 20.500 ;
        RECT 1311.070 20.440 1311.390 20.500 ;
      LAYER via ;
        RECT 1311.100 461.760 1311.360 462.020 ;
        RECT 1314.780 461.760 1315.040 462.020 ;
        RECT 1263.720 20.440 1263.980 20.700 ;
        RECT 1311.100 20.440 1311.360 20.700 ;
      LAYER met2 ;
        RECT 1316.750 510.410 1317.030 514.000 ;
        RECT 1314.840 510.270 1317.030 510.410 ;
        RECT 1314.840 462.050 1314.980 510.270 ;
        RECT 1316.750 510.000 1317.030 510.270 ;
        RECT 1311.100 461.730 1311.360 462.050 ;
        RECT 1314.780 461.730 1315.040 462.050 ;
        RECT 1311.160 20.730 1311.300 461.730 ;
        RECT 1263.720 20.410 1263.980 20.730 ;
        RECT 1311.100 20.410 1311.360 20.730 ;
        RECT 1263.780 10.610 1263.920 20.410 ;
        RECT 1263.320 10.470 1263.920 10.610 ;
        RECT 1263.320 2.400 1263.460 10.470 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1324.870 472.840 1325.190 472.900 ;
        RECT 1327.630 472.840 1327.950 472.900 ;
        RECT 1324.870 472.700 1327.950 472.840 ;
        RECT 1324.870 472.640 1325.190 472.700 ;
        RECT 1327.630 472.640 1327.950 472.700 ;
        RECT 1281.170 18.940 1281.490 19.000 ;
        RECT 1324.870 18.940 1325.190 19.000 ;
        RECT 1281.170 18.800 1325.190 18.940 ;
        RECT 1281.170 18.740 1281.490 18.800 ;
        RECT 1324.870 18.740 1325.190 18.800 ;
      LAYER via ;
        RECT 1324.900 472.640 1325.160 472.900 ;
        RECT 1327.660 472.640 1327.920 472.900 ;
        RECT 1281.200 18.740 1281.460 19.000 ;
        RECT 1324.900 18.740 1325.160 19.000 ;
      LAYER met2 ;
        RECT 1329.170 510.410 1329.450 514.000 ;
        RECT 1327.720 510.270 1329.450 510.410 ;
        RECT 1327.720 472.930 1327.860 510.270 ;
        RECT 1329.170 510.000 1329.450 510.270 ;
        RECT 1324.900 472.610 1325.160 472.930 ;
        RECT 1327.660 472.610 1327.920 472.930 ;
        RECT 1324.960 19.030 1325.100 472.610 ;
        RECT 1281.200 18.710 1281.460 19.030 ;
        RECT 1324.900 18.710 1325.160 19.030 ;
        RECT 1281.260 2.400 1281.400 18.710 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 19.620 1299.430 19.680 ;
        RECT 1338.670 19.620 1338.990 19.680 ;
        RECT 1299.110 19.480 1338.990 19.620 ;
        RECT 1299.110 19.420 1299.430 19.480 ;
        RECT 1338.670 19.420 1338.990 19.480 ;
      LAYER via ;
        RECT 1299.140 19.420 1299.400 19.680 ;
        RECT 1338.700 19.420 1338.960 19.680 ;
      LAYER met2 ;
        RECT 1342.050 510.410 1342.330 514.000 ;
        RECT 1338.760 510.270 1342.330 510.410 ;
        RECT 1338.760 19.710 1338.900 510.270 ;
        RECT 1342.050 510.000 1342.330 510.270 ;
        RECT 1299.140 19.390 1299.400 19.710 ;
        RECT 1338.700 19.390 1338.960 19.710 ;
        RECT 1299.200 2.400 1299.340 19.390 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1317.050 17.780 1322.800 17.920 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
        RECT 1322.660 17.580 1322.800 17.780 ;
        RECT 1352.930 17.580 1353.250 17.640 ;
        RECT 1322.660 17.440 1353.250 17.580 ;
        RECT 1352.930 17.380 1353.250 17.440 ;
      LAYER via ;
        RECT 1317.080 17.720 1317.340 17.980 ;
        RECT 1352.960 17.380 1353.220 17.640 ;
      LAYER met2 ;
        RECT 1354.930 510.410 1355.210 514.000 ;
        RECT 1353.020 510.270 1355.210 510.410 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1317.140 2.400 1317.280 17.690 ;
        RECT 1353.020 17.670 1353.160 510.270 ;
        RECT 1354.930 510.000 1355.210 510.270 ;
        RECT 1352.960 17.350 1353.220 17.670 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 17.240 1335.310 17.300 ;
        RECT 1366.730 17.240 1367.050 17.300 ;
        RECT 1334.990 17.100 1367.050 17.240 ;
        RECT 1334.990 17.040 1335.310 17.100 ;
        RECT 1366.730 17.040 1367.050 17.100 ;
      LAYER via ;
        RECT 1335.020 17.040 1335.280 17.300 ;
        RECT 1366.760 17.040 1367.020 17.300 ;
      LAYER met2 ;
        RECT 1367.810 510.410 1368.090 514.000 ;
        RECT 1366.820 510.270 1368.090 510.410 ;
        RECT 1366.820 17.330 1366.960 510.270 ;
        RECT 1367.810 510.000 1368.090 510.270 ;
        RECT 1335.020 17.010 1335.280 17.330 ;
        RECT 1366.760 17.010 1367.020 17.330 ;
        RECT 1335.080 2.400 1335.220 17.010 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.510 451.760 696.830 451.820 ;
        RECT 903.970 451.760 904.290 451.820 ;
        RECT 696.510 451.620 904.290 451.760 ;
        RECT 696.510 451.560 696.830 451.620 ;
        RECT 903.970 451.560 904.290 451.620 ;
        RECT 692.370 16.900 692.690 16.960 ;
        RECT 696.510 16.900 696.830 16.960 ;
        RECT 692.370 16.760 696.830 16.900 ;
        RECT 692.370 16.700 692.690 16.760 ;
        RECT 696.510 16.700 696.830 16.760 ;
      LAYER via ;
        RECT 696.540 451.560 696.800 451.820 ;
        RECT 904.000 451.560 904.260 451.820 ;
        RECT 692.400 16.700 692.660 16.960 ;
        RECT 696.540 16.700 696.800 16.960 ;
      LAYER met2 ;
        RECT 906.890 510.410 907.170 514.000 ;
        RECT 904.060 510.270 907.170 510.410 ;
        RECT 904.060 451.850 904.200 510.270 ;
        RECT 906.890 510.000 907.170 510.270 ;
        RECT 696.540 451.530 696.800 451.850 ;
        RECT 904.000 451.530 904.260 451.850 ;
        RECT 696.600 16.990 696.740 451.530 ;
        RECT 692.400 16.670 692.660 16.990 ;
        RECT 696.540 16.670 696.800 16.990 ;
        RECT 692.460 2.400 692.600 16.670 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 16.900 1352.790 16.960 ;
        RECT 1380.530 16.900 1380.850 16.960 ;
        RECT 1352.470 16.760 1380.850 16.900 ;
        RECT 1352.470 16.700 1352.790 16.760 ;
        RECT 1380.530 16.700 1380.850 16.760 ;
      LAYER via ;
        RECT 1352.500 16.700 1352.760 16.960 ;
        RECT 1380.560 16.700 1380.820 16.960 ;
      LAYER met2 ;
        RECT 1380.690 510.340 1380.970 514.000 ;
        RECT 1380.620 510.000 1380.970 510.340 ;
        RECT 1380.620 16.990 1380.760 510.000 ;
        RECT 1352.500 16.670 1352.760 16.990 ;
        RECT 1380.560 16.670 1380.820 16.990 ;
        RECT 1352.560 2.400 1352.700 16.670 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1387.890 386.480 1388.210 386.540 ;
        RECT 1388.350 386.480 1388.670 386.540 ;
        RECT 1387.890 386.340 1388.670 386.480 ;
        RECT 1387.890 386.280 1388.210 386.340 ;
        RECT 1388.350 386.280 1388.670 386.340 ;
        RECT 1387.890 352.140 1388.210 352.200 ;
        RECT 1387.520 352.000 1388.210 352.140 ;
        RECT 1387.520 351.860 1387.660 352.000 ;
        RECT 1387.890 351.940 1388.210 352.000 ;
        RECT 1387.430 351.600 1387.750 351.860 ;
        RECT 1387.430 304.540 1387.750 304.600 ;
        RECT 1387.430 304.400 1388.120 304.540 ;
        RECT 1387.430 304.340 1387.750 304.400 ;
        RECT 1387.980 303.580 1388.120 304.400 ;
        RECT 1387.890 303.320 1388.210 303.580 ;
        RECT 1370.410 15.200 1370.730 15.260 ;
        RECT 1387.890 15.200 1388.210 15.260 ;
        RECT 1370.410 15.060 1388.210 15.200 ;
        RECT 1370.410 15.000 1370.730 15.060 ;
        RECT 1387.890 15.000 1388.210 15.060 ;
      LAYER via ;
        RECT 1387.920 386.280 1388.180 386.540 ;
        RECT 1388.380 386.280 1388.640 386.540 ;
        RECT 1387.920 351.940 1388.180 352.200 ;
        RECT 1387.460 351.600 1387.720 351.860 ;
        RECT 1387.460 304.340 1387.720 304.600 ;
        RECT 1387.920 303.320 1388.180 303.580 ;
        RECT 1370.440 15.000 1370.700 15.260 ;
        RECT 1387.920 15.000 1388.180 15.260 ;
      LAYER met2 ;
        RECT 1393.570 511.090 1393.850 514.000 ;
        RECT 1389.820 510.950 1393.850 511.090 ;
        RECT 1389.820 449.210 1389.960 510.950 ;
        RECT 1393.570 510.000 1393.850 510.950 ;
        RECT 1388.440 449.070 1389.960 449.210 ;
        RECT 1388.440 386.570 1388.580 449.070 ;
        RECT 1387.920 386.250 1388.180 386.570 ;
        RECT 1388.380 386.250 1388.640 386.570 ;
        RECT 1387.980 352.230 1388.120 386.250 ;
        RECT 1387.920 351.910 1388.180 352.230 ;
        RECT 1387.460 351.570 1387.720 351.890 ;
        RECT 1387.520 304.630 1387.660 351.570 ;
        RECT 1387.460 304.310 1387.720 304.630 ;
        RECT 1387.920 303.290 1388.180 303.610 ;
        RECT 1387.980 207.130 1388.120 303.290 ;
        RECT 1387.520 206.990 1388.120 207.130 ;
        RECT 1387.520 206.450 1387.660 206.990 ;
        RECT 1387.520 206.310 1388.120 206.450 ;
        RECT 1387.980 110.570 1388.120 206.310 ;
        RECT 1387.520 110.430 1388.120 110.570 ;
        RECT 1387.520 109.890 1387.660 110.430 ;
        RECT 1387.520 109.750 1388.120 109.890 ;
        RECT 1387.980 15.290 1388.120 109.750 ;
        RECT 1370.440 14.970 1370.700 15.290 ;
        RECT 1387.920 14.970 1388.180 15.290 ;
        RECT 1370.500 2.400 1370.640 14.970 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1401.690 338.200 1402.010 338.260 ;
        RECT 1402.150 338.200 1402.470 338.260 ;
        RECT 1401.690 338.060 1402.470 338.200 ;
        RECT 1401.690 338.000 1402.010 338.060 ;
        RECT 1402.150 338.000 1402.470 338.060 ;
        RECT 1388.350 20.640 1388.670 20.700 ;
        RECT 1401.690 20.640 1402.010 20.700 ;
        RECT 1388.350 20.500 1402.010 20.640 ;
        RECT 1388.350 20.440 1388.670 20.500 ;
        RECT 1401.690 20.440 1402.010 20.500 ;
      LAYER via ;
        RECT 1401.720 338.000 1401.980 338.260 ;
        RECT 1402.180 338.000 1402.440 338.260 ;
        RECT 1388.380 20.440 1388.640 20.700 ;
        RECT 1401.720 20.440 1401.980 20.700 ;
      LAYER met2 ;
        RECT 1405.990 511.090 1406.270 514.000 ;
        RECT 1402.700 510.950 1406.270 511.090 ;
        RECT 1402.700 449.210 1402.840 510.950 ;
        RECT 1405.990 510.000 1406.270 510.950 ;
        RECT 1402.240 449.070 1402.840 449.210 ;
        RECT 1402.240 338.290 1402.380 449.070 ;
        RECT 1401.720 337.970 1401.980 338.290 ;
        RECT 1402.180 337.970 1402.440 338.290 ;
        RECT 1401.780 207.130 1401.920 337.970 ;
        RECT 1401.320 206.990 1401.920 207.130 ;
        RECT 1401.320 206.450 1401.460 206.990 ;
        RECT 1401.320 206.310 1401.920 206.450 ;
        RECT 1401.780 110.570 1401.920 206.310 ;
        RECT 1401.320 110.430 1401.920 110.570 ;
        RECT 1401.320 109.890 1401.460 110.430 ;
        RECT 1401.320 109.750 1401.920 109.890 ;
        RECT 1401.780 20.730 1401.920 109.750 ;
        RECT 1388.380 20.410 1388.640 20.730 ;
        RECT 1401.720 20.410 1401.980 20.730 ;
        RECT 1388.440 2.400 1388.580 20.410 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1415.565 289.765 1415.735 337.875 ;
      LAYER mcon ;
        RECT 1415.565 337.705 1415.735 337.875 ;
      LAYER met1 ;
        RECT 1415.490 337.860 1415.810 337.920 ;
        RECT 1415.295 337.720 1415.810 337.860 ;
        RECT 1415.490 337.660 1415.810 337.720 ;
        RECT 1415.490 289.920 1415.810 289.980 ;
        RECT 1415.295 289.780 1415.810 289.920 ;
        RECT 1415.490 289.720 1415.810 289.780 ;
        RECT 1406.290 15.200 1406.610 15.260 ;
        RECT 1415.490 15.200 1415.810 15.260 ;
        RECT 1406.290 15.060 1415.810 15.200 ;
        RECT 1406.290 15.000 1406.610 15.060 ;
        RECT 1415.490 15.000 1415.810 15.060 ;
      LAYER via ;
        RECT 1415.520 337.660 1415.780 337.920 ;
        RECT 1415.520 289.720 1415.780 289.980 ;
        RECT 1406.320 15.000 1406.580 15.260 ;
        RECT 1415.520 15.000 1415.780 15.260 ;
      LAYER met2 ;
        RECT 1418.870 510.410 1419.150 514.000 ;
        RECT 1416.960 510.270 1419.150 510.410 ;
        RECT 1416.960 449.210 1417.100 510.270 ;
        RECT 1418.870 510.000 1419.150 510.270 ;
        RECT 1416.040 449.070 1417.100 449.210 ;
        RECT 1416.040 351.290 1416.180 449.070 ;
        RECT 1415.580 351.150 1416.180 351.290 ;
        RECT 1415.580 337.950 1415.720 351.150 ;
        RECT 1415.520 337.630 1415.780 337.950 ;
        RECT 1415.520 289.690 1415.780 290.010 ;
        RECT 1415.580 207.130 1415.720 289.690 ;
        RECT 1415.120 206.990 1415.720 207.130 ;
        RECT 1415.120 206.450 1415.260 206.990 ;
        RECT 1415.120 206.310 1415.720 206.450 ;
        RECT 1415.580 110.570 1415.720 206.310 ;
        RECT 1415.120 110.430 1415.720 110.570 ;
        RECT 1415.120 109.890 1415.260 110.430 ;
        RECT 1415.120 109.750 1415.720 109.890 ;
        RECT 1415.580 15.290 1415.720 109.750 ;
        RECT 1406.320 14.970 1406.580 15.290 ;
        RECT 1415.520 14.970 1415.780 15.290 ;
        RECT 1406.380 2.400 1406.520 14.970 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.770 20.640 1424.090 20.700 ;
        RECT 1428.370 20.640 1428.690 20.700 ;
        RECT 1423.770 20.500 1428.690 20.640 ;
        RECT 1423.770 20.440 1424.090 20.500 ;
        RECT 1428.370 20.440 1428.690 20.500 ;
      LAYER via ;
        RECT 1423.800 20.440 1424.060 20.700 ;
        RECT 1428.400 20.440 1428.660 20.700 ;
      LAYER met2 ;
        RECT 1431.750 510.410 1432.030 514.000 ;
        RECT 1428.460 510.270 1432.030 510.410 ;
        RECT 1428.460 20.730 1428.600 510.270 ;
        RECT 1431.750 510.000 1432.030 510.270 ;
        RECT 1423.800 20.410 1424.060 20.730 ;
        RECT 1428.400 20.410 1428.660 20.730 ;
        RECT 1423.860 2.400 1424.000 20.410 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.630 510.410 1444.910 514.000 ;
        RECT 1442.260 510.270 1444.910 510.410 ;
        RECT 1442.260 20.300 1442.400 510.270 ;
        RECT 1444.630 510.000 1444.910 510.270 ;
        RECT 1441.800 20.160 1442.400 20.300 ;
        RECT 1441.800 2.400 1441.940 20.160 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1456.430 20.640 1456.750 20.700 ;
        RECT 1459.650 20.640 1459.970 20.700 ;
        RECT 1456.430 20.500 1459.970 20.640 ;
        RECT 1456.430 20.440 1456.750 20.500 ;
        RECT 1459.650 20.440 1459.970 20.500 ;
      LAYER via ;
        RECT 1456.460 20.440 1456.720 20.700 ;
        RECT 1459.680 20.440 1459.940 20.700 ;
      LAYER met2 ;
        RECT 1457.510 510.410 1457.790 514.000 ;
        RECT 1456.520 510.270 1457.790 510.410 ;
        RECT 1456.520 20.730 1456.660 510.270 ;
        RECT 1457.510 510.000 1457.790 510.270 ;
        RECT 1456.460 20.410 1456.720 20.730 ;
        RECT 1459.680 20.410 1459.940 20.730 ;
        RECT 1459.740 2.400 1459.880 20.410 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1470.230 496.980 1470.550 497.040 ;
        RECT 1475.750 496.980 1476.070 497.040 ;
        RECT 1470.230 496.840 1476.070 496.980 ;
        RECT 1470.230 496.780 1470.550 496.840 ;
        RECT 1475.750 496.780 1476.070 496.840 ;
      LAYER via ;
        RECT 1470.260 496.780 1470.520 497.040 ;
        RECT 1475.780 496.780 1476.040 497.040 ;
      LAYER met2 ;
        RECT 1470.390 510.340 1470.670 514.000 ;
        RECT 1470.320 510.000 1470.670 510.340 ;
        RECT 1470.320 497.070 1470.460 510.000 ;
        RECT 1470.260 496.750 1470.520 497.070 ;
        RECT 1475.780 496.750 1476.040 497.070 ;
        RECT 1475.840 17.410 1475.980 496.750 ;
        RECT 1475.840 17.270 1477.820 17.410 ;
        RECT 1477.680 2.400 1477.820 17.270 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1482.650 14.520 1482.970 14.580 ;
        RECT 1495.530 14.520 1495.850 14.580 ;
        RECT 1482.650 14.380 1495.850 14.520 ;
        RECT 1482.650 14.320 1482.970 14.380 ;
        RECT 1495.530 14.320 1495.850 14.380 ;
      LAYER via ;
        RECT 1482.680 14.320 1482.940 14.580 ;
        RECT 1495.560 14.320 1495.820 14.580 ;
      LAYER met2 ;
        RECT 1482.810 510.340 1483.090 514.000 ;
        RECT 1482.740 510.000 1483.090 510.340 ;
        RECT 1482.740 14.610 1482.880 510.000 ;
        RECT 1482.680 14.290 1482.940 14.610 ;
        RECT 1495.560 14.290 1495.820 14.610 ;
        RECT 1495.620 2.400 1495.760 14.290 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.450 16.900 1496.770 16.960 ;
        RECT 1513.010 16.900 1513.330 16.960 ;
        RECT 1496.450 16.760 1513.330 16.900 ;
        RECT 1496.450 16.700 1496.770 16.760 ;
        RECT 1513.010 16.700 1513.330 16.760 ;
      LAYER via ;
        RECT 1496.480 16.700 1496.740 16.960 ;
        RECT 1513.040 16.700 1513.300 16.960 ;
      LAYER met2 ;
        RECT 1495.690 510.410 1495.970 514.000 ;
        RECT 1495.690 510.270 1496.680 510.410 ;
        RECT 1495.690 510.000 1495.970 510.270 ;
        RECT 1496.540 16.990 1496.680 510.270 ;
        RECT 1496.480 16.670 1496.740 16.990 ;
        RECT 1513.040 16.670 1513.300 16.990 ;
        RECT 1513.100 2.400 1513.240 16.670 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 893.390 500.040 893.710 500.100 ;
        RECT 919.610 500.040 919.930 500.100 ;
        RECT 893.390 499.900 919.930 500.040 ;
        RECT 893.390 499.840 893.710 499.900 ;
        RECT 919.610 499.840 919.930 499.900 ;
        RECT 710.310 141.340 710.630 141.400 ;
        RECT 893.390 141.340 893.710 141.400 ;
        RECT 710.310 141.200 893.710 141.340 ;
        RECT 710.310 141.140 710.630 141.200 ;
        RECT 893.390 141.140 893.710 141.200 ;
      LAYER via ;
        RECT 893.420 499.840 893.680 500.100 ;
        RECT 919.640 499.840 919.900 500.100 ;
        RECT 710.340 141.140 710.600 141.400 ;
        RECT 893.420 141.140 893.680 141.400 ;
      LAYER met2 ;
        RECT 919.770 510.340 920.050 514.000 ;
        RECT 919.700 510.000 920.050 510.340 ;
        RECT 919.700 500.130 919.840 510.000 ;
        RECT 893.420 499.810 893.680 500.130 ;
        RECT 919.640 499.810 919.900 500.130 ;
        RECT 893.480 141.430 893.620 499.810 ;
        RECT 710.340 141.110 710.600 141.430 ;
        RECT 893.420 141.110 893.680 141.430 ;
        RECT 710.400 2.400 710.540 141.110 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.250 16.560 1510.570 16.620 ;
        RECT 1530.950 16.560 1531.270 16.620 ;
        RECT 1510.250 16.420 1531.270 16.560 ;
        RECT 1510.250 16.360 1510.570 16.420 ;
        RECT 1530.950 16.360 1531.270 16.420 ;
      LAYER via ;
        RECT 1510.280 16.360 1510.540 16.620 ;
        RECT 1530.980 16.360 1531.240 16.620 ;
      LAYER met2 ;
        RECT 1508.570 510.410 1508.850 514.000 ;
        RECT 1508.570 510.270 1510.480 510.410 ;
        RECT 1508.570 510.000 1508.850 510.270 ;
        RECT 1510.340 16.650 1510.480 510.270 ;
        RECT 1510.280 16.330 1510.540 16.650 ;
        RECT 1530.980 16.330 1531.240 16.650 ;
        RECT 1531.040 2.400 1531.180 16.330 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.510 19.960 1524.830 20.020 ;
        RECT 1548.890 19.960 1549.210 20.020 ;
        RECT 1524.510 19.820 1549.210 19.960 ;
        RECT 1524.510 19.760 1524.830 19.820 ;
        RECT 1548.890 19.760 1549.210 19.820 ;
      LAYER via ;
        RECT 1524.540 19.760 1524.800 20.020 ;
        RECT 1548.920 19.760 1549.180 20.020 ;
      LAYER met2 ;
        RECT 1521.450 510.410 1521.730 514.000 ;
        RECT 1521.450 510.270 1524.740 510.410 ;
        RECT 1521.450 510.000 1521.730 510.270 ;
        RECT 1524.600 20.050 1524.740 510.270 ;
        RECT 1524.540 19.730 1524.800 20.050 ;
        RECT 1548.920 19.730 1549.180 20.050 ;
        RECT 1548.980 2.400 1549.120 19.730 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1537.850 14.860 1538.170 14.920 ;
        RECT 1566.830 14.860 1567.150 14.920 ;
        RECT 1537.850 14.720 1567.150 14.860 ;
        RECT 1537.850 14.660 1538.170 14.720 ;
        RECT 1566.830 14.660 1567.150 14.720 ;
      LAYER via ;
        RECT 1537.880 14.660 1538.140 14.920 ;
        RECT 1566.860 14.660 1567.120 14.920 ;
      LAYER met2 ;
        RECT 1534.330 510.410 1534.610 514.000 ;
        RECT 1534.330 510.270 1538.080 510.410 ;
        RECT 1534.330 510.000 1534.610 510.270 ;
        RECT 1537.940 14.950 1538.080 510.270 ;
        RECT 1537.880 14.630 1538.140 14.950 ;
        RECT 1566.860 14.630 1567.120 14.950 ;
        RECT 1566.920 2.400 1567.060 14.630 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1547.050 503.440 1547.370 503.500 ;
        RECT 1552.110 503.440 1552.430 503.500 ;
        RECT 1547.050 503.300 1552.430 503.440 ;
        RECT 1547.050 503.240 1547.370 503.300 ;
        RECT 1552.110 503.240 1552.430 503.300 ;
        RECT 1552.110 13.500 1552.430 13.560 ;
        RECT 1584.770 13.500 1585.090 13.560 ;
        RECT 1552.110 13.360 1585.090 13.500 ;
        RECT 1552.110 13.300 1552.430 13.360 ;
        RECT 1584.770 13.300 1585.090 13.360 ;
      LAYER via ;
        RECT 1547.080 503.240 1547.340 503.500 ;
        RECT 1552.140 503.240 1552.400 503.500 ;
        RECT 1552.140 13.300 1552.400 13.560 ;
        RECT 1584.800 13.300 1585.060 13.560 ;
      LAYER met2 ;
        RECT 1547.210 510.340 1547.490 514.000 ;
        RECT 1547.140 510.000 1547.490 510.340 ;
        RECT 1547.140 503.530 1547.280 510.000 ;
        RECT 1547.080 503.210 1547.340 503.530 ;
        RECT 1552.140 503.210 1552.400 503.530 ;
        RECT 1552.200 13.590 1552.340 503.210 ;
        RECT 1552.140 13.270 1552.400 13.590 ;
        RECT 1584.800 13.270 1585.060 13.590 ;
        RECT 1584.860 2.400 1585.000 13.270 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.470 503.440 1559.790 503.500 ;
        RECT 1565.450 503.440 1565.770 503.500 ;
        RECT 1559.470 503.300 1565.770 503.440 ;
        RECT 1559.470 503.240 1559.790 503.300 ;
        RECT 1565.450 503.240 1565.770 503.300 ;
        RECT 1565.450 19.960 1565.770 20.020 ;
        RECT 1602.250 19.960 1602.570 20.020 ;
        RECT 1565.450 19.820 1602.570 19.960 ;
        RECT 1565.450 19.760 1565.770 19.820 ;
        RECT 1602.250 19.760 1602.570 19.820 ;
      LAYER via ;
        RECT 1559.500 503.240 1559.760 503.500 ;
        RECT 1565.480 503.240 1565.740 503.500 ;
        RECT 1565.480 19.760 1565.740 20.020 ;
        RECT 1602.280 19.760 1602.540 20.020 ;
      LAYER met2 ;
        RECT 1559.630 510.340 1559.910 514.000 ;
        RECT 1559.560 510.000 1559.910 510.340 ;
        RECT 1559.560 503.530 1559.700 510.000 ;
        RECT 1559.500 503.210 1559.760 503.530 ;
        RECT 1565.480 503.210 1565.740 503.530 ;
        RECT 1565.540 20.050 1565.680 503.210 ;
        RECT 1565.480 19.730 1565.740 20.050 ;
        RECT 1602.280 19.730 1602.540 20.050 ;
        RECT 1602.340 2.400 1602.480 19.730 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.350 17.240 1572.670 17.300 ;
        RECT 1620.190 17.240 1620.510 17.300 ;
        RECT 1572.350 17.100 1620.510 17.240 ;
        RECT 1572.350 17.040 1572.670 17.100 ;
        RECT 1620.190 17.040 1620.510 17.100 ;
      LAYER via ;
        RECT 1572.380 17.040 1572.640 17.300 ;
        RECT 1620.220 17.040 1620.480 17.300 ;
      LAYER met2 ;
        RECT 1572.510 510.340 1572.790 514.000 ;
        RECT 1572.440 510.000 1572.790 510.340 ;
        RECT 1572.440 17.330 1572.580 510.000 ;
        RECT 1572.380 17.010 1572.640 17.330 ;
        RECT 1620.220 17.010 1620.480 17.330 ;
        RECT 1620.280 2.400 1620.420 17.010 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 18.940 1586.930 19.000 ;
        RECT 1638.130 18.940 1638.450 19.000 ;
        RECT 1586.610 18.800 1638.450 18.940 ;
        RECT 1586.610 18.740 1586.930 18.800 ;
        RECT 1638.130 18.740 1638.450 18.800 ;
      LAYER via ;
        RECT 1586.640 18.740 1586.900 19.000 ;
        RECT 1638.160 18.740 1638.420 19.000 ;
      LAYER met2 ;
        RECT 1585.390 510.410 1585.670 514.000 ;
        RECT 1585.390 510.270 1586.840 510.410 ;
        RECT 1585.390 510.000 1585.670 510.270 ;
        RECT 1586.700 19.030 1586.840 510.270 ;
        RECT 1586.640 18.710 1586.900 19.030 ;
        RECT 1638.160 18.710 1638.420 19.030 ;
        RECT 1638.220 2.400 1638.360 18.710 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.410 18.260 1600.730 18.320 ;
        RECT 1656.070 18.260 1656.390 18.320 ;
        RECT 1600.410 18.120 1656.390 18.260 ;
        RECT 1600.410 18.060 1600.730 18.120 ;
        RECT 1656.070 18.060 1656.390 18.120 ;
      LAYER via ;
        RECT 1600.440 18.060 1600.700 18.320 ;
        RECT 1656.100 18.060 1656.360 18.320 ;
      LAYER met2 ;
        RECT 1598.270 510.410 1598.550 514.000 ;
        RECT 1598.270 510.270 1600.640 510.410 ;
        RECT 1598.270 510.000 1598.550 510.270 ;
        RECT 1600.500 18.350 1600.640 510.270 ;
        RECT 1600.440 18.030 1600.700 18.350 ;
        RECT 1656.100 18.030 1656.360 18.350 ;
        RECT 1656.160 2.400 1656.300 18.030 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1614.670 17.920 1614.990 17.980 ;
        RECT 1673.550 17.920 1673.870 17.980 ;
        RECT 1614.670 17.780 1673.870 17.920 ;
        RECT 1614.670 17.720 1614.990 17.780 ;
        RECT 1673.550 17.720 1673.870 17.780 ;
      LAYER via ;
        RECT 1614.700 17.720 1614.960 17.980 ;
        RECT 1673.580 17.720 1673.840 17.980 ;
      LAYER met2 ;
        RECT 1611.150 510.410 1611.430 514.000 ;
        RECT 1611.150 510.270 1614.440 510.410 ;
        RECT 1611.150 510.000 1611.430 510.270 ;
        RECT 1614.300 20.810 1614.440 510.270 ;
        RECT 1614.300 20.670 1614.900 20.810 ;
        RECT 1614.760 18.010 1614.900 20.670 ;
        RECT 1614.700 17.690 1614.960 18.010 ;
        RECT 1673.580 17.690 1673.840 18.010 ;
        RECT 1673.640 2.400 1673.780 17.690 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1623.870 503.440 1624.190 503.500 ;
        RECT 1627.550 503.440 1627.870 503.500 ;
        RECT 1623.870 503.300 1627.870 503.440 ;
        RECT 1623.870 503.240 1624.190 503.300 ;
        RECT 1627.550 503.240 1627.870 503.300 ;
        RECT 1627.550 17.580 1627.870 17.640 ;
        RECT 1691.490 17.580 1691.810 17.640 ;
        RECT 1627.550 17.440 1691.810 17.580 ;
        RECT 1627.550 17.380 1627.870 17.440 ;
        RECT 1691.490 17.380 1691.810 17.440 ;
      LAYER via ;
        RECT 1623.900 503.240 1624.160 503.500 ;
        RECT 1627.580 503.240 1627.840 503.500 ;
        RECT 1627.580 17.380 1627.840 17.640 ;
        RECT 1691.520 17.380 1691.780 17.640 ;
      LAYER met2 ;
        RECT 1624.030 510.340 1624.310 514.000 ;
        RECT 1623.960 510.000 1624.310 510.340 ;
        RECT 1623.960 503.530 1624.100 510.000 ;
        RECT 1623.900 503.210 1624.160 503.530 ;
        RECT 1627.580 503.210 1627.840 503.530 ;
        RECT 1627.640 17.670 1627.780 503.210 ;
        RECT 1627.580 17.350 1627.840 17.670 ;
        RECT 1691.520 17.350 1691.780 17.670 ;
        RECT 1691.580 2.400 1691.720 17.350 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 731.010 148.140 731.330 148.200 ;
        RECT 931.570 148.140 931.890 148.200 ;
        RECT 731.010 148.000 931.890 148.140 ;
        RECT 731.010 147.940 731.330 148.000 ;
        RECT 931.570 147.940 931.890 148.000 ;
        RECT 728.250 17.580 728.570 17.640 ;
        RECT 731.010 17.580 731.330 17.640 ;
        RECT 728.250 17.440 731.330 17.580 ;
        RECT 728.250 17.380 728.570 17.440 ;
        RECT 731.010 17.380 731.330 17.440 ;
      LAYER via ;
        RECT 731.040 147.940 731.300 148.200 ;
        RECT 931.600 147.940 931.860 148.200 ;
        RECT 728.280 17.380 728.540 17.640 ;
        RECT 731.040 17.380 731.300 17.640 ;
      LAYER met2 ;
        RECT 932.190 510.410 932.470 514.000 ;
        RECT 931.660 510.270 932.470 510.410 ;
        RECT 931.660 148.230 931.800 510.270 ;
        RECT 932.190 510.000 932.470 510.270 ;
        RECT 731.040 147.910 731.300 148.230 ;
        RECT 931.600 147.910 931.860 148.230 ;
        RECT 731.100 17.670 731.240 147.910 ;
        RECT 728.280 17.350 728.540 17.670 ;
        RECT 731.040 17.350 731.300 17.670 ;
        RECT 728.340 2.400 728.480 17.350 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1636.290 503.440 1636.610 503.500 ;
        RECT 1641.810 503.440 1642.130 503.500 ;
        RECT 1636.290 503.300 1642.130 503.440 ;
        RECT 1636.290 503.240 1636.610 503.300 ;
        RECT 1641.810 503.240 1642.130 503.300 ;
        RECT 1641.810 19.280 1642.130 19.340 ;
        RECT 1709.430 19.280 1709.750 19.340 ;
        RECT 1641.810 19.140 1709.750 19.280 ;
        RECT 1641.810 19.080 1642.130 19.140 ;
        RECT 1709.430 19.080 1709.750 19.140 ;
      LAYER via ;
        RECT 1636.320 503.240 1636.580 503.500 ;
        RECT 1641.840 503.240 1642.100 503.500 ;
        RECT 1641.840 19.080 1642.100 19.340 ;
        RECT 1709.460 19.080 1709.720 19.340 ;
      LAYER met2 ;
        RECT 1636.450 510.340 1636.730 514.000 ;
        RECT 1636.380 510.000 1636.730 510.340 ;
        RECT 1636.380 503.530 1636.520 510.000 ;
        RECT 1636.320 503.210 1636.580 503.530 ;
        RECT 1641.840 503.210 1642.100 503.530 ;
        RECT 1641.900 19.370 1642.040 503.210 ;
        RECT 1641.840 19.050 1642.100 19.370 ;
        RECT 1709.460 19.050 1709.720 19.370 ;
        RECT 1709.520 2.400 1709.660 19.050 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1649.170 503.440 1649.490 503.500 ;
        RECT 1655.150 503.440 1655.470 503.500 ;
        RECT 1649.170 503.300 1655.470 503.440 ;
        RECT 1649.170 503.240 1649.490 503.300 ;
        RECT 1655.150 503.240 1655.470 503.300 ;
        RECT 1655.150 58.720 1655.470 58.780 ;
        RECT 1725.070 58.720 1725.390 58.780 ;
        RECT 1655.150 58.580 1725.390 58.720 ;
        RECT 1655.150 58.520 1655.470 58.580 ;
        RECT 1725.070 58.520 1725.390 58.580 ;
      LAYER via ;
        RECT 1649.200 503.240 1649.460 503.500 ;
        RECT 1655.180 503.240 1655.440 503.500 ;
        RECT 1655.180 58.520 1655.440 58.780 ;
        RECT 1725.100 58.520 1725.360 58.780 ;
      LAYER met2 ;
        RECT 1649.330 510.340 1649.610 514.000 ;
        RECT 1649.260 510.000 1649.610 510.340 ;
        RECT 1649.260 503.530 1649.400 510.000 ;
        RECT 1649.200 503.210 1649.460 503.530 ;
        RECT 1655.180 503.210 1655.440 503.530 ;
        RECT 1655.240 58.810 1655.380 503.210 ;
        RECT 1655.180 58.490 1655.440 58.810 ;
        RECT 1725.100 58.490 1725.360 58.810 ;
        RECT 1725.160 3.130 1725.300 58.490 ;
        RECT 1725.160 2.990 1727.600 3.130 ;
        RECT 1727.460 2.400 1727.600 2.990 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1661.665 282.965 1661.835 331.075 ;
        RECT 1661.665 234.685 1661.835 241.995 ;
      LAYER mcon ;
        RECT 1661.665 330.905 1661.835 331.075 ;
        RECT 1661.665 241.825 1661.835 241.995 ;
      LAYER met1 ;
        RECT 1661.590 448.700 1661.910 448.760 ;
        RECT 1662.510 448.700 1662.830 448.760 ;
        RECT 1661.590 448.560 1662.830 448.700 ;
        RECT 1661.590 448.500 1661.910 448.560 ;
        RECT 1662.510 448.500 1662.830 448.560 ;
        RECT 1662.510 400.420 1662.830 400.480 ;
        RECT 1662.140 400.280 1662.830 400.420 ;
        RECT 1662.140 400.140 1662.280 400.280 ;
        RECT 1662.510 400.220 1662.830 400.280 ;
        RECT 1662.050 399.880 1662.370 400.140 ;
        RECT 1662.050 362.340 1662.370 362.400 ;
        RECT 1662.970 362.340 1663.290 362.400 ;
        RECT 1662.050 362.200 1663.290 362.340 ;
        RECT 1662.050 362.140 1662.370 362.200 ;
        RECT 1662.970 362.140 1663.290 362.200 ;
        RECT 1661.590 331.060 1661.910 331.120 ;
        RECT 1661.395 330.920 1661.910 331.060 ;
        RECT 1661.590 330.860 1661.910 330.920 ;
        RECT 1661.605 283.120 1661.895 283.165 ;
        RECT 1662.050 283.120 1662.370 283.180 ;
        RECT 1661.605 282.980 1662.370 283.120 ;
        RECT 1661.605 282.935 1661.895 282.980 ;
        RECT 1662.050 282.920 1662.370 282.980 ;
        RECT 1661.605 241.980 1661.895 242.025 ;
        RECT 1662.050 241.980 1662.370 242.040 ;
        RECT 1661.605 241.840 1662.370 241.980 ;
        RECT 1661.605 241.795 1661.895 241.840 ;
        RECT 1662.050 241.780 1662.370 241.840 ;
        RECT 1661.590 234.840 1661.910 234.900 ;
        RECT 1661.395 234.700 1661.910 234.840 ;
        RECT 1661.590 234.640 1661.910 234.700 ;
        RECT 1661.590 234.160 1661.910 234.220 ;
        RECT 1662.050 234.160 1662.370 234.220 ;
        RECT 1661.590 234.020 1662.370 234.160 ;
        RECT 1661.590 233.960 1661.910 234.020 ;
        RECT 1662.050 233.960 1662.370 234.020 ;
        RECT 1662.050 159.020 1662.370 159.080 ;
        RECT 1661.680 158.880 1662.370 159.020 ;
        RECT 1661.680 158.740 1661.820 158.880 ;
        RECT 1662.050 158.820 1662.370 158.880 ;
        RECT 1661.590 158.480 1661.910 158.740 ;
        RECT 1661.590 110.540 1661.910 110.800 ;
        RECT 1661.680 110.120 1661.820 110.540 ;
        RECT 1661.590 109.860 1661.910 110.120 ;
        RECT 1661.590 65.520 1661.910 65.580 ;
        RECT 1738.870 65.520 1739.190 65.580 ;
        RECT 1661.590 65.380 1739.190 65.520 ;
        RECT 1661.590 65.320 1661.910 65.380 ;
        RECT 1738.870 65.320 1739.190 65.380 ;
        RECT 1738.870 17.920 1739.190 17.980 ;
        RECT 1745.310 17.920 1745.630 17.980 ;
        RECT 1738.870 17.780 1745.630 17.920 ;
        RECT 1738.870 17.720 1739.190 17.780 ;
        RECT 1745.310 17.720 1745.630 17.780 ;
      LAYER via ;
        RECT 1661.620 448.500 1661.880 448.760 ;
        RECT 1662.540 448.500 1662.800 448.760 ;
        RECT 1662.540 400.220 1662.800 400.480 ;
        RECT 1662.080 399.880 1662.340 400.140 ;
        RECT 1662.080 362.140 1662.340 362.400 ;
        RECT 1663.000 362.140 1663.260 362.400 ;
        RECT 1661.620 330.860 1661.880 331.120 ;
        RECT 1662.080 282.920 1662.340 283.180 ;
        RECT 1662.080 241.780 1662.340 242.040 ;
        RECT 1661.620 234.640 1661.880 234.900 ;
        RECT 1661.620 233.960 1661.880 234.220 ;
        RECT 1662.080 233.960 1662.340 234.220 ;
        RECT 1662.080 158.820 1662.340 159.080 ;
        RECT 1661.620 158.480 1661.880 158.740 ;
        RECT 1661.620 110.540 1661.880 110.800 ;
        RECT 1661.620 109.860 1661.880 110.120 ;
        RECT 1661.620 65.320 1661.880 65.580 ;
        RECT 1738.900 65.320 1739.160 65.580 ;
        RECT 1738.900 17.720 1739.160 17.980 ;
        RECT 1745.340 17.720 1745.600 17.980 ;
      LAYER met2 ;
        RECT 1662.210 510.410 1662.490 514.000 ;
        RECT 1661.680 510.270 1662.490 510.410 ;
        RECT 1661.680 483.325 1661.820 510.270 ;
        RECT 1662.210 510.000 1662.490 510.270 ;
        RECT 1661.610 482.955 1661.890 483.325 ;
        RECT 1662.530 482.955 1662.810 483.325 ;
        RECT 1662.600 448.790 1662.740 482.955 ;
        RECT 1661.620 448.530 1661.880 448.790 ;
        RECT 1662.540 448.530 1662.800 448.790 ;
        RECT 1661.620 448.470 1662.800 448.530 ;
        RECT 1661.680 448.390 1662.740 448.470 ;
        RECT 1662.600 400.510 1662.740 448.390 ;
        RECT 1662.540 400.190 1662.800 400.510 ;
        RECT 1662.080 399.850 1662.340 400.170 ;
        RECT 1662.140 362.430 1662.280 399.850 ;
        RECT 1662.080 362.110 1662.340 362.430 ;
        RECT 1663.000 362.110 1663.260 362.430 ;
        RECT 1663.060 338.485 1663.200 362.110 ;
        RECT 1662.070 338.370 1662.350 338.485 ;
        RECT 1661.680 338.230 1662.350 338.370 ;
        RECT 1661.680 331.150 1661.820 338.230 ;
        RECT 1662.070 338.115 1662.350 338.230 ;
        RECT 1662.990 338.115 1663.270 338.485 ;
        RECT 1661.620 330.830 1661.880 331.150 ;
        RECT 1662.080 282.890 1662.340 283.210 ;
        RECT 1662.140 242.070 1662.280 282.890 ;
        RECT 1662.080 241.750 1662.340 242.070 ;
        RECT 1661.620 234.610 1661.880 234.930 ;
        RECT 1661.680 234.250 1661.820 234.610 ;
        RECT 1661.620 233.930 1661.880 234.250 ;
        RECT 1662.080 233.930 1662.340 234.250 ;
        RECT 1662.140 159.110 1662.280 233.930 ;
        RECT 1662.080 158.790 1662.340 159.110 ;
        RECT 1661.620 158.450 1661.880 158.770 ;
        RECT 1661.680 110.830 1661.820 158.450 ;
        RECT 1661.620 110.510 1661.880 110.830 ;
        RECT 1661.620 109.830 1661.880 110.150 ;
        RECT 1661.680 65.610 1661.820 109.830 ;
        RECT 1661.620 65.290 1661.880 65.610 ;
        RECT 1738.900 65.290 1739.160 65.610 ;
        RECT 1738.960 18.010 1739.100 65.290 ;
        RECT 1738.900 17.690 1739.160 18.010 ;
        RECT 1745.340 17.690 1745.600 18.010 ;
        RECT 1745.400 2.400 1745.540 17.690 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 1661.610 483.000 1661.890 483.280 ;
        RECT 1662.530 483.000 1662.810 483.280 ;
        RECT 1662.070 338.160 1662.350 338.440 ;
        RECT 1662.990 338.160 1663.270 338.440 ;
      LAYER met3 ;
        RECT 1661.585 483.290 1661.915 483.305 ;
        RECT 1662.505 483.290 1662.835 483.305 ;
        RECT 1661.585 482.990 1662.835 483.290 ;
        RECT 1661.585 482.975 1661.915 482.990 ;
        RECT 1662.505 482.975 1662.835 482.990 ;
        RECT 1662.045 338.450 1662.375 338.465 ;
        RECT 1662.965 338.450 1663.295 338.465 ;
        RECT 1662.045 338.150 1663.295 338.450 ;
        RECT 1662.045 338.135 1662.375 338.150 ;
        RECT 1662.965 338.135 1663.295 338.150 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1675.850 79.460 1676.170 79.520 ;
        RECT 1759.570 79.460 1759.890 79.520 ;
        RECT 1675.850 79.320 1759.890 79.460 ;
        RECT 1675.850 79.260 1676.170 79.320 ;
        RECT 1759.570 79.260 1759.890 79.320 ;
        RECT 1759.570 2.960 1759.890 3.020 ;
        RECT 1762.790 2.960 1763.110 3.020 ;
        RECT 1759.570 2.820 1763.110 2.960 ;
        RECT 1759.570 2.760 1759.890 2.820 ;
        RECT 1762.790 2.760 1763.110 2.820 ;
      LAYER via ;
        RECT 1675.880 79.260 1676.140 79.520 ;
        RECT 1759.600 79.260 1759.860 79.520 ;
        RECT 1759.600 2.760 1759.860 3.020 ;
        RECT 1762.820 2.760 1763.080 3.020 ;
      LAYER met2 ;
        RECT 1675.090 510.410 1675.370 514.000 ;
        RECT 1675.090 510.270 1676.080 510.410 ;
        RECT 1675.090 510.000 1675.370 510.270 ;
        RECT 1675.940 79.550 1676.080 510.270 ;
        RECT 1675.880 79.230 1676.140 79.550 ;
        RECT 1759.600 79.230 1759.860 79.550 ;
        RECT 1759.660 3.050 1759.800 79.230 ;
        RECT 1759.600 2.730 1759.860 3.050 ;
        RECT 1762.820 2.730 1763.080 3.050 ;
        RECT 1762.880 2.400 1763.020 2.730 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1687.810 500.720 1688.130 500.780 ;
        RECT 1693.790 500.720 1694.110 500.780 ;
        RECT 1687.810 500.580 1694.110 500.720 ;
        RECT 1687.810 500.520 1688.130 500.580 ;
        RECT 1693.790 500.520 1694.110 500.580 ;
        RECT 1693.790 44.780 1694.110 44.840 ;
        RECT 1780.730 44.780 1781.050 44.840 ;
        RECT 1693.790 44.640 1781.050 44.780 ;
        RECT 1693.790 44.580 1694.110 44.640 ;
        RECT 1780.730 44.580 1781.050 44.640 ;
      LAYER via ;
        RECT 1687.840 500.520 1688.100 500.780 ;
        RECT 1693.820 500.520 1694.080 500.780 ;
        RECT 1693.820 44.580 1694.080 44.840 ;
        RECT 1780.760 44.580 1781.020 44.840 ;
      LAYER met2 ;
        RECT 1687.970 510.340 1688.250 514.000 ;
        RECT 1687.900 510.000 1688.250 510.340 ;
        RECT 1687.900 500.810 1688.040 510.000 ;
        RECT 1687.840 500.490 1688.100 500.810 ;
        RECT 1693.820 500.490 1694.080 500.810 ;
        RECT 1693.880 44.870 1694.020 500.490 ;
        RECT 1693.820 44.550 1694.080 44.870 ;
        RECT 1780.760 44.550 1781.020 44.870 ;
        RECT 1780.820 2.400 1780.960 44.550 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1798.745 2.805 1798.915 48.195 ;
      LAYER mcon ;
        RECT 1798.745 48.025 1798.915 48.195 ;
      LAYER met1 ;
        RECT 1703.910 86.260 1704.230 86.320 ;
        RECT 1794.070 86.260 1794.390 86.320 ;
        RECT 1703.910 86.120 1794.390 86.260 ;
        RECT 1703.910 86.060 1704.230 86.120 ;
        RECT 1794.070 86.060 1794.390 86.120 ;
        RECT 1794.070 48.180 1794.390 48.240 ;
        RECT 1798.685 48.180 1798.975 48.225 ;
        RECT 1794.070 48.040 1798.975 48.180 ;
        RECT 1794.070 47.980 1794.390 48.040 ;
        RECT 1798.685 47.995 1798.975 48.040 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1798.475 2.820 1798.990 2.960 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 1703.940 86.060 1704.200 86.320 ;
        RECT 1794.100 86.060 1794.360 86.320 ;
        RECT 1794.100 47.980 1794.360 48.240 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 1700.850 510.410 1701.130 514.000 ;
        RECT 1700.850 510.270 1704.140 510.410 ;
        RECT 1700.850 510.000 1701.130 510.270 ;
        RECT 1704.000 86.350 1704.140 510.270 ;
        RECT 1703.940 86.030 1704.200 86.350 ;
        RECT 1794.100 86.030 1794.360 86.350 ;
        RECT 1794.160 48.270 1794.300 86.030 ;
        RECT 1794.100 47.950 1794.360 48.270 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1713.110 503.100 1713.430 503.160 ;
        RECT 1735.190 503.100 1735.510 503.160 ;
        RECT 1713.110 502.960 1735.510 503.100 ;
        RECT 1713.110 502.900 1713.430 502.960 ;
        RECT 1735.190 502.900 1735.510 502.960 ;
        RECT 1735.190 58.720 1735.510 58.780 ;
        RECT 1814.770 58.720 1815.090 58.780 ;
        RECT 1735.190 58.580 1815.090 58.720 ;
        RECT 1735.190 58.520 1735.510 58.580 ;
        RECT 1814.770 58.520 1815.090 58.580 ;
      LAYER via ;
        RECT 1713.140 502.900 1713.400 503.160 ;
        RECT 1735.220 502.900 1735.480 503.160 ;
        RECT 1735.220 58.520 1735.480 58.780 ;
        RECT 1814.800 58.520 1815.060 58.780 ;
      LAYER met2 ;
        RECT 1713.270 510.340 1713.550 514.000 ;
        RECT 1713.200 510.000 1713.550 510.340 ;
        RECT 1713.200 503.190 1713.340 510.000 ;
        RECT 1713.140 502.870 1713.400 503.190 ;
        RECT 1735.220 502.870 1735.480 503.190 ;
        RECT 1735.280 58.810 1735.420 502.870 ;
        RECT 1735.220 58.490 1735.480 58.810 ;
        RECT 1814.800 58.490 1815.060 58.810 ;
        RECT 1814.860 16.050 1815.000 58.490 ;
        RECT 1814.860 15.910 1816.840 16.050 ;
        RECT 1816.700 2.400 1816.840 15.910 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1725.990 503.440 1726.310 503.500 ;
        RECT 1731.050 503.440 1731.370 503.500 ;
        RECT 1725.990 503.300 1731.370 503.440 ;
        RECT 1725.990 503.240 1726.310 503.300 ;
        RECT 1731.050 503.240 1731.370 503.300 ;
        RECT 1731.050 93.060 1731.370 93.120 ;
        RECT 1828.570 93.060 1828.890 93.120 ;
        RECT 1731.050 92.920 1828.890 93.060 ;
        RECT 1731.050 92.860 1731.370 92.920 ;
        RECT 1828.570 92.860 1828.890 92.920 ;
        RECT 1828.570 19.280 1828.890 19.340 ;
        RECT 1834.550 19.280 1834.870 19.340 ;
        RECT 1828.570 19.140 1834.870 19.280 ;
        RECT 1828.570 19.080 1828.890 19.140 ;
        RECT 1834.550 19.080 1834.870 19.140 ;
      LAYER via ;
        RECT 1726.020 503.240 1726.280 503.500 ;
        RECT 1731.080 503.240 1731.340 503.500 ;
        RECT 1731.080 92.860 1731.340 93.120 ;
        RECT 1828.600 92.860 1828.860 93.120 ;
        RECT 1828.600 19.080 1828.860 19.340 ;
        RECT 1834.580 19.080 1834.840 19.340 ;
      LAYER met2 ;
        RECT 1726.150 510.340 1726.430 514.000 ;
        RECT 1726.080 510.000 1726.430 510.340 ;
        RECT 1726.080 503.530 1726.220 510.000 ;
        RECT 1726.020 503.210 1726.280 503.530 ;
        RECT 1731.080 503.210 1731.340 503.530 ;
        RECT 1731.140 93.150 1731.280 503.210 ;
        RECT 1731.080 92.830 1731.340 93.150 ;
        RECT 1828.600 92.830 1828.860 93.150 ;
        RECT 1828.660 19.370 1828.800 92.830 ;
        RECT 1828.600 19.050 1828.860 19.370 ;
        RECT 1834.580 19.050 1834.840 19.370 ;
        RECT 1834.640 2.400 1834.780 19.050 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.870 503.100 1739.190 503.160 ;
        RECT 1744.850 503.100 1745.170 503.160 ;
        RECT 1738.870 502.960 1745.170 503.100 ;
        RECT 1738.870 502.900 1739.190 502.960 ;
        RECT 1744.850 502.900 1745.170 502.960 ;
        RECT 1744.850 107.000 1745.170 107.060 ;
        RECT 1849.270 107.000 1849.590 107.060 ;
        RECT 1744.850 106.860 1849.590 107.000 ;
        RECT 1744.850 106.800 1745.170 106.860 ;
        RECT 1849.270 106.800 1849.590 106.860 ;
      LAYER via ;
        RECT 1738.900 502.900 1739.160 503.160 ;
        RECT 1744.880 502.900 1745.140 503.160 ;
        RECT 1744.880 106.800 1745.140 107.060 ;
        RECT 1849.300 106.800 1849.560 107.060 ;
      LAYER met2 ;
        RECT 1739.030 510.340 1739.310 514.000 ;
        RECT 1738.960 510.000 1739.310 510.340 ;
        RECT 1738.960 503.190 1739.100 510.000 ;
        RECT 1738.900 502.870 1739.160 503.190 ;
        RECT 1744.880 502.870 1745.140 503.190 ;
        RECT 1744.940 107.090 1745.080 502.870 ;
        RECT 1744.880 106.770 1745.140 107.090 ;
        RECT 1849.300 106.770 1849.560 107.090 ;
        RECT 1849.360 17.410 1849.500 106.770 ;
        RECT 1849.360 17.270 1852.260 17.410 ;
        RECT 1852.120 2.400 1852.260 17.270 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1750.905 379.525 1751.075 400.775 ;
        RECT 1750.905 319.345 1751.075 331.075 ;
        RECT 1751.825 158.185 1751.995 220.575 ;
      LAYER mcon ;
        RECT 1750.905 400.605 1751.075 400.775 ;
        RECT 1750.905 330.905 1751.075 331.075 ;
        RECT 1751.825 220.405 1751.995 220.575 ;
      LAYER met1 ;
        RECT 1750.845 400.760 1751.135 400.805 ;
        RECT 1751.290 400.760 1751.610 400.820 ;
        RECT 1750.845 400.620 1751.610 400.760 ;
        RECT 1750.845 400.575 1751.135 400.620 ;
        RECT 1751.290 400.560 1751.610 400.620 ;
        RECT 1750.830 379.680 1751.150 379.740 ;
        RECT 1750.635 379.540 1751.150 379.680 ;
        RECT 1750.830 379.480 1751.150 379.540 ;
        RECT 1750.830 338.200 1751.150 338.260 ;
        RECT 1751.750 338.200 1752.070 338.260 ;
        RECT 1750.830 338.060 1752.070 338.200 ;
        RECT 1750.830 338.000 1751.150 338.060 ;
        RECT 1751.750 338.000 1752.070 338.060 ;
        RECT 1750.845 331.060 1751.135 331.105 ;
        RECT 1751.750 331.060 1752.070 331.120 ;
        RECT 1750.845 330.920 1752.070 331.060 ;
        RECT 1750.845 330.875 1751.135 330.920 ;
        RECT 1751.750 330.860 1752.070 330.920 ;
        RECT 1750.845 319.500 1751.135 319.545 ;
        RECT 1751.750 319.500 1752.070 319.560 ;
        RECT 1750.845 319.360 1752.070 319.500 ;
        RECT 1750.845 319.315 1751.135 319.360 ;
        RECT 1751.750 319.300 1752.070 319.360 ;
        RECT 1751.750 221.240 1752.070 221.300 ;
        RECT 1752.670 221.240 1752.990 221.300 ;
        RECT 1751.750 221.100 1752.990 221.240 ;
        RECT 1751.750 221.040 1752.070 221.100 ;
        RECT 1752.670 221.040 1752.990 221.100 ;
        RECT 1751.750 220.560 1752.070 220.620 ;
        RECT 1751.555 220.420 1752.070 220.560 ;
        RECT 1751.750 220.360 1752.070 220.420 ;
        RECT 1751.750 158.340 1752.070 158.400 ;
        RECT 1751.555 158.200 1752.070 158.340 ;
        RECT 1751.750 158.140 1752.070 158.200 ;
        RECT 1751.290 83.200 1751.610 83.260 ;
        RECT 1751.750 83.200 1752.070 83.260 ;
        RECT 1751.290 83.060 1752.070 83.200 ;
        RECT 1751.290 83.000 1751.610 83.060 ;
        RECT 1751.750 83.000 1752.070 83.060 ;
        RECT 1751.290 65.520 1751.610 65.580 ;
        RECT 1870.430 65.520 1870.750 65.580 ;
        RECT 1751.290 65.380 1870.750 65.520 ;
        RECT 1751.290 65.320 1751.610 65.380 ;
        RECT 1870.430 65.320 1870.750 65.380 ;
      LAYER via ;
        RECT 1751.320 400.560 1751.580 400.820 ;
        RECT 1750.860 379.480 1751.120 379.740 ;
        RECT 1750.860 338.000 1751.120 338.260 ;
        RECT 1751.780 338.000 1752.040 338.260 ;
        RECT 1751.780 330.860 1752.040 331.120 ;
        RECT 1751.780 319.300 1752.040 319.560 ;
        RECT 1751.780 221.040 1752.040 221.300 ;
        RECT 1752.700 221.040 1752.960 221.300 ;
        RECT 1751.780 220.360 1752.040 220.620 ;
        RECT 1751.780 158.140 1752.040 158.400 ;
        RECT 1751.320 83.000 1751.580 83.260 ;
        RECT 1751.780 83.000 1752.040 83.260 ;
        RECT 1751.320 65.320 1751.580 65.580 ;
        RECT 1870.460 65.320 1870.720 65.580 ;
      LAYER met2 ;
        RECT 1751.910 511.090 1752.190 514.000 ;
        RECT 1751.910 510.950 1752.900 511.090 ;
        RECT 1751.910 510.000 1752.190 510.950 ;
        RECT 1752.760 483.210 1752.900 510.950 ;
        RECT 1752.300 483.070 1752.900 483.210 ;
        RECT 1752.300 435.045 1752.440 483.070 ;
        RECT 1751.310 434.675 1751.590 435.045 ;
        RECT 1752.230 434.675 1752.510 435.045 ;
        RECT 1751.380 400.850 1751.520 434.675 ;
        RECT 1751.320 400.530 1751.580 400.850 ;
        RECT 1750.860 379.450 1751.120 379.770 ;
        RECT 1750.920 338.290 1751.060 379.450 ;
        RECT 1750.860 337.970 1751.120 338.290 ;
        RECT 1751.780 337.970 1752.040 338.290 ;
        RECT 1751.840 331.150 1751.980 337.970 ;
        RECT 1751.780 330.830 1752.040 331.150 ;
        RECT 1751.780 319.270 1752.040 319.590 ;
        RECT 1751.840 270.485 1751.980 319.270 ;
        RECT 1751.770 270.115 1752.050 270.485 ;
        RECT 1751.770 269.435 1752.050 269.805 ;
        RECT 1751.840 269.125 1751.980 269.435 ;
        RECT 1751.770 268.755 1752.050 269.125 ;
        RECT 1752.690 268.755 1752.970 269.125 ;
        RECT 1752.760 221.330 1752.900 268.755 ;
        RECT 1751.780 221.010 1752.040 221.330 ;
        RECT 1752.700 221.010 1752.960 221.330 ;
        RECT 1751.840 220.650 1751.980 221.010 ;
        RECT 1751.780 220.330 1752.040 220.650 ;
        RECT 1751.780 158.110 1752.040 158.430 ;
        RECT 1751.840 83.290 1751.980 158.110 ;
        RECT 1751.320 82.970 1751.580 83.290 ;
        RECT 1751.780 82.970 1752.040 83.290 ;
        RECT 1751.380 65.610 1751.520 82.970 ;
        RECT 1751.320 65.290 1751.580 65.610 ;
        RECT 1870.460 65.290 1870.720 65.610 ;
        RECT 1870.520 7.210 1870.660 65.290 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
      LAYER via2 ;
        RECT 1751.310 434.720 1751.590 435.000 ;
        RECT 1752.230 434.720 1752.510 435.000 ;
        RECT 1751.770 270.160 1752.050 270.440 ;
        RECT 1751.770 269.480 1752.050 269.760 ;
        RECT 1751.770 268.800 1752.050 269.080 ;
        RECT 1752.690 268.800 1752.970 269.080 ;
      LAYER met3 ;
        RECT 1751.285 435.010 1751.615 435.025 ;
        RECT 1752.205 435.010 1752.535 435.025 ;
        RECT 1751.285 434.710 1752.535 435.010 ;
        RECT 1751.285 434.695 1751.615 434.710 ;
        RECT 1752.205 434.695 1752.535 434.710 ;
        RECT 1751.745 270.450 1752.075 270.465 ;
        RECT 1751.070 270.150 1752.075 270.450 ;
        RECT 1751.070 269.770 1751.370 270.150 ;
        RECT 1751.745 270.135 1752.075 270.150 ;
        RECT 1751.745 269.770 1752.075 269.785 ;
        RECT 1751.070 269.470 1752.075 269.770 ;
        RECT 1751.745 269.455 1752.075 269.470 ;
        RECT 1751.745 269.090 1752.075 269.105 ;
        RECT 1752.665 269.090 1752.995 269.105 ;
        RECT 1751.745 268.790 1752.995 269.090 ;
        RECT 1751.745 268.775 1752.075 268.790 ;
        RECT 1752.665 268.775 1752.995 268.790 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 155.280 752.030 155.340 ;
        RECT 938.930 155.280 939.250 155.340 ;
        RECT 751.710 155.140 939.250 155.280 ;
        RECT 751.710 155.080 752.030 155.140 ;
        RECT 938.930 155.080 939.250 155.140 ;
        RECT 746.190 20.640 746.510 20.700 ;
        RECT 751.710 20.640 752.030 20.700 ;
        RECT 746.190 20.500 752.030 20.640 ;
        RECT 746.190 20.440 746.510 20.500 ;
        RECT 751.710 20.440 752.030 20.500 ;
      LAYER via ;
        RECT 751.740 155.080 752.000 155.340 ;
        RECT 938.960 155.080 939.220 155.340 ;
        RECT 746.220 20.440 746.480 20.700 ;
        RECT 751.740 20.440 752.000 20.700 ;
      LAYER met2 ;
        RECT 945.070 511.090 945.350 514.000 ;
        RECT 941.780 510.950 945.350 511.090 ;
        RECT 941.780 490.010 941.920 510.950 ;
        RECT 945.070 510.000 945.350 510.950 ;
        RECT 939.020 489.870 941.920 490.010 ;
        RECT 939.020 155.370 939.160 489.870 ;
        RECT 751.740 155.050 752.000 155.370 ;
        RECT 938.960 155.050 939.220 155.370 ;
        RECT 751.800 20.730 751.940 155.050 ;
        RECT 746.220 20.410 746.480 20.730 ;
        RECT 751.740 20.410 752.000 20.730 ;
        RECT 746.280 2.400 746.420 20.410 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1765.550 113.800 1765.870 113.860 ;
        RECT 1883.770 113.800 1884.090 113.860 ;
        RECT 1765.550 113.660 1884.090 113.800 ;
        RECT 1765.550 113.600 1765.870 113.660 ;
        RECT 1883.770 113.600 1884.090 113.660 ;
      LAYER via ;
        RECT 1765.580 113.600 1765.840 113.860 ;
        RECT 1883.800 113.600 1884.060 113.860 ;
      LAYER met2 ;
        RECT 1764.790 510.410 1765.070 514.000 ;
        RECT 1764.790 510.270 1765.780 510.410 ;
        RECT 1764.790 510.000 1765.070 510.270 ;
        RECT 1765.640 113.890 1765.780 510.270 ;
        RECT 1765.580 113.570 1765.840 113.890 ;
        RECT 1883.800 113.570 1884.060 113.890 ;
        RECT 1883.860 16.730 1884.000 113.570 ;
        RECT 1883.860 16.590 1888.140 16.730 ;
        RECT 1888.000 2.400 1888.140 16.590 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 79.460 1780.130 79.520 ;
        RECT 1904.470 79.460 1904.790 79.520 ;
        RECT 1779.810 79.320 1904.790 79.460 ;
        RECT 1779.810 79.260 1780.130 79.320 ;
        RECT 1904.470 79.260 1904.790 79.320 ;
      LAYER via ;
        RECT 1779.840 79.260 1780.100 79.520 ;
        RECT 1904.500 79.260 1904.760 79.520 ;
      LAYER met2 ;
        RECT 1777.670 510.410 1777.950 514.000 ;
        RECT 1777.670 510.270 1780.040 510.410 ;
        RECT 1777.670 510.000 1777.950 510.270 ;
        RECT 1779.900 79.550 1780.040 510.270 ;
        RECT 1779.840 79.230 1780.100 79.550 ;
        RECT 1904.500 79.230 1904.760 79.550 ;
        RECT 1904.560 16.730 1904.700 79.230 ;
        RECT 1904.560 16.590 1906.080 16.730 ;
        RECT 1905.940 2.400 1906.080 16.590 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1793.610 72.320 1793.930 72.380 ;
        RECT 1918.270 72.320 1918.590 72.380 ;
        RECT 1793.610 72.180 1918.590 72.320 ;
        RECT 1793.610 72.120 1793.930 72.180 ;
        RECT 1918.270 72.120 1918.590 72.180 ;
      LAYER via ;
        RECT 1793.640 72.120 1793.900 72.380 ;
        RECT 1918.300 72.120 1918.560 72.380 ;
      LAYER met2 ;
        RECT 1790.090 510.410 1790.370 514.000 ;
        RECT 1790.090 510.270 1793.840 510.410 ;
        RECT 1790.090 510.000 1790.370 510.270 ;
        RECT 1793.700 72.410 1793.840 510.270 ;
        RECT 1793.640 72.090 1793.900 72.410 ;
        RECT 1918.300 72.090 1918.560 72.410 ;
        RECT 1918.360 17.410 1918.500 72.090 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1802.810 500.380 1803.130 500.440 ;
        RECT 1852.490 500.380 1852.810 500.440 ;
        RECT 1802.810 500.240 1852.810 500.380 ;
        RECT 1802.810 500.180 1803.130 500.240 ;
        RECT 1852.490 500.180 1852.810 500.240 ;
        RECT 1852.490 99.860 1852.810 99.920 ;
        RECT 1938.970 99.860 1939.290 99.920 ;
        RECT 1852.490 99.720 1939.290 99.860 ;
        RECT 1852.490 99.660 1852.810 99.720 ;
        RECT 1938.970 99.660 1939.290 99.720 ;
      LAYER via ;
        RECT 1802.840 500.180 1803.100 500.440 ;
        RECT 1852.520 500.180 1852.780 500.440 ;
        RECT 1852.520 99.660 1852.780 99.920 ;
        RECT 1939.000 99.660 1939.260 99.920 ;
      LAYER met2 ;
        RECT 1802.970 510.340 1803.250 514.000 ;
        RECT 1802.900 510.000 1803.250 510.340 ;
        RECT 1802.900 500.470 1803.040 510.000 ;
        RECT 1802.840 500.150 1803.100 500.470 ;
        RECT 1852.520 500.150 1852.780 500.470 ;
        RECT 1852.580 99.950 1852.720 500.150 ;
        RECT 1852.520 99.630 1852.780 99.950 ;
        RECT 1939.000 99.630 1939.260 99.950 ;
        RECT 1939.060 17.410 1939.200 99.630 ;
        RECT 1939.060 17.270 1941.500 17.410 ;
        RECT 1941.360 2.400 1941.500 17.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1815.690 496.980 1816.010 497.040 ;
        RECT 1820.750 496.980 1821.070 497.040 ;
        RECT 1815.690 496.840 1821.070 496.980 ;
        RECT 1815.690 496.780 1816.010 496.840 ;
        RECT 1820.750 496.780 1821.070 496.840 ;
        RECT 1820.750 86.260 1821.070 86.320 ;
        RECT 1952.770 86.260 1953.090 86.320 ;
        RECT 1820.750 86.120 1953.090 86.260 ;
        RECT 1820.750 86.060 1821.070 86.120 ;
        RECT 1952.770 86.060 1953.090 86.120 ;
        RECT 1952.770 38.320 1953.090 38.380 ;
        RECT 1959.210 38.320 1959.530 38.380 ;
        RECT 1952.770 38.180 1959.530 38.320 ;
        RECT 1952.770 38.120 1953.090 38.180 ;
        RECT 1959.210 38.120 1959.530 38.180 ;
      LAYER via ;
        RECT 1815.720 496.780 1815.980 497.040 ;
        RECT 1820.780 496.780 1821.040 497.040 ;
        RECT 1820.780 86.060 1821.040 86.320 ;
        RECT 1952.800 86.060 1953.060 86.320 ;
        RECT 1952.800 38.120 1953.060 38.380 ;
        RECT 1959.240 38.120 1959.500 38.380 ;
      LAYER met2 ;
        RECT 1815.850 510.340 1816.130 514.000 ;
        RECT 1815.780 510.000 1816.130 510.340 ;
        RECT 1815.780 497.070 1815.920 510.000 ;
        RECT 1815.720 496.750 1815.980 497.070 ;
        RECT 1820.780 496.750 1821.040 497.070 ;
        RECT 1820.840 86.350 1820.980 496.750 ;
        RECT 1820.780 86.030 1821.040 86.350 ;
        RECT 1952.800 86.030 1953.060 86.350 ;
        RECT 1952.860 38.410 1953.000 86.030 ;
        RECT 1952.800 38.090 1953.060 38.410 ;
        RECT 1959.240 38.090 1959.500 38.410 ;
        RECT 1959.300 2.400 1959.440 38.090 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1977.225 48.365 1977.395 93.075 ;
      LAYER mcon ;
        RECT 1977.225 92.905 1977.395 93.075 ;
      LAYER met1 ;
        RECT 1828.570 496.980 1828.890 497.040 ;
        RECT 1835.010 496.980 1835.330 497.040 ;
        RECT 1828.570 496.840 1835.330 496.980 ;
        RECT 1828.570 496.780 1828.890 496.840 ;
        RECT 1835.010 496.780 1835.330 496.840 ;
        RECT 1835.010 93.060 1835.330 93.120 ;
        RECT 1977.165 93.060 1977.455 93.105 ;
        RECT 1835.010 92.920 1977.455 93.060 ;
        RECT 1835.010 92.860 1835.330 92.920 ;
        RECT 1977.165 92.875 1977.455 92.920 ;
        RECT 1977.150 48.520 1977.470 48.580 ;
        RECT 1976.955 48.380 1977.470 48.520 ;
        RECT 1977.150 48.320 1977.470 48.380 ;
      LAYER via ;
        RECT 1828.600 496.780 1828.860 497.040 ;
        RECT 1835.040 496.780 1835.300 497.040 ;
        RECT 1835.040 92.860 1835.300 93.120 ;
        RECT 1977.180 48.320 1977.440 48.580 ;
      LAYER met2 ;
        RECT 1828.730 510.340 1829.010 514.000 ;
        RECT 1828.660 510.000 1829.010 510.340 ;
        RECT 1828.660 497.070 1828.800 510.000 ;
        RECT 1828.600 496.750 1828.860 497.070 ;
        RECT 1835.040 496.750 1835.300 497.070 ;
        RECT 1835.100 93.150 1835.240 496.750 ;
        RECT 1835.040 92.830 1835.300 93.150 ;
        RECT 1977.180 48.290 1977.440 48.610 ;
        RECT 1977.240 2.400 1977.380 48.290 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1841.450 120.600 1841.770 120.660 ;
        RECT 1994.170 120.600 1994.490 120.660 ;
        RECT 1841.450 120.460 1994.490 120.600 ;
        RECT 1841.450 120.400 1841.770 120.460 ;
        RECT 1994.170 120.400 1994.490 120.460 ;
        RECT 1994.170 62.260 1994.490 62.520 ;
        RECT 1994.260 61.780 1994.400 62.260 ;
        RECT 1995.090 61.780 1995.410 61.840 ;
        RECT 1994.260 61.640 1995.410 61.780 ;
        RECT 1995.090 61.580 1995.410 61.640 ;
        RECT 1995.090 47.980 1995.410 48.240 ;
        RECT 1995.180 47.560 1995.320 47.980 ;
        RECT 1995.090 47.300 1995.410 47.560 ;
      LAYER via ;
        RECT 1841.480 120.400 1841.740 120.660 ;
        RECT 1994.200 120.400 1994.460 120.660 ;
        RECT 1994.200 62.260 1994.460 62.520 ;
        RECT 1995.120 61.580 1995.380 61.840 ;
        RECT 1995.120 47.980 1995.380 48.240 ;
        RECT 1995.120 47.300 1995.380 47.560 ;
      LAYER met2 ;
        RECT 1841.610 510.340 1841.890 514.000 ;
        RECT 1841.540 510.000 1841.890 510.340 ;
        RECT 1841.540 120.690 1841.680 510.000 ;
        RECT 1841.480 120.370 1841.740 120.690 ;
        RECT 1994.200 120.370 1994.460 120.690 ;
        RECT 1994.260 62.550 1994.400 120.370 ;
        RECT 1994.200 62.230 1994.460 62.550 ;
        RECT 1995.120 61.550 1995.380 61.870 ;
        RECT 1995.180 48.270 1995.320 61.550 ;
        RECT 1995.120 47.950 1995.380 48.270 ;
        RECT 1995.120 47.270 1995.380 47.590 ;
        RECT 1995.180 2.400 1995.320 47.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 107.000 1856.030 107.060 ;
        RECT 2007.970 107.000 2008.290 107.060 ;
        RECT 1855.710 106.860 2008.290 107.000 ;
        RECT 1855.710 106.800 1856.030 106.860 ;
        RECT 2007.970 106.800 2008.290 106.860 ;
        RECT 2007.970 62.120 2008.290 62.180 ;
        RECT 2012.570 62.120 2012.890 62.180 ;
        RECT 2007.970 61.980 2012.890 62.120 ;
        RECT 2007.970 61.920 2008.290 61.980 ;
        RECT 2012.570 61.920 2012.890 61.980 ;
      LAYER via ;
        RECT 1855.740 106.800 1856.000 107.060 ;
        RECT 2008.000 106.800 2008.260 107.060 ;
        RECT 2008.000 61.920 2008.260 62.180 ;
        RECT 2012.600 61.920 2012.860 62.180 ;
      LAYER met2 ;
        RECT 1854.490 510.410 1854.770 514.000 ;
        RECT 1854.490 510.270 1855.940 510.410 ;
        RECT 1854.490 510.000 1854.770 510.270 ;
        RECT 1855.800 107.090 1855.940 510.270 ;
        RECT 1855.740 106.770 1856.000 107.090 ;
        RECT 2008.000 106.770 2008.260 107.090 ;
        RECT 2008.060 62.210 2008.200 106.770 ;
        RECT 2008.000 61.890 2008.260 62.210 ;
        RECT 2012.600 61.890 2012.860 62.210 ;
        RECT 2012.660 2.400 2012.800 61.890 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2030.585 2.805 2030.755 48.195 ;
      LAYER mcon ;
        RECT 2030.585 48.025 2030.755 48.195 ;
      LAYER met1 ;
        RECT 1869.510 127.740 1869.830 127.800 ;
        RECT 2028.670 127.740 2028.990 127.800 ;
        RECT 1869.510 127.600 2028.990 127.740 ;
        RECT 1869.510 127.540 1869.830 127.600 ;
        RECT 2028.670 127.540 2028.990 127.600 ;
        RECT 2030.510 48.180 2030.830 48.240 ;
        RECT 2030.315 48.040 2030.830 48.180 ;
        RECT 2030.510 47.980 2030.830 48.040 ;
        RECT 2030.510 2.960 2030.830 3.020 ;
        RECT 2030.315 2.820 2030.830 2.960 ;
        RECT 2030.510 2.760 2030.830 2.820 ;
      LAYER via ;
        RECT 1869.540 127.540 1869.800 127.800 ;
        RECT 2028.700 127.540 2028.960 127.800 ;
        RECT 2030.540 47.980 2030.800 48.240 ;
        RECT 2030.540 2.760 2030.800 3.020 ;
      LAYER met2 ;
        RECT 1866.910 510.410 1867.190 514.000 ;
        RECT 1866.910 510.270 1869.740 510.410 ;
        RECT 1866.910 510.000 1867.190 510.270 ;
        RECT 1869.600 127.830 1869.740 510.270 ;
        RECT 1869.540 127.510 1869.800 127.830 ;
        RECT 2028.700 127.510 2028.960 127.830 ;
        RECT 2028.760 72.490 2028.900 127.510 ;
        RECT 2028.760 72.350 2029.360 72.490 ;
        RECT 2029.220 61.610 2029.360 72.350 ;
        RECT 2029.220 61.470 2030.740 61.610 ;
        RECT 2030.600 48.270 2030.740 61.470 ;
        RECT 2030.540 47.950 2030.800 48.270 ;
        RECT 2030.540 2.730 2030.800 3.050 ;
        RECT 2030.600 2.400 2030.740 2.730 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1879.630 500.040 1879.950 500.100 ;
        RECT 1886.990 500.040 1887.310 500.100 ;
        RECT 1879.630 499.900 1887.310 500.040 ;
        RECT 1879.630 499.840 1879.950 499.900 ;
        RECT 1886.990 499.840 1887.310 499.900 ;
        RECT 1886.990 113.800 1887.310 113.860 ;
        RECT 2042.470 113.800 2042.790 113.860 ;
        RECT 1886.990 113.660 2042.790 113.800 ;
        RECT 1886.990 113.600 1887.310 113.660 ;
        RECT 2042.470 113.600 2042.790 113.660 ;
        RECT 2042.470 38.320 2042.790 38.380 ;
        RECT 2048.450 38.320 2048.770 38.380 ;
        RECT 2042.470 38.180 2048.770 38.320 ;
        RECT 2042.470 38.120 2042.790 38.180 ;
        RECT 2048.450 38.120 2048.770 38.180 ;
      LAYER via ;
        RECT 1879.660 499.840 1879.920 500.100 ;
        RECT 1887.020 499.840 1887.280 500.100 ;
        RECT 1887.020 113.600 1887.280 113.860 ;
        RECT 2042.500 113.600 2042.760 113.860 ;
        RECT 2042.500 38.120 2042.760 38.380 ;
        RECT 2048.480 38.120 2048.740 38.380 ;
      LAYER met2 ;
        RECT 1879.790 510.340 1880.070 514.000 ;
        RECT 1879.720 510.000 1880.070 510.340 ;
        RECT 1879.720 500.130 1879.860 510.000 ;
        RECT 1879.660 499.810 1879.920 500.130 ;
        RECT 1887.020 499.810 1887.280 500.130 ;
        RECT 1887.080 113.890 1887.220 499.810 ;
        RECT 1887.020 113.570 1887.280 113.890 ;
        RECT 2042.500 113.570 2042.760 113.890 ;
        RECT 2042.560 38.410 2042.700 113.570 ;
        RECT 2042.500 38.090 2042.760 38.410 ;
        RECT 2048.480 38.090 2048.740 38.410 ;
        RECT 2048.540 2.400 2048.680 38.090 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.510 162.080 765.830 162.140 ;
        RECT 952.730 162.080 953.050 162.140 ;
        RECT 765.510 161.940 953.050 162.080 ;
        RECT 765.510 161.880 765.830 161.940 ;
        RECT 952.730 161.880 953.050 161.940 ;
      LAYER via ;
        RECT 765.540 161.880 765.800 162.140 ;
        RECT 952.760 161.880 953.020 162.140 ;
      LAYER met2 ;
        RECT 957.950 511.090 958.230 514.000 ;
        RECT 954.660 510.950 958.230 511.090 ;
        RECT 954.660 490.010 954.800 510.950 ;
        RECT 957.950 510.000 958.230 510.950 ;
        RECT 952.820 489.870 954.800 490.010 ;
        RECT 952.820 162.170 952.960 489.870 ;
        RECT 765.540 161.850 765.800 162.170 ;
        RECT 952.760 161.850 953.020 162.170 ;
        RECT 765.600 3.130 765.740 161.850 ;
        RECT 763.760 2.990 765.740 3.130 ;
        RECT 763.760 2.400 763.900 2.990 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1892.510 472.500 1892.830 472.560 ;
        RECT 2063.170 472.500 2063.490 472.560 ;
        RECT 1892.510 472.360 2063.490 472.500 ;
        RECT 1892.510 472.300 1892.830 472.360 ;
        RECT 2063.170 472.300 2063.490 472.360 ;
        RECT 2063.170 62.120 2063.490 62.180 ;
        RECT 2066.390 62.120 2066.710 62.180 ;
        RECT 2063.170 61.980 2066.710 62.120 ;
        RECT 2063.170 61.920 2063.490 61.980 ;
        RECT 2066.390 61.920 2066.710 61.980 ;
      LAYER via ;
        RECT 1892.540 472.300 1892.800 472.560 ;
        RECT 2063.200 472.300 2063.460 472.560 ;
        RECT 2063.200 61.920 2063.460 62.180 ;
        RECT 2066.420 61.920 2066.680 62.180 ;
      LAYER met2 ;
        RECT 1892.670 510.340 1892.950 514.000 ;
        RECT 1892.600 510.000 1892.950 510.340 ;
        RECT 1892.600 472.590 1892.740 510.000 ;
        RECT 1892.540 472.270 1892.800 472.590 ;
        RECT 2063.200 472.270 2063.460 472.590 ;
        RECT 2063.260 62.210 2063.400 472.270 ;
        RECT 2063.200 61.890 2063.460 62.210 ;
        RECT 2066.420 61.890 2066.680 62.210 ;
        RECT 2066.480 2.400 2066.620 61.890 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1905.390 499.360 1905.710 499.420 ;
        RECT 1910.910 499.360 1911.230 499.420 ;
        RECT 1905.390 499.220 1911.230 499.360 ;
        RECT 1905.390 499.160 1905.710 499.220 ;
        RECT 1910.910 499.160 1911.230 499.220 ;
        RECT 1910.910 134.540 1911.230 134.600 ;
        RECT 2084.330 134.540 2084.650 134.600 ;
        RECT 1910.910 134.400 2084.650 134.540 ;
        RECT 1910.910 134.340 1911.230 134.400 ;
        RECT 2084.330 134.340 2084.650 134.400 ;
      LAYER via ;
        RECT 1905.420 499.160 1905.680 499.420 ;
        RECT 1910.940 499.160 1911.200 499.420 ;
        RECT 1910.940 134.340 1911.200 134.600 ;
        RECT 2084.360 134.340 2084.620 134.600 ;
      LAYER met2 ;
        RECT 1905.550 510.340 1905.830 514.000 ;
        RECT 1905.480 510.000 1905.830 510.340 ;
        RECT 1905.480 499.450 1905.620 510.000 ;
        RECT 1905.420 499.130 1905.680 499.450 ;
        RECT 1910.940 499.130 1911.200 499.450 ;
        RECT 1911.000 134.630 1911.140 499.130 ;
        RECT 1910.940 134.310 1911.200 134.630 ;
        RECT 2084.360 134.310 2084.620 134.630 ;
        RECT 2084.420 2.400 2084.560 134.310 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1918.270 503.440 1918.590 503.500 ;
        RECT 1924.710 503.440 1925.030 503.500 ;
        RECT 1918.270 503.300 1925.030 503.440 ;
        RECT 1918.270 503.240 1918.590 503.300 ;
        RECT 1924.710 503.240 1925.030 503.300 ;
        RECT 1924.710 141.340 1925.030 141.400 ;
        RECT 2097.670 141.340 2097.990 141.400 ;
        RECT 1924.710 141.200 2097.990 141.340 ;
        RECT 1924.710 141.140 1925.030 141.200 ;
        RECT 2097.670 141.140 2097.990 141.200 ;
        RECT 2097.670 62.120 2097.990 62.180 ;
        RECT 2101.810 62.120 2102.130 62.180 ;
        RECT 2097.670 61.980 2102.130 62.120 ;
        RECT 2097.670 61.920 2097.990 61.980 ;
        RECT 2101.810 61.920 2102.130 61.980 ;
      LAYER via ;
        RECT 1918.300 503.240 1918.560 503.500 ;
        RECT 1924.740 503.240 1925.000 503.500 ;
        RECT 1924.740 141.140 1925.000 141.400 ;
        RECT 2097.700 141.140 2097.960 141.400 ;
        RECT 2097.700 61.920 2097.960 62.180 ;
        RECT 2101.840 61.920 2102.100 62.180 ;
      LAYER met2 ;
        RECT 1918.430 510.340 1918.710 514.000 ;
        RECT 1918.360 510.000 1918.710 510.340 ;
        RECT 1918.360 503.530 1918.500 510.000 ;
        RECT 1918.300 503.210 1918.560 503.530 ;
        RECT 1924.740 503.210 1925.000 503.530 ;
        RECT 1924.800 141.430 1924.940 503.210 ;
        RECT 1924.740 141.110 1925.000 141.430 ;
        RECT 2097.700 141.110 2097.960 141.430 ;
        RECT 2097.760 62.210 2097.900 141.110 ;
        RECT 2097.700 61.890 2097.960 62.210 ;
        RECT 2101.840 61.890 2102.100 62.210 ;
        RECT 2101.900 2.400 2102.040 61.890 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1930.765 241.485 1930.935 280.075 ;
        RECT 1931.225 147.985 1931.395 193.035 ;
      LAYER mcon ;
        RECT 1930.765 279.905 1930.935 280.075 ;
        RECT 1931.225 192.865 1931.395 193.035 ;
      LAYER met1 ;
        RECT 1930.690 496.640 1931.010 496.700 ;
        RECT 1931.610 496.640 1931.930 496.700 ;
        RECT 1930.690 496.500 1931.930 496.640 ;
        RECT 1930.690 496.440 1931.010 496.500 ;
        RECT 1931.610 496.440 1931.930 496.500 ;
        RECT 1930.690 379.680 1931.010 379.740 ;
        RECT 1931.610 379.680 1931.930 379.740 ;
        RECT 1930.690 379.540 1931.930 379.680 ;
        RECT 1930.690 379.480 1931.010 379.540 ;
        RECT 1931.610 379.480 1931.930 379.540 ;
        RECT 1930.690 280.060 1931.010 280.120 ;
        RECT 1930.495 279.920 1931.010 280.060 ;
        RECT 1930.690 279.860 1931.010 279.920 ;
        RECT 1930.705 241.640 1930.995 241.685 ;
        RECT 1931.610 241.640 1931.930 241.700 ;
        RECT 1930.705 241.500 1931.930 241.640 ;
        RECT 1930.705 241.455 1930.995 241.500 ;
        RECT 1931.610 241.440 1931.930 241.500 ;
        RECT 1931.610 207.300 1931.930 207.360 ;
        RECT 1931.240 207.160 1931.930 207.300 ;
        RECT 1931.240 207.020 1931.380 207.160 ;
        RECT 1931.610 207.100 1931.930 207.160 ;
        RECT 1931.150 206.760 1931.470 207.020 ;
        RECT 1931.150 193.020 1931.470 193.080 ;
        RECT 1930.955 192.880 1931.470 193.020 ;
        RECT 1931.150 192.820 1931.470 192.880 ;
        RECT 1931.165 148.140 1931.455 148.185 ;
        RECT 2118.370 148.140 2118.690 148.200 ;
        RECT 1931.165 148.000 2118.690 148.140 ;
        RECT 1931.165 147.955 1931.455 148.000 ;
        RECT 2118.370 147.940 2118.690 148.000 ;
      LAYER via ;
        RECT 1930.720 496.440 1930.980 496.700 ;
        RECT 1931.640 496.440 1931.900 496.700 ;
        RECT 1930.720 379.480 1930.980 379.740 ;
        RECT 1931.640 379.480 1931.900 379.740 ;
        RECT 1930.720 279.860 1930.980 280.120 ;
        RECT 1931.640 241.440 1931.900 241.700 ;
        RECT 1931.640 207.100 1931.900 207.360 ;
        RECT 1931.180 206.760 1931.440 207.020 ;
        RECT 1931.180 192.820 1931.440 193.080 ;
        RECT 2118.400 147.940 2118.660 148.200 ;
      LAYER met2 ;
        RECT 1931.310 510.410 1931.590 514.000 ;
        RECT 1930.780 510.270 1931.590 510.410 ;
        RECT 1930.780 496.730 1930.920 510.270 ;
        RECT 1931.310 510.000 1931.590 510.270 ;
        RECT 1930.720 496.410 1930.980 496.730 ;
        RECT 1931.640 496.410 1931.900 496.730 ;
        RECT 1931.700 379.770 1931.840 496.410 ;
        RECT 1930.720 379.450 1930.980 379.770 ;
        RECT 1931.640 379.450 1931.900 379.770 ;
        RECT 1930.780 280.150 1930.920 379.450 ;
        RECT 1930.720 279.830 1930.980 280.150 ;
        RECT 1931.640 241.410 1931.900 241.730 ;
        RECT 1931.700 207.390 1931.840 241.410 ;
        RECT 1931.640 207.070 1931.900 207.390 ;
        RECT 1931.180 206.730 1931.440 207.050 ;
        RECT 1931.240 193.110 1931.380 206.730 ;
        RECT 1931.180 192.790 1931.440 193.110 ;
        RECT 2118.400 147.910 2118.660 148.230 ;
        RECT 2118.460 3.130 2118.600 147.910 ;
        RECT 2118.460 2.990 2119.980 3.130 ;
        RECT 2119.840 2.400 2119.980 2.990 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1944.950 155.280 1945.270 155.340 ;
        RECT 2132.170 155.280 2132.490 155.340 ;
        RECT 1944.950 155.140 2132.490 155.280 ;
        RECT 1944.950 155.080 1945.270 155.140 ;
        RECT 2132.170 155.080 2132.490 155.140 ;
        RECT 2132.170 62.120 2132.490 62.180 ;
        RECT 2137.690 62.120 2138.010 62.180 ;
        RECT 2132.170 61.980 2138.010 62.120 ;
        RECT 2132.170 61.920 2132.490 61.980 ;
        RECT 2137.690 61.920 2138.010 61.980 ;
      LAYER via ;
        RECT 1944.980 155.080 1945.240 155.340 ;
        RECT 2132.200 155.080 2132.460 155.340 ;
        RECT 2132.200 61.920 2132.460 62.180 ;
        RECT 2137.720 61.920 2137.980 62.180 ;
      LAYER met2 ;
        RECT 1943.730 510.410 1944.010 514.000 ;
        RECT 1943.730 510.270 1945.180 510.410 ;
        RECT 1943.730 510.000 1944.010 510.270 ;
        RECT 1945.040 155.370 1945.180 510.270 ;
        RECT 1944.980 155.050 1945.240 155.370 ;
        RECT 2132.200 155.050 2132.460 155.370 ;
        RECT 2132.260 62.210 2132.400 155.050 ;
        RECT 2132.200 61.890 2132.460 62.210 ;
        RECT 2137.720 61.890 2137.980 62.210 ;
        RECT 2137.780 2.400 2137.920 61.890 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2155.705 2.805 2155.875 48.195 ;
      LAYER mcon ;
        RECT 2155.705 48.025 2155.875 48.195 ;
      LAYER met1 ;
        RECT 1959.210 168.880 1959.530 168.940 ;
        RECT 2152.870 168.880 2153.190 168.940 ;
        RECT 1959.210 168.740 2153.190 168.880 ;
        RECT 1959.210 168.680 1959.530 168.740 ;
        RECT 2152.870 168.680 2153.190 168.740 ;
        RECT 2152.870 62.120 2153.190 62.180 ;
        RECT 2155.630 62.120 2155.950 62.180 ;
        RECT 2152.870 61.980 2155.950 62.120 ;
        RECT 2152.870 61.920 2153.190 61.980 ;
        RECT 2155.630 61.920 2155.950 61.980 ;
        RECT 2155.630 48.180 2155.950 48.240 ;
        RECT 2155.435 48.040 2155.950 48.180 ;
        RECT 2155.630 47.980 2155.950 48.040 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2155.435 2.820 2155.950 2.960 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1959.240 168.680 1959.500 168.940 ;
        RECT 2152.900 168.680 2153.160 168.940 ;
        RECT 2152.900 61.920 2153.160 62.180 ;
        RECT 2155.660 61.920 2155.920 62.180 ;
        RECT 2155.660 47.980 2155.920 48.240 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1956.610 510.410 1956.890 514.000 ;
        RECT 1956.610 510.270 1959.440 510.410 ;
        RECT 1956.610 510.000 1956.890 510.270 ;
        RECT 1959.300 168.970 1959.440 510.270 ;
        RECT 1959.240 168.650 1959.500 168.970 ;
        RECT 2152.900 168.650 2153.160 168.970 ;
        RECT 2152.960 62.210 2153.100 168.650 ;
        RECT 2152.900 61.890 2153.160 62.210 ;
        RECT 2155.660 61.890 2155.920 62.210 ;
        RECT 2155.720 48.270 2155.860 61.890 ;
        RECT 2155.660 47.950 2155.920 48.270 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 176.020 1973.330 176.080 ;
        RECT 2166.670 176.020 2166.990 176.080 ;
        RECT 1973.010 175.880 2166.990 176.020 ;
        RECT 1973.010 175.820 1973.330 175.880 ;
        RECT 2166.670 175.820 2166.990 175.880 ;
        RECT 2166.670 30.160 2166.990 30.220 ;
        RECT 2173.110 30.160 2173.430 30.220 ;
        RECT 2166.670 30.020 2173.430 30.160 ;
        RECT 2166.670 29.960 2166.990 30.020 ;
        RECT 2173.110 29.960 2173.430 30.020 ;
      LAYER via ;
        RECT 1973.040 175.820 1973.300 176.080 ;
        RECT 2166.700 175.820 2166.960 176.080 ;
        RECT 2166.700 29.960 2166.960 30.220 ;
        RECT 2173.140 29.960 2173.400 30.220 ;
      LAYER met2 ;
        RECT 1969.490 510.410 1969.770 514.000 ;
        RECT 1969.490 510.270 1973.240 510.410 ;
        RECT 1969.490 510.000 1969.770 510.270 ;
        RECT 1973.100 176.110 1973.240 510.270 ;
        RECT 1973.040 175.790 1973.300 176.110 ;
        RECT 2166.700 175.790 2166.960 176.110 ;
        RECT 2166.760 30.250 2166.900 175.790 ;
        RECT 2166.700 29.930 2166.960 30.250 ;
        RECT 2173.140 29.930 2173.400 30.250 ;
        RECT 2173.200 2.400 2173.340 29.930 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1982.210 496.980 1982.530 497.040 ;
        RECT 1986.810 496.980 1987.130 497.040 ;
        RECT 1982.210 496.840 1987.130 496.980 ;
        RECT 1982.210 496.780 1982.530 496.840 ;
        RECT 1986.810 496.780 1987.130 496.840 ;
        RECT 1986.810 444.960 1987.130 445.020 ;
        RECT 2187.370 444.960 2187.690 445.020 ;
        RECT 1986.810 444.820 2187.690 444.960 ;
        RECT 1986.810 444.760 1987.130 444.820 ;
        RECT 2187.370 444.760 2187.690 444.820 ;
      LAYER via ;
        RECT 1982.240 496.780 1982.500 497.040 ;
        RECT 1986.840 496.780 1987.100 497.040 ;
        RECT 1986.840 444.760 1987.100 445.020 ;
        RECT 2187.400 444.760 2187.660 445.020 ;
      LAYER met2 ;
        RECT 1982.370 510.340 1982.650 514.000 ;
        RECT 1982.300 510.000 1982.650 510.340 ;
        RECT 1982.300 497.070 1982.440 510.000 ;
        RECT 1982.240 496.750 1982.500 497.070 ;
        RECT 1986.840 496.750 1987.100 497.070 ;
        RECT 1986.900 445.050 1987.040 496.750 ;
        RECT 1986.840 444.730 1987.100 445.050 ;
        RECT 2187.400 444.730 2187.660 445.050 ;
        RECT 2187.460 17.410 2187.600 444.730 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 496.980 1995.410 497.040 ;
        RECT 2000.150 496.980 2000.470 497.040 ;
        RECT 1995.090 496.840 2000.470 496.980 ;
        RECT 1995.090 496.780 1995.410 496.840 ;
        RECT 2000.150 496.780 2000.470 496.840 ;
        RECT 2000.150 451.760 2000.470 451.820 ;
        RECT 2208.070 451.760 2208.390 451.820 ;
        RECT 2000.150 451.620 2208.390 451.760 ;
        RECT 2000.150 451.560 2000.470 451.620 ;
        RECT 2208.070 451.560 2208.390 451.620 ;
      LAYER via ;
        RECT 1995.120 496.780 1995.380 497.040 ;
        RECT 2000.180 496.780 2000.440 497.040 ;
        RECT 2000.180 451.560 2000.440 451.820 ;
        RECT 2208.100 451.560 2208.360 451.820 ;
      LAYER met2 ;
        RECT 1995.250 510.340 1995.530 514.000 ;
        RECT 1995.180 510.000 1995.530 510.340 ;
        RECT 1995.180 497.070 1995.320 510.000 ;
        RECT 1995.120 496.750 1995.380 497.070 ;
        RECT 2000.180 496.750 2000.440 497.070 ;
        RECT 2000.240 451.850 2000.380 496.750 ;
        RECT 2000.180 451.530 2000.440 451.850 ;
        RECT 2208.100 451.530 2208.360 451.850 ;
        RECT 2208.160 17.410 2208.300 451.530 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.970 496.980 2008.290 497.040 ;
        RECT 2013.950 496.980 2014.270 497.040 ;
        RECT 2007.970 496.840 2014.270 496.980 ;
        RECT 2007.970 496.780 2008.290 496.840 ;
        RECT 2013.950 496.780 2014.270 496.840 ;
        RECT 2013.950 196.760 2014.270 196.820 ;
        RECT 2221.870 196.760 2222.190 196.820 ;
        RECT 2013.950 196.620 2222.190 196.760 ;
        RECT 2013.950 196.560 2014.270 196.620 ;
        RECT 2221.870 196.560 2222.190 196.620 ;
      LAYER via ;
        RECT 2008.000 496.780 2008.260 497.040 ;
        RECT 2013.980 496.780 2014.240 497.040 ;
        RECT 2013.980 196.560 2014.240 196.820 ;
        RECT 2221.900 196.560 2222.160 196.820 ;
      LAYER met2 ;
        RECT 2008.130 510.340 2008.410 514.000 ;
        RECT 2008.060 510.000 2008.410 510.340 ;
        RECT 2008.060 497.070 2008.200 510.000 ;
        RECT 2008.000 496.750 2008.260 497.070 ;
        RECT 2013.980 496.750 2014.240 497.070 ;
        RECT 2014.040 196.850 2014.180 496.750 ;
        RECT 2013.980 196.530 2014.240 196.850 ;
        RECT 2221.900 196.530 2222.160 196.850 ;
        RECT 2221.960 17.410 2222.100 196.530 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 168.880 786.530 168.940 ;
        RECT 966.530 168.880 966.850 168.940 ;
        RECT 786.210 168.740 966.850 168.880 ;
        RECT 786.210 168.680 786.530 168.740 ;
        RECT 966.530 168.680 966.850 168.740 ;
        RECT 781.610 14.520 781.930 14.580 ;
        RECT 786.210 14.520 786.530 14.580 ;
        RECT 781.610 14.380 786.530 14.520 ;
        RECT 781.610 14.320 781.930 14.380 ;
        RECT 786.210 14.320 786.530 14.380 ;
      LAYER via ;
        RECT 786.240 168.680 786.500 168.940 ;
        RECT 966.560 168.680 966.820 168.940 ;
        RECT 781.640 14.320 781.900 14.580 ;
        RECT 786.240 14.320 786.500 14.580 ;
      LAYER met2 ;
        RECT 970.830 511.090 971.110 514.000 ;
        RECT 967.540 510.950 971.110 511.090 ;
        RECT 967.540 490.010 967.680 510.950 ;
        RECT 970.830 510.000 971.110 510.950 ;
        RECT 966.620 489.870 967.680 490.010 ;
        RECT 966.620 168.970 966.760 489.870 ;
        RECT 786.240 168.650 786.500 168.970 ;
        RECT 966.560 168.650 966.820 168.970 ;
        RECT 786.300 14.610 786.440 168.650 ;
        RECT 781.640 14.290 781.900 14.610 ;
        RECT 786.240 14.290 786.500 14.610 ;
        RECT 781.700 2.400 781.840 14.290 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2021.310 65.520 2021.630 65.580 ;
        RECT 2242.570 65.520 2242.890 65.580 ;
        RECT 2021.310 65.380 2242.890 65.520 ;
        RECT 2021.310 65.320 2021.630 65.380 ;
        RECT 2242.570 65.320 2242.890 65.380 ;
      LAYER via ;
        RECT 2021.340 65.320 2021.600 65.580 ;
        RECT 2242.600 65.320 2242.860 65.580 ;
      LAYER met2 ;
        RECT 2020.550 510.410 2020.830 514.000 ;
        RECT 2020.550 510.270 2021.540 510.410 ;
        RECT 2020.550 510.000 2020.830 510.270 ;
        RECT 2021.400 65.610 2021.540 510.270 ;
        RECT 2021.340 65.290 2021.600 65.610 ;
        RECT 2242.600 65.290 2242.860 65.610 ;
        RECT 2242.660 17.410 2242.800 65.290 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2034.650 203.560 2034.970 203.620 ;
        RECT 2256.370 203.560 2256.690 203.620 ;
        RECT 2034.650 203.420 2256.690 203.560 ;
        RECT 2034.650 203.360 2034.970 203.420 ;
        RECT 2256.370 203.360 2256.690 203.420 ;
        RECT 2256.370 16.900 2256.690 16.960 ;
        RECT 2262.350 16.900 2262.670 16.960 ;
        RECT 2256.370 16.760 2262.670 16.900 ;
        RECT 2256.370 16.700 2256.690 16.760 ;
        RECT 2262.350 16.700 2262.670 16.760 ;
      LAYER via ;
        RECT 2034.680 203.360 2034.940 203.620 ;
        RECT 2256.400 203.360 2256.660 203.620 ;
        RECT 2256.400 16.700 2256.660 16.960 ;
        RECT 2262.380 16.700 2262.640 16.960 ;
      LAYER met2 ;
        RECT 2033.430 510.410 2033.710 514.000 ;
        RECT 2033.430 510.270 2034.880 510.410 ;
        RECT 2033.430 510.000 2033.710 510.270 ;
        RECT 2034.740 203.650 2034.880 510.270 ;
        RECT 2034.680 203.330 2034.940 203.650 ;
        RECT 2256.400 203.330 2256.660 203.650 ;
        RECT 2256.460 16.990 2256.600 203.330 ;
        RECT 2256.400 16.670 2256.660 16.990 ;
        RECT 2262.380 16.670 2262.640 16.990 ;
        RECT 2262.440 2.400 2262.580 16.670 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2048.910 217.160 2049.230 217.220 ;
        RECT 2277.070 217.160 2277.390 217.220 ;
        RECT 2048.910 217.020 2277.390 217.160 ;
        RECT 2048.910 216.960 2049.230 217.020 ;
        RECT 2277.070 216.960 2277.390 217.020 ;
      LAYER via ;
        RECT 2048.940 216.960 2049.200 217.220 ;
        RECT 2277.100 216.960 2277.360 217.220 ;
      LAYER met2 ;
        RECT 2046.310 510.410 2046.590 514.000 ;
        RECT 2046.310 510.270 2049.140 510.410 ;
        RECT 2046.310 510.000 2046.590 510.270 ;
        RECT 2049.000 217.250 2049.140 510.270 ;
        RECT 2048.940 216.930 2049.200 217.250 ;
        RECT 2277.100 216.930 2277.360 217.250 ;
        RECT 2277.160 17.410 2277.300 216.930 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2059.030 496.980 2059.350 497.040 ;
        RECT 2062.710 496.980 2063.030 497.040 ;
        RECT 2059.030 496.840 2063.030 496.980 ;
        RECT 2059.030 496.780 2059.350 496.840 ;
        RECT 2062.710 496.780 2063.030 496.840 ;
        RECT 2062.710 231.100 2063.030 231.160 ;
        RECT 2298.230 231.100 2298.550 231.160 ;
        RECT 2062.710 230.960 2298.550 231.100 ;
        RECT 2062.710 230.900 2063.030 230.960 ;
        RECT 2298.230 230.900 2298.550 230.960 ;
      LAYER via ;
        RECT 2059.060 496.780 2059.320 497.040 ;
        RECT 2062.740 496.780 2063.000 497.040 ;
        RECT 2062.740 230.900 2063.000 231.160 ;
        RECT 2298.260 230.900 2298.520 231.160 ;
      LAYER met2 ;
        RECT 2059.190 510.340 2059.470 514.000 ;
        RECT 2059.120 510.000 2059.470 510.340 ;
        RECT 2059.120 497.070 2059.260 510.000 ;
        RECT 2059.060 496.750 2059.320 497.070 ;
        RECT 2062.740 496.750 2063.000 497.070 ;
        RECT 2062.800 231.190 2062.940 496.750 ;
        RECT 2062.740 230.870 2063.000 231.190 ;
        RECT 2298.260 230.870 2298.520 231.190 ;
        RECT 2298.320 2.400 2298.460 230.870 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2071.910 472.500 2072.230 472.560 ;
        RECT 2311.570 472.500 2311.890 472.560 ;
        RECT 2071.910 472.360 2311.890 472.500 ;
        RECT 2071.910 472.300 2072.230 472.360 ;
        RECT 2311.570 472.300 2311.890 472.360 ;
      LAYER via ;
        RECT 2071.940 472.300 2072.200 472.560 ;
        RECT 2311.600 472.300 2311.860 472.560 ;
      LAYER met2 ;
        RECT 2072.070 510.340 2072.350 514.000 ;
        RECT 2072.000 510.000 2072.350 510.340 ;
        RECT 2072.000 472.590 2072.140 510.000 ;
        RECT 2071.940 472.270 2072.200 472.590 ;
        RECT 2311.600 472.270 2311.860 472.590 ;
        RECT 2311.660 17.410 2311.800 472.270 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2084.790 496.980 2085.110 497.040 ;
        RECT 2089.850 496.980 2090.170 497.040 ;
        RECT 2084.790 496.840 2090.170 496.980 ;
        RECT 2084.790 496.780 2085.110 496.840 ;
        RECT 2089.850 496.780 2090.170 496.840 ;
        RECT 2089.850 245.040 2090.170 245.100 ;
        RECT 2332.270 245.040 2332.590 245.100 ;
        RECT 2089.850 244.900 2332.590 245.040 ;
        RECT 2089.850 244.840 2090.170 244.900 ;
        RECT 2332.270 244.840 2332.590 244.900 ;
      LAYER via ;
        RECT 2084.820 496.780 2085.080 497.040 ;
        RECT 2089.880 496.780 2090.140 497.040 ;
        RECT 2089.880 244.840 2090.140 245.100 ;
        RECT 2332.300 244.840 2332.560 245.100 ;
      LAYER met2 ;
        RECT 2084.950 510.340 2085.230 514.000 ;
        RECT 2084.880 510.000 2085.230 510.340 ;
        RECT 2084.880 497.070 2085.020 510.000 ;
        RECT 2084.820 496.750 2085.080 497.070 ;
        RECT 2089.880 496.750 2090.140 497.070 ;
        RECT 2089.940 245.130 2090.080 496.750 ;
        RECT 2089.880 244.810 2090.140 245.130 ;
        RECT 2332.300 244.810 2332.560 245.130 ;
        RECT 2332.360 17.410 2332.500 244.810 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2097.210 252.180 2097.530 252.240 ;
        RECT 2346.070 252.180 2346.390 252.240 ;
        RECT 2097.210 252.040 2346.390 252.180 ;
        RECT 2097.210 251.980 2097.530 252.040 ;
        RECT 2346.070 251.980 2346.390 252.040 ;
      LAYER via ;
        RECT 2097.240 251.980 2097.500 252.240 ;
        RECT 2346.100 251.980 2346.360 252.240 ;
      LAYER met2 ;
        RECT 2097.370 510.340 2097.650 514.000 ;
        RECT 2097.300 510.000 2097.650 510.340 ;
        RECT 2097.300 252.270 2097.440 510.000 ;
        RECT 2097.240 251.950 2097.500 252.270 ;
        RECT 2346.100 251.950 2346.360 252.270 ;
        RECT 2346.160 17.410 2346.300 251.950 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2110.625 414.545 2110.795 462.315 ;
        RECT 2110.165 317.645 2110.335 406.895 ;
      LAYER mcon ;
        RECT 2110.625 462.145 2110.795 462.315 ;
        RECT 2110.165 406.725 2110.335 406.895 ;
      LAYER met1 ;
        RECT 2110.550 462.300 2110.870 462.360 ;
        RECT 2110.355 462.160 2110.870 462.300 ;
        RECT 2110.550 462.100 2110.870 462.160 ;
        RECT 2109.630 414.700 2109.950 414.760 ;
        RECT 2110.565 414.700 2110.855 414.745 ;
        RECT 2109.630 414.560 2110.855 414.700 ;
        RECT 2109.630 414.500 2109.950 414.560 ;
        RECT 2110.565 414.515 2110.855 414.560 ;
        RECT 2110.090 406.880 2110.410 406.940 ;
        RECT 2109.895 406.740 2110.410 406.880 ;
        RECT 2110.090 406.680 2110.410 406.740 ;
        RECT 2110.090 317.800 2110.410 317.860 ;
        RECT 2109.895 317.660 2110.410 317.800 ;
        RECT 2110.090 317.600 2110.410 317.660 ;
        RECT 2109.630 269.180 2109.950 269.240 ;
        RECT 2110.090 269.180 2110.410 269.240 ;
        RECT 2109.630 269.040 2110.410 269.180 ;
        RECT 2109.630 268.980 2109.950 269.040 ;
        RECT 2110.090 268.980 2110.410 269.040 ;
        RECT 2109.630 258.980 2109.950 259.040 ;
        RECT 2366.770 258.980 2367.090 259.040 ;
        RECT 2109.630 258.840 2367.090 258.980 ;
        RECT 2109.630 258.780 2109.950 258.840 ;
        RECT 2366.770 258.780 2367.090 258.840 ;
      LAYER via ;
        RECT 2110.580 462.100 2110.840 462.360 ;
        RECT 2109.660 414.500 2109.920 414.760 ;
        RECT 2110.120 406.680 2110.380 406.940 ;
        RECT 2110.120 317.600 2110.380 317.860 ;
        RECT 2109.660 268.980 2109.920 269.240 ;
        RECT 2110.120 268.980 2110.380 269.240 ;
        RECT 2109.660 258.780 2109.920 259.040 ;
        RECT 2366.800 258.780 2367.060 259.040 ;
      LAYER met2 ;
        RECT 2110.250 510.410 2110.530 514.000 ;
        RECT 2109.720 510.270 2110.530 510.410 ;
        RECT 2109.720 483.325 2109.860 510.270 ;
        RECT 2110.250 510.000 2110.530 510.270 ;
        RECT 2109.650 482.955 2109.930 483.325 ;
        RECT 2110.570 482.955 2110.850 483.325 ;
        RECT 2110.640 462.390 2110.780 482.955 ;
        RECT 2110.580 462.070 2110.840 462.390 ;
        RECT 2109.660 414.530 2109.920 414.790 ;
        RECT 2109.660 414.470 2110.320 414.530 ;
        RECT 2109.720 414.390 2110.320 414.470 ;
        RECT 2110.180 406.970 2110.320 414.390 ;
        RECT 2110.120 406.650 2110.380 406.970 ;
        RECT 2110.120 317.570 2110.380 317.890 ;
        RECT 2110.180 269.270 2110.320 317.570 ;
        RECT 2109.660 268.950 2109.920 269.270 ;
        RECT 2110.120 268.950 2110.380 269.270 ;
        RECT 2109.720 259.070 2109.860 268.950 ;
        RECT 2109.660 258.750 2109.920 259.070 ;
        RECT 2366.800 258.750 2367.060 259.070 ;
        RECT 2366.860 16.730 2367.000 258.750 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
      LAYER via2 ;
        RECT 2109.650 483.000 2109.930 483.280 ;
        RECT 2110.570 483.000 2110.850 483.280 ;
      LAYER met3 ;
        RECT 2109.625 483.290 2109.955 483.305 ;
        RECT 2110.545 483.290 2110.875 483.305 ;
        RECT 2109.625 482.990 2110.875 483.290 ;
        RECT 2109.625 482.975 2109.955 482.990 ;
        RECT 2110.545 482.975 2110.875 482.990 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.350 265.780 2124.670 265.840 ;
        RECT 2387.930 265.780 2388.250 265.840 ;
        RECT 2124.350 265.640 2388.250 265.780 ;
        RECT 2124.350 265.580 2124.670 265.640 ;
        RECT 2387.930 265.580 2388.250 265.640 ;
      LAYER via ;
        RECT 2124.380 265.580 2124.640 265.840 ;
        RECT 2387.960 265.580 2388.220 265.840 ;
      LAYER met2 ;
        RECT 2123.130 510.410 2123.410 514.000 ;
        RECT 2123.130 510.270 2124.580 510.410 ;
        RECT 2123.130 510.000 2123.410 510.270 ;
        RECT 2124.440 265.870 2124.580 510.270 ;
        RECT 2124.380 265.550 2124.640 265.870 ;
        RECT 2387.960 265.550 2388.220 265.870 ;
        RECT 2388.020 17.410 2388.160 265.550 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2135.850 497.320 2136.170 497.380 ;
        RECT 2156.090 497.320 2156.410 497.380 ;
        RECT 2135.850 497.180 2156.410 497.320 ;
        RECT 2135.850 497.120 2136.170 497.180 ;
        RECT 2156.090 497.120 2156.410 497.180 ;
        RECT 2156.090 272.580 2156.410 272.640 ;
        RECT 2401.270 272.580 2401.590 272.640 ;
        RECT 2156.090 272.440 2401.590 272.580 ;
        RECT 2156.090 272.380 2156.410 272.440 ;
        RECT 2401.270 272.380 2401.590 272.440 ;
      LAYER via ;
        RECT 2135.880 497.120 2136.140 497.380 ;
        RECT 2156.120 497.120 2156.380 497.380 ;
        RECT 2156.120 272.380 2156.380 272.640 ;
        RECT 2401.300 272.380 2401.560 272.640 ;
      LAYER met2 ;
        RECT 2136.010 510.340 2136.290 514.000 ;
        RECT 2135.940 510.000 2136.290 510.340 ;
        RECT 2135.940 497.410 2136.080 510.000 ;
        RECT 2135.880 497.090 2136.140 497.410 ;
        RECT 2156.120 497.090 2156.380 497.410 ;
        RECT 2156.180 272.670 2156.320 497.090 ;
        RECT 2156.120 272.350 2156.380 272.670 ;
        RECT 2401.300 272.350 2401.560 272.670 ;
        RECT 2401.360 16.730 2401.500 272.350 ;
        RECT 2401.360 16.590 2405.640 16.730 ;
        RECT 2405.500 2.400 2405.640 16.590 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 979.945 386.325 980.115 434.775 ;
      LAYER mcon ;
        RECT 979.945 434.605 980.115 434.775 ;
      LAYER met1 ;
        RECT 979.885 434.760 980.175 434.805 ;
        RECT 980.330 434.760 980.650 434.820 ;
        RECT 979.885 434.620 980.650 434.760 ;
        RECT 979.885 434.575 980.175 434.620 ;
        RECT 980.330 434.560 980.650 434.620 ;
        RECT 979.870 386.480 980.190 386.540 ;
        RECT 979.675 386.340 980.190 386.480 ;
        RECT 979.870 386.280 980.190 386.340 ;
        RECT 800.010 176.020 800.330 176.080 ;
        RECT 979.870 176.020 980.190 176.080 ;
        RECT 800.010 175.880 980.190 176.020 ;
        RECT 800.010 175.820 800.330 175.880 ;
        RECT 979.870 175.820 980.190 175.880 ;
      LAYER via ;
        RECT 980.360 434.560 980.620 434.820 ;
        RECT 979.900 386.280 980.160 386.540 ;
        RECT 800.040 175.820 800.300 176.080 ;
        RECT 979.900 175.820 980.160 176.080 ;
      LAYER met2 ;
        RECT 983.710 510.410 983.990 514.000 ;
        RECT 981.800 510.270 983.990 510.410 ;
        RECT 981.800 449.210 981.940 510.270 ;
        RECT 983.710 510.000 983.990 510.270 ;
        RECT 980.880 449.070 981.940 449.210 ;
        RECT 980.880 448.530 981.020 449.070 ;
        RECT 980.420 448.390 981.020 448.530 ;
        RECT 980.420 434.850 980.560 448.390 ;
        RECT 980.360 434.530 980.620 434.850 ;
        RECT 979.900 386.250 980.160 386.570 ;
        RECT 979.960 176.110 980.100 386.250 ;
        RECT 800.040 175.790 800.300 176.110 ;
        RECT 979.900 175.790 980.160 176.110 ;
        RECT 800.100 20.130 800.240 175.790 ;
        RECT 799.640 19.990 800.240 20.130 ;
        RECT 799.640 2.400 799.780 19.990 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 127.740 648.530 127.800 ;
        RECT 869.470 127.740 869.790 127.800 ;
        RECT 648.210 127.600 869.790 127.740 ;
        RECT 648.210 127.540 648.530 127.600 ;
        RECT 869.470 127.540 869.790 127.600 ;
        RECT 644.990 16.900 645.310 16.960 ;
        RECT 648.210 16.900 648.530 16.960 ;
        RECT 644.990 16.760 648.530 16.900 ;
        RECT 644.990 16.700 645.310 16.760 ;
        RECT 648.210 16.700 648.530 16.760 ;
      LAYER via ;
        RECT 648.240 127.540 648.500 127.800 ;
        RECT 869.500 127.540 869.760 127.800 ;
        RECT 645.020 16.700 645.280 16.960 ;
        RECT 648.240 16.700 648.500 16.960 ;
      LAYER met2 ;
        RECT 872.850 510.410 873.130 514.000 ;
        RECT 869.560 510.270 873.130 510.410 ;
        RECT 869.560 127.830 869.700 510.270 ;
        RECT 872.850 510.000 873.130 510.270 ;
        RECT 648.240 127.510 648.500 127.830 ;
        RECT 869.500 127.510 869.760 127.830 ;
        RECT 648.300 16.990 648.440 127.510 ;
        RECT 645.020 16.670 645.280 16.990 ;
        RECT 648.240 16.670 648.500 16.990 ;
        RECT 645.080 2.400 645.220 16.670 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.870 503.440 2153.190 503.500 ;
        RECT 2159.310 503.440 2159.630 503.500 ;
        RECT 2152.870 503.300 2159.630 503.440 ;
        RECT 2152.870 503.240 2153.190 503.300 ;
        RECT 2159.310 503.240 2159.630 503.300 ;
        RECT 2159.310 279.380 2159.630 279.440 ;
        RECT 2428.870 279.380 2429.190 279.440 ;
        RECT 2159.310 279.240 2429.190 279.380 ;
        RECT 2159.310 279.180 2159.630 279.240 ;
        RECT 2428.870 279.180 2429.190 279.240 ;
      LAYER via ;
        RECT 2152.900 503.240 2153.160 503.500 ;
        RECT 2159.340 503.240 2159.600 503.500 ;
        RECT 2159.340 279.180 2159.600 279.440 ;
        RECT 2428.900 279.180 2429.160 279.440 ;
      LAYER met2 ;
        RECT 2153.030 510.340 2153.310 514.000 ;
        RECT 2152.960 510.000 2153.310 510.340 ;
        RECT 2152.960 503.530 2153.100 510.000 ;
        RECT 2152.900 503.210 2153.160 503.530 ;
        RECT 2159.340 503.210 2159.600 503.530 ;
        RECT 2159.400 279.470 2159.540 503.210 ;
        RECT 2159.340 279.150 2159.600 279.470 ;
        RECT 2428.900 279.150 2429.160 279.470 ;
        RECT 2428.960 2.400 2429.100 279.150 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2165.290 400.420 2165.610 400.480 ;
        RECT 2166.210 400.420 2166.530 400.480 ;
        RECT 2165.290 400.280 2166.530 400.420 ;
        RECT 2165.290 400.220 2165.610 400.280 ;
        RECT 2166.210 400.220 2166.530 400.280 ;
        RECT 2166.210 286.180 2166.530 286.240 ;
        RECT 2442.670 286.180 2442.990 286.240 ;
        RECT 2166.210 286.040 2442.990 286.180 ;
        RECT 2166.210 285.980 2166.530 286.040 ;
        RECT 2442.670 285.980 2442.990 286.040 ;
      LAYER via ;
        RECT 2165.320 400.220 2165.580 400.480 ;
        RECT 2166.240 400.220 2166.500 400.480 ;
        RECT 2166.240 285.980 2166.500 286.240 ;
        RECT 2442.700 285.980 2442.960 286.240 ;
      LAYER met2 ;
        RECT 2165.910 510.410 2166.190 514.000 ;
        RECT 2165.380 510.270 2166.190 510.410 ;
        RECT 2165.380 483.325 2165.520 510.270 ;
        RECT 2165.910 510.000 2166.190 510.270 ;
        RECT 2165.310 482.955 2165.590 483.325 ;
        RECT 2166.230 482.955 2166.510 483.325 ;
        RECT 2166.300 448.530 2166.440 482.955 ;
        RECT 2165.380 448.390 2166.440 448.530 ;
        RECT 2165.380 400.510 2165.520 448.390 ;
        RECT 2166.300 400.510 2166.440 400.665 ;
        RECT 2165.320 400.250 2165.580 400.510 ;
        RECT 2166.240 400.250 2166.500 400.510 ;
        RECT 2165.320 400.190 2166.500 400.250 ;
        RECT 2165.380 400.110 2166.440 400.190 ;
        RECT 2165.380 351.970 2165.520 400.110 ;
        RECT 2165.380 351.830 2166.440 351.970 ;
        RECT 2166.300 286.270 2166.440 351.830 ;
        RECT 2166.240 285.950 2166.500 286.270 ;
        RECT 2442.700 285.950 2442.960 286.270 ;
        RECT 2442.760 16.730 2442.900 285.950 ;
        RECT 2442.760 16.590 2447.040 16.730 ;
        RECT 2446.900 2.400 2447.040 16.590 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
      LAYER via2 ;
        RECT 2165.310 483.000 2165.590 483.280 ;
        RECT 2166.230 483.000 2166.510 483.280 ;
      LAYER met3 ;
        RECT 2165.285 483.290 2165.615 483.305 ;
        RECT 2166.205 483.290 2166.535 483.305 ;
        RECT 2165.285 482.990 2166.535 483.290 ;
        RECT 2165.285 482.975 2165.615 482.990 ;
        RECT 2166.205 482.975 2166.535 482.990 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2179.550 293.320 2179.870 293.380 ;
        RECT 2463.370 293.320 2463.690 293.380 ;
        RECT 2179.550 293.180 2463.690 293.320 ;
        RECT 2179.550 293.120 2179.870 293.180 ;
        RECT 2463.370 293.120 2463.690 293.180 ;
      LAYER via ;
        RECT 2179.580 293.120 2179.840 293.380 ;
        RECT 2463.400 293.120 2463.660 293.380 ;
      LAYER met2 ;
        RECT 2178.790 510.410 2179.070 514.000 ;
        RECT 2178.790 510.270 2179.780 510.410 ;
        RECT 2178.790 510.000 2179.070 510.270 ;
        RECT 2179.640 293.410 2179.780 510.270 ;
        RECT 2179.580 293.090 2179.840 293.410 ;
        RECT 2463.400 293.090 2463.660 293.410 ;
        RECT 2463.460 17.410 2463.600 293.090 ;
        RECT 2463.460 17.270 2464.980 17.410 ;
        RECT 2464.840 2.400 2464.980 17.270 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2193.810 417.420 2194.130 417.480 ;
        RECT 2477.170 417.420 2477.490 417.480 ;
        RECT 2193.810 417.280 2477.490 417.420 ;
        RECT 2193.810 417.220 2194.130 417.280 ;
        RECT 2477.170 417.220 2477.490 417.280 ;
      LAYER via ;
        RECT 2193.840 417.220 2194.100 417.480 ;
        RECT 2477.200 417.220 2477.460 417.480 ;
      LAYER met2 ;
        RECT 2191.670 510.410 2191.950 514.000 ;
        RECT 2191.670 510.270 2194.040 510.410 ;
        RECT 2191.670 510.000 2191.950 510.270 ;
        RECT 2193.900 417.510 2194.040 510.270 ;
        RECT 2193.840 417.190 2194.100 417.510 ;
        RECT 2477.200 417.190 2477.460 417.510 ;
        RECT 2477.260 17.410 2477.400 417.190 ;
        RECT 2477.260 17.270 2482.920 17.410 ;
        RECT 2482.780 2.400 2482.920 17.270 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2207.610 300.120 2207.930 300.180 ;
        RECT 2497.870 300.120 2498.190 300.180 ;
        RECT 2207.610 299.980 2498.190 300.120 ;
        RECT 2207.610 299.920 2207.930 299.980 ;
        RECT 2497.870 299.920 2498.190 299.980 ;
      LAYER via ;
        RECT 2207.640 299.920 2207.900 300.180 ;
        RECT 2497.900 299.920 2498.160 300.180 ;
      LAYER met2 ;
        RECT 2204.090 510.410 2204.370 514.000 ;
        RECT 2204.090 510.270 2207.840 510.410 ;
        RECT 2204.090 510.000 2204.370 510.270 ;
        RECT 2207.700 300.210 2207.840 510.270 ;
        RECT 2207.640 299.890 2207.900 300.210 ;
        RECT 2497.900 299.890 2498.160 300.210 ;
        RECT 2497.960 16.730 2498.100 299.890 ;
        RECT 2497.960 16.590 2500.860 16.730 ;
        RECT 2500.720 2.400 2500.860 16.590 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2216.810 497.320 2217.130 497.380 ;
        RECT 2238.890 497.320 2239.210 497.380 ;
        RECT 2216.810 497.180 2239.210 497.320 ;
        RECT 2216.810 497.120 2217.130 497.180 ;
        RECT 2238.890 497.120 2239.210 497.180 ;
        RECT 2238.890 86.260 2239.210 86.320 ;
        RECT 2512.130 86.260 2512.450 86.320 ;
        RECT 2238.890 86.120 2512.450 86.260 ;
        RECT 2238.890 86.060 2239.210 86.120 ;
        RECT 2512.130 86.060 2512.450 86.120 ;
        RECT 2512.130 20.980 2512.450 21.040 ;
        RECT 2518.110 20.980 2518.430 21.040 ;
        RECT 2512.130 20.840 2518.430 20.980 ;
        RECT 2512.130 20.780 2512.450 20.840 ;
        RECT 2518.110 20.780 2518.430 20.840 ;
      LAYER via ;
        RECT 2216.840 497.120 2217.100 497.380 ;
        RECT 2238.920 497.120 2239.180 497.380 ;
        RECT 2238.920 86.060 2239.180 86.320 ;
        RECT 2512.160 86.060 2512.420 86.320 ;
        RECT 2512.160 20.780 2512.420 21.040 ;
        RECT 2518.140 20.780 2518.400 21.040 ;
      LAYER met2 ;
        RECT 2216.970 510.340 2217.250 514.000 ;
        RECT 2216.900 510.000 2217.250 510.340 ;
        RECT 2216.900 497.410 2217.040 510.000 ;
        RECT 2216.840 497.090 2217.100 497.410 ;
        RECT 2238.920 497.090 2239.180 497.410 ;
        RECT 2238.980 86.350 2239.120 497.090 ;
        RECT 2238.920 86.030 2239.180 86.350 ;
        RECT 2512.160 86.030 2512.420 86.350 ;
        RECT 2512.220 21.070 2512.360 86.030 ;
        RECT 2512.160 20.750 2512.420 21.070 ;
        RECT 2518.140 20.750 2518.400 21.070 ;
        RECT 2518.200 2.400 2518.340 20.750 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2229.690 503.440 2230.010 503.500 ;
        RECT 2234.750 503.440 2235.070 503.500 ;
        RECT 2229.690 503.300 2235.070 503.440 ;
        RECT 2229.690 503.240 2230.010 503.300 ;
        RECT 2234.750 503.240 2235.070 503.300 ;
        RECT 2234.750 306.920 2235.070 306.980 ;
        RECT 2532.370 306.920 2532.690 306.980 ;
        RECT 2234.750 306.780 2532.690 306.920 ;
        RECT 2234.750 306.720 2235.070 306.780 ;
        RECT 2532.370 306.720 2532.690 306.780 ;
      LAYER via ;
        RECT 2229.720 503.240 2229.980 503.500 ;
        RECT 2234.780 503.240 2235.040 503.500 ;
        RECT 2234.780 306.720 2235.040 306.980 ;
        RECT 2532.400 306.720 2532.660 306.980 ;
      LAYER met2 ;
        RECT 2229.850 510.340 2230.130 514.000 ;
        RECT 2229.780 510.000 2230.130 510.340 ;
        RECT 2229.780 503.530 2229.920 510.000 ;
        RECT 2229.720 503.210 2229.980 503.530 ;
        RECT 2234.780 503.210 2235.040 503.530 ;
        RECT 2234.840 307.010 2234.980 503.210 ;
        RECT 2234.780 306.690 2235.040 307.010 ;
        RECT 2532.400 306.690 2532.660 307.010 ;
        RECT 2532.460 16.730 2532.600 306.690 ;
        RECT 2532.460 16.590 2536.280 16.730 ;
        RECT 2536.140 2.400 2536.280 16.590 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.570 503.440 2242.890 503.500 ;
        RECT 2248.550 503.440 2248.870 503.500 ;
        RECT 2242.570 503.300 2248.870 503.440 ;
        RECT 2242.570 503.240 2242.890 503.300 ;
        RECT 2248.550 503.240 2248.870 503.300 ;
        RECT 2248.550 362.340 2248.870 362.400 ;
        RECT 2553.070 362.340 2553.390 362.400 ;
        RECT 2248.550 362.200 2553.390 362.340 ;
        RECT 2248.550 362.140 2248.870 362.200 ;
        RECT 2553.070 362.140 2553.390 362.200 ;
      LAYER via ;
        RECT 2242.600 503.240 2242.860 503.500 ;
        RECT 2248.580 503.240 2248.840 503.500 ;
        RECT 2248.580 362.140 2248.840 362.400 ;
        RECT 2553.100 362.140 2553.360 362.400 ;
      LAYER met2 ;
        RECT 2242.730 510.340 2243.010 514.000 ;
        RECT 2242.660 510.000 2243.010 510.340 ;
        RECT 2242.660 503.530 2242.800 510.000 ;
        RECT 2242.600 503.210 2242.860 503.530 ;
        RECT 2248.580 503.210 2248.840 503.530 ;
        RECT 2248.640 362.430 2248.780 503.210 ;
        RECT 2248.580 362.110 2248.840 362.430 ;
        RECT 2553.100 362.110 2553.360 362.430 ;
        RECT 2553.160 17.410 2553.300 362.110 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2254.990 448.700 2255.310 448.760 ;
        RECT 2255.910 448.700 2256.230 448.760 ;
        RECT 2254.990 448.560 2256.230 448.700 ;
        RECT 2254.990 448.500 2255.310 448.560 ;
        RECT 2255.910 448.500 2256.230 448.560 ;
        RECT 2254.990 355.200 2255.310 355.260 ;
        RECT 2566.870 355.200 2567.190 355.260 ;
        RECT 2254.990 355.060 2567.190 355.200 ;
        RECT 2254.990 355.000 2255.310 355.060 ;
        RECT 2566.870 355.000 2567.190 355.060 ;
      LAYER via ;
        RECT 2255.020 448.500 2255.280 448.760 ;
        RECT 2255.940 448.500 2256.200 448.760 ;
        RECT 2255.020 355.000 2255.280 355.260 ;
        RECT 2566.900 355.000 2567.160 355.260 ;
      LAYER met2 ;
        RECT 2255.610 510.410 2255.890 514.000 ;
        RECT 2255.080 510.270 2255.890 510.410 ;
        RECT 2255.080 483.325 2255.220 510.270 ;
        RECT 2255.610 510.000 2255.890 510.270 ;
        RECT 2255.010 482.955 2255.290 483.325 ;
        RECT 2255.930 482.955 2256.210 483.325 ;
        RECT 2256.000 448.790 2256.140 482.955 ;
        RECT 2255.020 448.470 2255.280 448.790 ;
        RECT 2255.940 448.470 2256.200 448.790 ;
        RECT 2255.080 355.290 2255.220 448.470 ;
        RECT 2255.020 354.970 2255.280 355.290 ;
        RECT 2566.900 354.970 2567.160 355.290 ;
        RECT 2566.960 17.410 2567.100 354.970 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.400 2572.160 17.270 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
      LAYER via2 ;
        RECT 2255.010 483.000 2255.290 483.280 ;
        RECT 2255.930 483.000 2256.210 483.280 ;
      LAYER met3 ;
        RECT 2254.985 483.290 2255.315 483.305 ;
        RECT 2255.905 483.290 2256.235 483.305 ;
        RECT 2254.985 482.990 2256.235 483.290 ;
        RECT 2254.985 482.975 2255.315 482.990 ;
        RECT 2255.905 482.975 2256.235 482.990 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 314.060 2270.030 314.120 ;
        RECT 2587.570 314.060 2587.890 314.120 ;
        RECT 2269.710 313.920 2587.890 314.060 ;
        RECT 2269.710 313.860 2270.030 313.920 ;
        RECT 2587.570 313.860 2587.890 313.920 ;
      LAYER via ;
        RECT 2269.740 313.860 2270.000 314.120 ;
        RECT 2587.600 313.860 2587.860 314.120 ;
      LAYER met2 ;
        RECT 2268.490 510.410 2268.770 514.000 ;
        RECT 2268.490 510.270 2269.940 510.410 ;
        RECT 2268.490 510.000 2268.770 510.270 ;
        RECT 2269.800 314.150 2269.940 510.270 ;
        RECT 2269.740 313.830 2270.000 314.150 ;
        RECT 2587.600 313.830 2587.860 314.150 ;
        RECT 2587.660 17.410 2587.800 313.830 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1001.565 386.325 1001.735 434.775 ;
      LAYER mcon ;
        RECT 1001.565 434.605 1001.735 434.775 ;
      LAYER met1 ;
        RECT 1001.490 434.760 1001.810 434.820 ;
        RECT 1001.295 434.620 1001.810 434.760 ;
        RECT 1001.490 434.560 1001.810 434.620 ;
        RECT 1001.490 386.480 1001.810 386.540 ;
        RECT 1001.295 386.340 1001.810 386.480 ;
        RECT 1001.490 386.280 1001.810 386.340 ;
        RECT 827.610 182.820 827.930 182.880 ;
        RECT 1001.490 182.820 1001.810 182.880 ;
        RECT 827.610 182.680 1001.810 182.820 ;
        RECT 827.610 182.620 827.930 182.680 ;
        RECT 1001.490 182.620 1001.810 182.680 ;
        RECT 823.470 17.580 823.790 17.640 ;
        RECT 827.610 17.580 827.930 17.640 ;
        RECT 823.470 17.440 827.930 17.580 ;
        RECT 823.470 17.380 823.790 17.440 ;
        RECT 827.610 17.380 827.930 17.440 ;
      LAYER via ;
        RECT 1001.520 434.560 1001.780 434.820 ;
        RECT 1001.520 386.280 1001.780 386.540 ;
        RECT 827.640 182.620 827.900 182.880 ;
        RECT 1001.520 182.620 1001.780 182.880 ;
        RECT 823.500 17.380 823.760 17.640 ;
        RECT 827.640 17.380 827.900 17.640 ;
      LAYER met2 ;
        RECT 1000.730 510.410 1001.010 514.000 ;
        RECT 1000.200 510.270 1001.010 510.410 ;
        RECT 1000.200 483.325 1000.340 510.270 ;
        RECT 1000.730 510.000 1001.010 510.270 ;
        RECT 1000.130 482.955 1000.410 483.325 ;
        RECT 1001.510 482.955 1001.790 483.325 ;
        RECT 1001.580 434.850 1001.720 482.955 ;
        RECT 1001.520 434.530 1001.780 434.850 ;
        RECT 1001.520 386.250 1001.780 386.570 ;
        RECT 1001.580 182.910 1001.720 386.250 ;
        RECT 827.640 182.590 827.900 182.910 ;
        RECT 1001.520 182.590 1001.780 182.910 ;
        RECT 827.700 17.670 827.840 182.590 ;
        RECT 823.500 17.350 823.760 17.670 ;
        RECT 827.640 17.350 827.900 17.670 ;
        RECT 823.560 2.400 823.700 17.350 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 1000.130 483.000 1000.410 483.280 ;
        RECT 1001.510 483.000 1001.790 483.280 ;
      LAYER met3 ;
        RECT 1000.105 483.290 1000.435 483.305 ;
        RECT 1001.485 483.290 1001.815 483.305 ;
        RECT 1000.105 482.990 1001.815 483.290 ;
        RECT 1000.105 482.975 1000.435 482.990 ;
        RECT 1001.485 482.975 1001.815 482.990 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2283.510 327.660 2283.830 327.720 ;
        RECT 2601.830 327.660 2602.150 327.720 ;
        RECT 2283.510 327.520 2602.150 327.660 ;
        RECT 2283.510 327.460 2283.830 327.520 ;
        RECT 2601.830 327.460 2602.150 327.520 ;
      LAYER via ;
        RECT 2283.540 327.460 2283.800 327.720 ;
        RECT 2601.860 327.460 2602.120 327.720 ;
      LAYER met2 ;
        RECT 2280.910 510.410 2281.190 514.000 ;
        RECT 2280.910 510.270 2283.740 510.410 ;
        RECT 2280.910 510.000 2281.190 510.270 ;
        RECT 2283.600 327.750 2283.740 510.270 ;
        RECT 2283.540 327.430 2283.800 327.750 ;
        RECT 2601.860 327.430 2602.120 327.750 ;
        RECT 2601.920 17.410 2602.060 327.430 ;
        RECT 2601.920 17.270 2607.580 17.410 ;
        RECT 2607.440 2.400 2607.580 17.270 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2293.630 496.980 2293.950 497.040 ;
        RECT 2297.310 496.980 2297.630 497.040 ;
        RECT 2293.630 496.840 2297.630 496.980 ;
        RECT 2293.630 496.780 2293.950 496.840 ;
        RECT 2297.310 496.780 2297.630 496.840 ;
        RECT 2297.310 348.400 2297.630 348.460 ;
        RECT 2622.070 348.400 2622.390 348.460 ;
        RECT 2297.310 348.260 2622.390 348.400 ;
        RECT 2297.310 348.200 2297.630 348.260 ;
        RECT 2622.070 348.200 2622.390 348.260 ;
      LAYER via ;
        RECT 2293.660 496.780 2293.920 497.040 ;
        RECT 2297.340 496.780 2297.600 497.040 ;
        RECT 2297.340 348.200 2297.600 348.460 ;
        RECT 2622.100 348.200 2622.360 348.460 ;
      LAYER met2 ;
        RECT 2293.790 510.340 2294.070 514.000 ;
        RECT 2293.720 510.000 2294.070 510.340 ;
        RECT 2293.720 497.070 2293.860 510.000 ;
        RECT 2293.660 496.750 2293.920 497.070 ;
        RECT 2297.340 496.750 2297.600 497.070 ;
        RECT 2297.400 348.490 2297.540 496.750 ;
        RECT 2297.340 348.170 2297.600 348.490 ;
        RECT 2622.100 348.170 2622.360 348.490 ;
        RECT 2622.160 17.410 2622.300 348.170 ;
        RECT 2622.160 17.270 2625.520 17.410 ;
        RECT 2625.380 2.400 2625.520 17.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2306.510 496.980 2306.830 497.040 ;
        RECT 2311.110 496.980 2311.430 497.040 ;
        RECT 2306.510 496.840 2311.430 496.980 ;
        RECT 2306.510 496.780 2306.830 496.840 ;
        RECT 2311.110 496.780 2311.430 496.840 ;
        RECT 2311.110 334.460 2311.430 334.520 ;
        RECT 2643.230 334.460 2643.550 334.520 ;
        RECT 2311.110 334.320 2643.550 334.460 ;
        RECT 2311.110 334.260 2311.430 334.320 ;
        RECT 2643.230 334.260 2643.550 334.320 ;
      LAYER via ;
        RECT 2306.540 496.780 2306.800 497.040 ;
        RECT 2311.140 496.780 2311.400 497.040 ;
        RECT 2311.140 334.260 2311.400 334.520 ;
        RECT 2643.260 334.260 2643.520 334.520 ;
      LAYER met2 ;
        RECT 2306.670 510.340 2306.950 514.000 ;
        RECT 2306.600 510.000 2306.950 510.340 ;
        RECT 2306.600 497.070 2306.740 510.000 ;
        RECT 2306.540 496.750 2306.800 497.070 ;
        RECT 2311.140 496.750 2311.400 497.070 ;
        RECT 2311.200 334.550 2311.340 496.750 ;
        RECT 2311.140 334.230 2311.400 334.550 ;
        RECT 2643.260 334.230 2643.520 334.550 ;
        RECT 2643.320 2.400 2643.460 334.230 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2319.390 496.980 2319.710 497.040 ;
        RECT 2324.450 496.980 2324.770 497.040 ;
        RECT 2319.390 496.840 2324.770 496.980 ;
        RECT 2319.390 496.780 2319.710 496.840 ;
        RECT 2324.450 496.780 2324.770 496.840 ;
        RECT 2324.450 341.600 2324.770 341.660 ;
        RECT 2656.570 341.600 2656.890 341.660 ;
        RECT 2324.450 341.460 2656.890 341.600 ;
        RECT 2324.450 341.400 2324.770 341.460 ;
        RECT 2656.570 341.400 2656.890 341.460 ;
      LAYER via ;
        RECT 2319.420 496.780 2319.680 497.040 ;
        RECT 2324.480 496.780 2324.740 497.040 ;
        RECT 2324.480 341.400 2324.740 341.660 ;
        RECT 2656.600 341.400 2656.860 341.660 ;
      LAYER met2 ;
        RECT 2319.550 510.340 2319.830 514.000 ;
        RECT 2319.480 510.000 2319.830 510.340 ;
        RECT 2319.480 497.070 2319.620 510.000 ;
        RECT 2319.420 496.750 2319.680 497.070 ;
        RECT 2324.480 496.750 2324.740 497.070 ;
        RECT 2324.540 341.690 2324.680 496.750 ;
        RECT 2324.480 341.370 2324.740 341.690 ;
        RECT 2656.600 341.370 2656.860 341.690 ;
        RECT 2656.660 17.410 2656.800 341.370 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2332.270 503.440 2332.590 503.500 ;
        RECT 2338.710 503.440 2339.030 503.500 ;
        RECT 2332.270 503.300 2339.030 503.440 ;
        RECT 2332.270 503.240 2332.590 503.300 ;
        RECT 2338.710 503.240 2339.030 503.300 ;
        RECT 2338.710 251.840 2339.030 251.900 ;
        RECT 2677.270 251.840 2677.590 251.900 ;
        RECT 2338.710 251.700 2677.590 251.840 ;
        RECT 2338.710 251.640 2339.030 251.700 ;
        RECT 2677.270 251.640 2677.590 251.700 ;
      LAYER via ;
        RECT 2332.300 503.240 2332.560 503.500 ;
        RECT 2338.740 503.240 2339.000 503.500 ;
        RECT 2338.740 251.640 2339.000 251.900 ;
        RECT 2677.300 251.640 2677.560 251.900 ;
      LAYER met2 ;
        RECT 2332.430 510.340 2332.710 514.000 ;
        RECT 2332.360 510.000 2332.710 510.340 ;
        RECT 2332.360 503.530 2332.500 510.000 ;
        RECT 2332.300 503.210 2332.560 503.530 ;
        RECT 2338.740 503.210 2339.000 503.530 ;
        RECT 2338.800 251.930 2338.940 503.210 ;
        RECT 2338.740 251.610 2339.000 251.930 ;
        RECT 2677.300 251.610 2677.560 251.930 ;
        RECT 2677.360 17.410 2677.500 251.610 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2344.305 448.205 2344.475 482.715 ;
        RECT 2344.765 338.045 2344.935 427.635 ;
      LAYER mcon ;
        RECT 2344.305 482.545 2344.475 482.715 ;
        RECT 2344.765 427.465 2344.935 427.635 ;
      LAYER met1 ;
        RECT 2343.770 483.380 2344.090 483.440 ;
        RECT 2344.230 483.380 2344.550 483.440 ;
        RECT 2343.770 483.240 2344.550 483.380 ;
        RECT 2343.770 483.180 2344.090 483.240 ;
        RECT 2344.230 483.180 2344.550 483.240 ;
        RECT 2344.230 482.700 2344.550 482.760 ;
        RECT 2344.035 482.560 2344.550 482.700 ;
        RECT 2344.230 482.500 2344.550 482.560 ;
        RECT 2344.245 448.360 2344.535 448.405 ;
        RECT 2345.150 448.360 2345.470 448.420 ;
        RECT 2344.245 448.220 2345.470 448.360 ;
        RECT 2344.245 448.175 2344.535 448.220 ;
        RECT 2345.150 448.160 2345.470 448.220 ;
        RECT 2344.705 427.620 2344.995 427.665 ;
        RECT 2345.150 427.620 2345.470 427.680 ;
        RECT 2344.705 427.480 2345.470 427.620 ;
        RECT 2344.705 427.435 2344.995 427.480 ;
        RECT 2345.150 427.420 2345.470 427.480 ;
        RECT 2344.690 338.200 2345.010 338.260 ;
        RECT 2344.495 338.060 2345.010 338.200 ;
        RECT 2344.690 338.000 2345.010 338.060 ;
        RECT 2345.610 258.640 2345.930 258.700 ;
        RECT 2691.070 258.640 2691.390 258.700 ;
        RECT 2345.610 258.500 2691.390 258.640 ;
        RECT 2345.610 258.440 2345.930 258.500 ;
        RECT 2691.070 258.440 2691.390 258.500 ;
      LAYER via ;
        RECT 2343.800 483.180 2344.060 483.440 ;
        RECT 2344.260 483.180 2344.520 483.440 ;
        RECT 2344.260 482.500 2344.520 482.760 ;
        RECT 2345.180 448.160 2345.440 448.420 ;
        RECT 2345.180 427.420 2345.440 427.680 ;
        RECT 2344.720 338.000 2344.980 338.260 ;
        RECT 2345.640 258.440 2345.900 258.700 ;
        RECT 2691.100 258.440 2691.360 258.700 ;
      LAYER met2 ;
        RECT 2345.310 511.090 2345.590 514.000 ;
        RECT 2343.860 510.950 2345.590 511.090 ;
        RECT 2343.860 483.470 2344.000 510.950 ;
        RECT 2345.310 510.000 2345.590 510.950 ;
        RECT 2343.800 483.150 2344.060 483.470 ;
        RECT 2344.260 483.150 2344.520 483.470 ;
        RECT 2344.320 482.790 2344.460 483.150 ;
        RECT 2344.260 482.470 2344.520 482.790 ;
        RECT 2345.180 448.130 2345.440 448.450 ;
        RECT 2345.240 427.710 2345.380 448.130 ;
        RECT 2345.180 427.390 2345.440 427.710 ;
        RECT 2344.720 337.970 2344.980 338.290 ;
        RECT 2344.780 303.690 2344.920 337.970 ;
        RECT 2344.780 303.550 2345.840 303.690 ;
        RECT 2345.700 258.730 2345.840 303.550 ;
        RECT 2345.640 258.410 2345.900 258.730 ;
        RECT 2691.100 258.410 2691.360 258.730 ;
        RECT 2691.160 16.730 2691.300 258.410 ;
        RECT 2691.160 16.590 2696.820 16.730 ;
        RECT 2696.680 2.400 2696.820 16.590 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2358.950 265.440 2359.270 265.500 ;
        RECT 2711.770 265.440 2712.090 265.500 ;
        RECT 2358.950 265.300 2712.090 265.440 ;
        RECT 2358.950 265.240 2359.270 265.300 ;
        RECT 2711.770 265.240 2712.090 265.300 ;
      LAYER via ;
        RECT 2358.980 265.240 2359.240 265.500 ;
        RECT 2711.800 265.240 2712.060 265.500 ;
      LAYER met2 ;
        RECT 2357.730 510.410 2358.010 514.000 ;
        RECT 2357.730 510.270 2359.180 510.410 ;
        RECT 2357.730 510.000 2358.010 510.270 ;
        RECT 2359.040 265.530 2359.180 510.270 ;
        RECT 2358.980 265.210 2359.240 265.530 ;
        RECT 2711.800 265.210 2712.060 265.530 ;
        RECT 2711.860 16.730 2712.000 265.210 ;
        RECT 2711.860 16.590 2714.760 16.730 ;
        RECT 2714.620 2.400 2714.760 16.590 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2373.210 20.640 2373.530 20.700 ;
        RECT 2732.470 20.640 2732.790 20.700 ;
        RECT 2373.210 20.500 2732.790 20.640 ;
        RECT 2373.210 20.440 2373.530 20.500 ;
        RECT 2732.470 20.440 2732.790 20.500 ;
      LAYER via ;
        RECT 2373.240 20.440 2373.500 20.700 ;
        RECT 2732.500 20.440 2732.760 20.700 ;
      LAYER met2 ;
        RECT 2370.610 510.410 2370.890 514.000 ;
        RECT 2370.610 510.270 2373.440 510.410 ;
        RECT 2370.610 510.000 2370.890 510.270 ;
        RECT 2373.300 20.730 2373.440 510.270 ;
        RECT 2373.240 20.410 2373.500 20.730 ;
        RECT 2732.500 20.410 2732.760 20.730 ;
        RECT 2732.560 2.400 2732.700 20.410 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.010 20.300 2387.330 20.360 ;
        RECT 2750.410 20.300 2750.730 20.360 ;
        RECT 2387.010 20.160 2750.730 20.300 ;
        RECT 2387.010 20.100 2387.330 20.160 ;
        RECT 2750.410 20.100 2750.730 20.160 ;
      LAYER via ;
        RECT 2387.040 20.100 2387.300 20.360 ;
        RECT 2750.440 20.100 2750.700 20.360 ;
      LAYER met2 ;
        RECT 2383.490 510.410 2383.770 514.000 ;
        RECT 2383.490 510.270 2387.240 510.410 ;
        RECT 2383.490 510.000 2383.770 510.270 ;
        RECT 2387.100 20.390 2387.240 510.270 ;
        RECT 2387.040 20.070 2387.300 20.390 ;
        RECT 2750.440 20.070 2750.700 20.390 ;
        RECT 2750.500 2.400 2750.640 20.070 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2396.210 496.980 2396.530 497.040 ;
        RECT 2400.810 496.980 2401.130 497.040 ;
        RECT 2396.210 496.840 2401.130 496.980 ;
        RECT 2396.210 496.780 2396.530 496.840 ;
        RECT 2400.810 496.780 2401.130 496.840 ;
        RECT 2400.810 19.960 2401.130 20.020 ;
        RECT 2767.890 19.960 2768.210 20.020 ;
        RECT 2400.810 19.820 2768.210 19.960 ;
        RECT 2400.810 19.760 2401.130 19.820 ;
        RECT 2767.890 19.760 2768.210 19.820 ;
      LAYER via ;
        RECT 2396.240 496.780 2396.500 497.040 ;
        RECT 2400.840 496.780 2401.100 497.040 ;
        RECT 2400.840 19.760 2401.100 20.020 ;
        RECT 2767.920 19.760 2768.180 20.020 ;
      LAYER met2 ;
        RECT 2396.370 510.340 2396.650 514.000 ;
        RECT 2396.300 510.000 2396.650 510.340 ;
        RECT 2396.300 497.070 2396.440 510.000 ;
        RECT 2396.240 496.750 2396.500 497.070 ;
        RECT 2400.840 496.750 2401.100 497.070 ;
        RECT 2400.900 20.050 2401.040 496.750 ;
        RECT 2400.840 19.730 2401.100 20.050 ;
        RECT 2767.920 19.730 2768.180 20.050 ;
        RECT 2767.980 2.400 2768.120 19.730 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 189.620 841.730 189.680 ;
        RECT 1007.930 189.620 1008.250 189.680 ;
        RECT 841.410 189.480 1008.250 189.620 ;
        RECT 841.410 189.420 841.730 189.480 ;
        RECT 1007.930 189.420 1008.250 189.480 ;
      LAYER via ;
        RECT 841.440 189.420 841.700 189.680 ;
        RECT 1007.960 189.420 1008.220 189.680 ;
      LAYER met2 ;
        RECT 1013.610 510.410 1013.890 514.000 ;
        RECT 1010.320 510.270 1013.890 510.410 ;
        RECT 1010.320 472.330 1010.460 510.270 ;
        RECT 1013.610 510.000 1013.890 510.270 ;
        RECT 1008.020 472.190 1010.460 472.330 ;
        RECT 1008.020 189.710 1008.160 472.190 ;
        RECT 841.440 189.390 841.700 189.710 ;
        RECT 1007.960 189.390 1008.220 189.710 ;
        RECT 841.500 20.130 841.640 189.390 ;
        RECT 841.040 19.990 841.640 20.130 ;
        RECT 841.040 2.400 841.180 19.990 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2409.090 496.980 2409.410 497.040 ;
        RECT 2414.610 496.980 2414.930 497.040 ;
        RECT 2409.090 496.840 2414.930 496.980 ;
        RECT 2409.090 496.780 2409.410 496.840 ;
        RECT 2414.610 496.780 2414.930 496.840 ;
        RECT 2414.610 19.620 2414.930 19.680 ;
        RECT 2785.830 19.620 2786.150 19.680 ;
        RECT 2414.610 19.480 2786.150 19.620 ;
        RECT 2414.610 19.420 2414.930 19.480 ;
        RECT 2785.830 19.420 2786.150 19.480 ;
      LAYER via ;
        RECT 2409.120 496.780 2409.380 497.040 ;
        RECT 2414.640 496.780 2414.900 497.040 ;
        RECT 2414.640 19.420 2414.900 19.680 ;
        RECT 2785.860 19.420 2786.120 19.680 ;
      LAYER met2 ;
        RECT 2409.250 510.340 2409.530 514.000 ;
        RECT 2409.180 510.000 2409.530 510.340 ;
        RECT 2409.180 497.070 2409.320 510.000 ;
        RECT 2409.120 496.750 2409.380 497.070 ;
        RECT 2414.640 496.750 2414.900 497.070 ;
        RECT 2414.700 19.710 2414.840 496.750 ;
        RECT 2414.640 19.390 2414.900 19.710 ;
        RECT 2785.860 19.390 2786.120 19.710 ;
        RECT 2785.920 2.400 2786.060 19.390 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2421.970 496.980 2422.290 497.040 ;
        RECT 2428.410 496.980 2428.730 497.040 ;
        RECT 2421.970 496.840 2428.730 496.980 ;
        RECT 2421.970 496.780 2422.290 496.840 ;
        RECT 2428.410 496.780 2428.730 496.840 ;
        RECT 2428.410 19.280 2428.730 19.340 ;
        RECT 2803.770 19.280 2804.090 19.340 ;
        RECT 2428.410 19.140 2804.090 19.280 ;
        RECT 2428.410 19.080 2428.730 19.140 ;
        RECT 2803.770 19.080 2804.090 19.140 ;
      LAYER via ;
        RECT 2422.000 496.780 2422.260 497.040 ;
        RECT 2428.440 496.780 2428.700 497.040 ;
        RECT 2428.440 19.080 2428.700 19.340 ;
        RECT 2803.800 19.080 2804.060 19.340 ;
      LAYER met2 ;
        RECT 2422.130 510.340 2422.410 514.000 ;
        RECT 2422.060 510.000 2422.410 510.340 ;
        RECT 2422.060 497.070 2422.200 510.000 ;
        RECT 2422.000 496.750 2422.260 497.070 ;
        RECT 2428.440 496.750 2428.700 497.070 ;
        RECT 2428.500 19.370 2428.640 496.750 ;
        RECT 2428.440 19.050 2428.700 19.370 ;
        RECT 2803.800 19.050 2804.060 19.370 ;
        RECT 2803.860 2.400 2804.000 19.050 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.310 18.940 2435.630 19.000 ;
        RECT 2821.710 18.940 2822.030 19.000 ;
        RECT 2435.310 18.800 2822.030 18.940 ;
        RECT 2435.310 18.740 2435.630 18.800 ;
        RECT 2821.710 18.740 2822.030 18.800 ;
      LAYER via ;
        RECT 2435.340 18.740 2435.600 19.000 ;
        RECT 2821.740 18.740 2822.000 19.000 ;
      LAYER met2 ;
        RECT 2434.550 510.410 2434.830 514.000 ;
        RECT 2434.550 510.270 2435.540 510.410 ;
        RECT 2434.550 510.000 2434.830 510.270 ;
        RECT 2435.400 19.030 2435.540 510.270 ;
        RECT 2435.340 18.710 2435.600 19.030 ;
        RECT 2821.740 18.710 2822.000 19.030 ;
        RECT 2821.800 2.400 2821.940 18.710 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2449.110 18.600 2449.430 18.660 ;
        RECT 2839.190 18.600 2839.510 18.660 ;
        RECT 2449.110 18.460 2839.510 18.600 ;
        RECT 2449.110 18.400 2449.430 18.460 ;
        RECT 2839.190 18.400 2839.510 18.460 ;
      LAYER via ;
        RECT 2449.140 18.400 2449.400 18.660 ;
        RECT 2839.220 18.400 2839.480 18.660 ;
      LAYER met2 ;
        RECT 2447.430 510.410 2447.710 514.000 ;
        RECT 2447.430 510.270 2449.340 510.410 ;
        RECT 2447.430 510.000 2447.710 510.270 ;
        RECT 2449.200 18.690 2449.340 510.270 ;
        RECT 2449.140 18.370 2449.400 18.690 ;
        RECT 2839.220 18.370 2839.480 18.690 ;
        RECT 2839.280 2.400 2839.420 18.370 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2462.910 18.260 2463.230 18.320 ;
        RECT 2856.670 18.260 2856.990 18.320 ;
        RECT 2462.910 18.120 2856.990 18.260 ;
        RECT 2462.910 18.060 2463.230 18.120 ;
        RECT 2856.670 18.060 2856.990 18.120 ;
      LAYER via ;
        RECT 2462.940 18.060 2463.200 18.320 ;
        RECT 2856.700 18.060 2856.960 18.320 ;
      LAYER met2 ;
        RECT 2460.310 510.410 2460.590 514.000 ;
        RECT 2460.310 510.270 2463.140 510.410 ;
        RECT 2460.310 510.000 2460.590 510.270 ;
        RECT 2463.000 18.350 2463.140 510.270 ;
        RECT 2462.940 18.030 2463.200 18.350 ;
        RECT 2856.700 18.030 2856.960 18.350 ;
        RECT 2856.760 17.410 2856.900 18.030 ;
        RECT 2856.760 17.270 2857.360 17.410 ;
        RECT 2857.220 2.400 2857.360 17.270 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2843.865 16.745 2844.035 17.935 ;
      LAYER mcon ;
        RECT 2843.865 17.765 2844.035 17.935 ;
      LAYER met1 ;
        RECT 2473.030 496.980 2473.350 497.040 ;
        RECT 2476.710 496.980 2477.030 497.040 ;
        RECT 2473.030 496.840 2477.030 496.980 ;
        RECT 2473.030 496.780 2473.350 496.840 ;
        RECT 2476.710 496.780 2477.030 496.840 ;
        RECT 2475.790 17.920 2476.110 17.980 ;
        RECT 2843.805 17.920 2844.095 17.965 ;
        RECT 2475.790 17.780 2844.095 17.920 ;
        RECT 2475.790 17.720 2476.110 17.780 ;
        RECT 2843.805 17.735 2844.095 17.780 ;
        RECT 2843.805 16.900 2844.095 16.945 ;
        RECT 2875.070 16.900 2875.390 16.960 ;
        RECT 2843.805 16.760 2875.390 16.900 ;
        RECT 2843.805 16.715 2844.095 16.760 ;
        RECT 2875.070 16.700 2875.390 16.760 ;
      LAYER via ;
        RECT 2473.060 496.780 2473.320 497.040 ;
        RECT 2476.740 496.780 2477.000 497.040 ;
        RECT 2475.820 17.720 2476.080 17.980 ;
        RECT 2875.100 16.700 2875.360 16.960 ;
      LAYER met2 ;
        RECT 2473.190 510.340 2473.470 514.000 ;
        RECT 2473.120 510.000 2473.470 510.340 ;
        RECT 2473.120 497.070 2473.260 510.000 ;
        RECT 2473.060 496.750 2473.320 497.070 ;
        RECT 2476.740 496.750 2477.000 497.070 ;
        RECT 2476.800 26.250 2476.940 496.750 ;
        RECT 2475.880 26.110 2476.940 26.250 ;
        RECT 2475.880 18.010 2476.020 26.110 ;
        RECT 2475.820 17.690 2476.080 18.010 ;
        RECT 2875.100 16.670 2875.360 16.990 ;
        RECT 2875.160 2.400 2875.300 16.670 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2485.910 496.980 2486.230 497.040 ;
        RECT 2490.510 496.980 2490.830 497.040 ;
        RECT 2485.910 496.840 2490.830 496.980 ;
        RECT 2485.910 496.780 2486.230 496.840 ;
        RECT 2490.510 496.780 2490.830 496.840 ;
        RECT 2490.510 17.580 2490.830 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2490.510 17.440 2893.330 17.580 ;
        RECT 2490.510 17.380 2490.830 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 2485.940 496.780 2486.200 497.040 ;
        RECT 2490.540 496.780 2490.800 497.040 ;
        RECT 2490.540 17.380 2490.800 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 2486.070 510.340 2486.350 514.000 ;
        RECT 2486.000 510.000 2486.350 510.340 ;
        RECT 2486.000 497.070 2486.140 510.000 ;
        RECT 2485.940 496.750 2486.200 497.070 ;
        RECT 2490.540 496.750 2490.800 497.070 ;
        RECT 2490.600 17.670 2490.740 496.750 ;
        RECT 2490.540 17.350 2490.800 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2498.790 496.980 2499.110 497.040 ;
        RECT 2504.310 496.980 2504.630 497.040 ;
        RECT 2498.790 496.840 2504.630 496.980 ;
        RECT 2498.790 496.780 2499.110 496.840 ;
        RECT 2504.310 496.780 2504.630 496.840 ;
        RECT 2504.310 17.240 2504.630 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2504.310 17.100 2911.270 17.240 ;
        RECT 2504.310 17.040 2504.630 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 2498.820 496.780 2499.080 497.040 ;
        RECT 2504.340 496.780 2504.600 497.040 ;
        RECT 2504.340 17.040 2504.600 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 2498.950 510.340 2499.230 514.000 ;
        RECT 2498.880 510.000 2499.230 510.340 ;
        RECT 2498.880 497.070 2499.020 510.000 ;
        RECT 2498.820 496.750 2499.080 497.070 ;
        RECT 2504.340 496.750 2504.600 497.070 ;
        RECT 2504.400 17.330 2504.540 496.750 ;
        RECT 2504.340 17.010 2504.600 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 17.240 859.210 17.300 ;
        RECT 1022.190 17.240 1022.510 17.300 ;
        RECT 858.890 17.100 1022.510 17.240 ;
        RECT 858.890 17.040 859.210 17.100 ;
        RECT 1022.190 17.040 1022.510 17.100 ;
      LAYER via ;
        RECT 858.920 17.040 859.180 17.300 ;
        RECT 1022.220 17.040 1022.480 17.300 ;
      LAYER met2 ;
        RECT 1026.490 510.410 1026.770 514.000 ;
        RECT 1022.740 510.270 1026.770 510.410 ;
        RECT 1022.740 449.210 1022.880 510.270 ;
        RECT 1026.490 510.000 1026.770 510.270 ;
        RECT 1022.280 449.070 1022.880 449.210 ;
        RECT 1022.280 17.330 1022.420 449.070 ;
        RECT 858.920 17.010 859.180 17.330 ;
        RECT 1022.220 17.010 1022.480 17.330 ;
        RECT 858.980 2.400 859.120 17.010 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1035.145 144.925 1035.315 193.035 ;
      LAYER mcon ;
        RECT 1035.145 192.865 1035.315 193.035 ;
      LAYER met1 ;
        RECT 1034.610 241.300 1034.930 241.360 ;
        RECT 1035.530 241.300 1035.850 241.360 ;
        RECT 1034.610 241.160 1035.850 241.300 ;
        RECT 1034.610 241.100 1034.930 241.160 ;
        RECT 1035.530 241.100 1035.850 241.160 ;
        RECT 1035.070 193.020 1035.390 193.080 ;
        RECT 1034.875 192.880 1035.390 193.020 ;
        RECT 1035.070 192.820 1035.390 192.880 ;
        RECT 1035.085 145.080 1035.375 145.125 ;
        RECT 1035.530 145.080 1035.850 145.140 ;
        RECT 1035.085 144.940 1035.850 145.080 ;
        RECT 1035.085 144.895 1035.375 144.940 ;
        RECT 1035.530 144.880 1035.850 144.940 ;
        RECT 1035.070 96.800 1035.390 96.860 ;
        RECT 1035.530 96.800 1035.850 96.860 ;
        RECT 1035.070 96.660 1035.850 96.800 ;
        RECT 1035.070 96.600 1035.390 96.660 ;
        RECT 1035.530 96.600 1035.850 96.660 ;
        RECT 876.830 17.920 877.150 17.980 ;
        RECT 1035.530 17.920 1035.850 17.980 ;
        RECT 876.830 17.780 1035.850 17.920 ;
        RECT 876.830 17.720 877.150 17.780 ;
        RECT 1035.530 17.720 1035.850 17.780 ;
      LAYER via ;
        RECT 1034.640 241.100 1034.900 241.360 ;
        RECT 1035.560 241.100 1035.820 241.360 ;
        RECT 1035.100 192.820 1035.360 193.080 ;
        RECT 1035.560 144.880 1035.820 145.140 ;
        RECT 1035.100 96.600 1035.360 96.860 ;
        RECT 1035.560 96.600 1035.820 96.860 ;
        RECT 876.860 17.720 877.120 17.980 ;
        RECT 1035.560 17.720 1035.820 17.980 ;
      LAYER met2 ;
        RECT 1038.910 510.340 1039.190 514.000 ;
        RECT 1038.840 510.000 1039.190 510.340 ;
        RECT 1038.840 483.325 1038.980 510.000 ;
        RECT 1036.470 482.955 1036.750 483.325 ;
        RECT 1038.770 482.955 1039.050 483.325 ;
        RECT 1036.540 434.930 1036.680 482.955 ;
        RECT 1036.080 434.790 1036.680 434.930 ;
        RECT 1036.080 386.765 1036.220 434.790 ;
        RECT 1035.090 386.395 1035.370 386.765 ;
        RECT 1036.010 386.395 1036.290 386.765 ;
        RECT 1035.160 355.370 1035.300 386.395 ;
        RECT 1035.160 355.230 1036.220 355.370 ;
        RECT 1036.080 265.610 1036.220 355.230 ;
        RECT 1035.620 265.470 1036.220 265.610 ;
        RECT 1035.620 241.390 1035.760 265.470 ;
        RECT 1034.640 241.070 1034.900 241.390 ;
        RECT 1035.560 241.070 1035.820 241.390 ;
        RECT 1034.700 193.530 1034.840 241.070 ;
        RECT 1034.700 193.390 1035.300 193.530 ;
        RECT 1035.160 193.110 1035.300 193.390 ;
        RECT 1035.100 192.790 1035.360 193.110 ;
        RECT 1035.560 144.850 1035.820 145.170 ;
        RECT 1035.620 96.890 1035.760 144.850 ;
        RECT 1035.100 96.570 1035.360 96.890 ;
        RECT 1035.560 96.570 1035.820 96.890 ;
        RECT 1035.160 48.010 1035.300 96.570 ;
        RECT 1035.160 47.870 1035.760 48.010 ;
        RECT 1035.620 18.010 1035.760 47.870 ;
        RECT 876.860 17.690 877.120 18.010 ;
        RECT 1035.560 17.690 1035.820 18.010 ;
        RECT 876.920 2.400 877.060 17.690 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1036.470 483.000 1036.750 483.280 ;
        RECT 1038.770 483.000 1039.050 483.280 ;
        RECT 1035.090 386.440 1035.370 386.720 ;
        RECT 1036.010 386.440 1036.290 386.720 ;
      LAYER met3 ;
        RECT 1036.445 483.290 1036.775 483.305 ;
        RECT 1038.745 483.290 1039.075 483.305 ;
        RECT 1036.445 482.990 1039.075 483.290 ;
        RECT 1036.445 482.975 1036.775 482.990 ;
        RECT 1038.745 482.975 1039.075 482.990 ;
        RECT 1035.065 386.730 1035.395 386.745 ;
        RECT 1035.985 386.730 1036.315 386.745 ;
        RECT 1035.065 386.430 1036.315 386.730 ;
        RECT 1035.065 386.415 1035.395 386.430 ;
        RECT 1035.985 386.415 1036.315 386.430 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 17.580 895.090 17.640 ;
        RECT 1049.790 17.580 1050.110 17.640 ;
        RECT 894.770 17.440 1050.110 17.580 ;
        RECT 894.770 17.380 895.090 17.440 ;
        RECT 1049.790 17.380 1050.110 17.440 ;
      LAYER via ;
        RECT 894.800 17.380 895.060 17.640 ;
        RECT 1049.820 17.380 1050.080 17.640 ;
      LAYER met2 ;
        RECT 1051.790 510.410 1052.070 514.000 ;
        RECT 1049.880 510.270 1052.070 510.410 ;
        RECT 1049.880 17.670 1050.020 510.270 ;
        RECT 1051.790 510.000 1052.070 510.270 ;
        RECT 894.800 17.350 895.060 17.670 ;
        RECT 1049.820 17.350 1050.080 17.670 ;
        RECT 894.860 2.400 895.000 17.350 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 18.260 913.030 18.320 ;
        RECT 1062.670 18.260 1062.990 18.320 ;
        RECT 912.710 18.120 1062.990 18.260 ;
        RECT 912.710 18.060 913.030 18.120 ;
        RECT 1062.670 18.060 1062.990 18.120 ;
      LAYER via ;
        RECT 912.740 18.060 913.000 18.320 ;
        RECT 1062.700 18.060 1062.960 18.320 ;
      LAYER met2 ;
        RECT 1064.670 510.410 1064.950 514.000 ;
        RECT 1062.760 510.270 1064.950 510.410 ;
        RECT 1062.760 18.350 1062.900 510.270 ;
        RECT 1064.670 510.000 1064.950 510.270 ;
        RECT 912.740 18.030 913.000 18.350 ;
        RECT 1062.700 18.030 1062.960 18.350 ;
        RECT 912.800 2.400 912.940 18.030 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 930.190 18.600 930.510 18.660 ;
        RECT 1076.470 18.600 1076.790 18.660 ;
        RECT 930.190 18.460 1076.790 18.600 ;
        RECT 930.190 18.400 930.510 18.460 ;
        RECT 1076.470 18.400 1076.790 18.460 ;
      LAYER via ;
        RECT 930.220 18.400 930.480 18.660 ;
        RECT 1076.500 18.400 1076.760 18.660 ;
      LAYER met2 ;
        RECT 1077.550 510.410 1077.830 514.000 ;
        RECT 1076.560 510.270 1077.830 510.410 ;
        RECT 1076.560 18.690 1076.700 510.270 ;
        RECT 1077.550 510.000 1077.830 510.270 ;
        RECT 930.220 18.370 930.480 18.690 ;
        RECT 1076.500 18.370 1076.760 18.690 ;
        RECT 930.280 2.400 930.420 18.370 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 18.940 948.450 19.000 ;
        RECT 1090.270 18.940 1090.590 19.000 ;
        RECT 948.130 18.800 1090.590 18.940 ;
        RECT 948.130 18.740 948.450 18.800 ;
        RECT 1090.270 18.740 1090.590 18.800 ;
      LAYER via ;
        RECT 948.160 18.740 948.420 19.000 ;
        RECT 1090.300 18.740 1090.560 19.000 ;
      LAYER met2 ;
        RECT 1090.430 510.340 1090.710 514.000 ;
        RECT 1090.360 510.000 1090.710 510.340 ;
        RECT 1090.360 19.030 1090.500 510.000 ;
        RECT 948.160 18.710 948.420 19.030 ;
        RECT 1090.300 18.710 1090.560 19.030 ;
        RECT 948.220 2.400 948.360 18.710 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1098.090 193.840 1098.410 194.100 ;
        RECT 1098.180 193.420 1098.320 193.840 ;
        RECT 1098.090 193.160 1098.410 193.420 ;
        RECT 1098.090 158.820 1098.410 159.080 ;
        RECT 1098.180 158.340 1098.320 158.820 ;
        RECT 1098.550 158.340 1098.870 158.400 ;
        RECT 1098.180 158.200 1098.870 158.340 ;
        RECT 1098.550 158.140 1098.870 158.200 ;
        RECT 966.070 19.620 966.390 19.680 ;
        RECT 1097.630 19.620 1097.950 19.680 ;
        RECT 966.070 19.480 1097.950 19.620 ;
        RECT 966.070 19.420 966.390 19.480 ;
        RECT 1097.630 19.420 1097.950 19.480 ;
      LAYER via ;
        RECT 1098.120 193.840 1098.380 194.100 ;
        RECT 1098.120 193.160 1098.380 193.420 ;
        RECT 1098.120 158.820 1098.380 159.080 ;
        RECT 1098.580 158.140 1098.840 158.400 ;
        RECT 966.100 19.420 966.360 19.680 ;
        RECT 1097.660 19.420 1097.920 19.680 ;
      LAYER met2 ;
        RECT 1103.310 510.410 1103.590 514.000 ;
        RECT 1101.400 510.270 1103.590 510.410 ;
        RECT 1101.400 472.330 1101.540 510.270 ;
        RECT 1103.310 510.000 1103.590 510.270 ;
        RECT 1098.180 472.190 1101.540 472.330 ;
        RECT 1098.180 303.690 1098.320 472.190 ;
        RECT 1097.720 303.550 1098.320 303.690 ;
        RECT 1097.720 303.010 1097.860 303.550 ;
        RECT 1097.720 302.870 1098.320 303.010 ;
        RECT 1098.180 194.130 1098.320 302.870 ;
        RECT 1098.120 193.810 1098.380 194.130 ;
        RECT 1098.120 193.130 1098.380 193.450 ;
        RECT 1098.180 159.110 1098.320 193.130 ;
        RECT 1098.120 158.790 1098.380 159.110 ;
        RECT 1098.580 158.110 1098.840 158.430 ;
        RECT 1098.640 110.570 1098.780 158.110 ;
        RECT 1097.720 110.430 1098.780 110.570 ;
        RECT 1097.720 19.710 1097.860 110.430 ;
        RECT 966.100 19.390 966.360 19.710 ;
        RECT 1097.660 19.390 1097.920 19.710 ;
        RECT 966.160 2.400 966.300 19.390 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 472.840 1111.290 472.900 ;
        RECT 1114.190 472.840 1114.510 472.900 ;
        RECT 1110.970 472.700 1114.510 472.840 ;
        RECT 1110.970 472.640 1111.290 472.700 ;
        RECT 1114.190 472.640 1114.510 472.700 ;
        RECT 984.010 19.280 984.330 19.340 ;
        RECT 1110.970 19.280 1111.290 19.340 ;
        RECT 984.010 19.140 1111.290 19.280 ;
        RECT 984.010 19.080 984.330 19.140 ;
        RECT 1110.970 19.080 1111.290 19.140 ;
      LAYER via ;
        RECT 1111.000 472.640 1111.260 472.900 ;
        RECT 1114.220 472.640 1114.480 472.900 ;
        RECT 984.040 19.080 984.300 19.340 ;
        RECT 1111.000 19.080 1111.260 19.340 ;
      LAYER met2 ;
        RECT 1115.730 510.410 1116.010 514.000 ;
        RECT 1114.280 510.270 1116.010 510.410 ;
        RECT 1114.280 472.930 1114.420 510.270 ;
        RECT 1115.730 510.000 1116.010 510.270 ;
        RECT 1111.000 472.610 1111.260 472.930 ;
        RECT 1114.220 472.610 1114.480 472.930 ;
        RECT 1111.060 19.370 1111.200 472.610 ;
        RECT 984.040 19.050 984.300 19.370 ;
        RECT 1111.000 19.050 1111.260 19.370 ;
        RECT 984.100 2.400 984.240 19.050 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.990 500.040 714.310 500.100 ;
        RECT 885.110 500.040 885.430 500.100 ;
        RECT 713.990 499.900 885.430 500.040 ;
        RECT 713.990 499.840 714.310 499.900 ;
        RECT 885.110 499.840 885.430 499.900 ;
        RECT 662.930 31.180 663.250 31.240 ;
        RECT 713.990 31.180 714.310 31.240 ;
        RECT 662.930 31.040 714.310 31.180 ;
        RECT 662.930 30.980 663.250 31.040 ;
        RECT 713.990 30.980 714.310 31.040 ;
      LAYER via ;
        RECT 714.020 499.840 714.280 500.100 ;
        RECT 885.140 499.840 885.400 500.100 ;
        RECT 662.960 30.980 663.220 31.240 ;
        RECT 714.020 30.980 714.280 31.240 ;
      LAYER met2 ;
        RECT 885.270 510.340 885.550 514.000 ;
        RECT 885.200 510.000 885.550 510.340 ;
        RECT 885.200 500.130 885.340 510.000 ;
        RECT 714.020 499.810 714.280 500.130 ;
        RECT 885.140 499.810 885.400 500.130 ;
        RECT 714.080 31.270 714.220 499.810 ;
        RECT 662.960 30.950 663.220 31.270 ;
        RECT 714.020 30.950 714.280 31.270 ;
        RECT 663.020 2.400 663.160 30.950 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1124.385 379.525 1124.555 427.635 ;
        RECT 1124.845 186.405 1125.015 234.515 ;
        RECT 1124.845 96.985 1125.015 144.755 ;
        RECT 1124.845 48.365 1125.015 96.475 ;
      LAYER mcon ;
        RECT 1124.385 427.465 1124.555 427.635 ;
        RECT 1124.845 234.345 1125.015 234.515 ;
        RECT 1124.845 144.585 1125.015 144.755 ;
        RECT 1124.845 96.305 1125.015 96.475 ;
      LAYER met1 ;
        RECT 1124.310 435.100 1124.630 435.160 ;
        RECT 1126.610 435.100 1126.930 435.160 ;
        RECT 1124.310 434.960 1126.930 435.100 ;
        RECT 1124.310 434.900 1124.630 434.960 ;
        RECT 1126.610 434.900 1126.930 434.960 ;
        RECT 1124.310 427.620 1124.630 427.680 ;
        RECT 1124.115 427.480 1124.630 427.620 ;
        RECT 1124.310 427.420 1124.630 427.480 ;
        RECT 1124.325 379.680 1124.615 379.725 ;
        RECT 1124.770 379.680 1125.090 379.740 ;
        RECT 1124.325 379.540 1125.090 379.680 ;
        RECT 1124.325 379.495 1124.615 379.540 ;
        RECT 1124.770 379.480 1125.090 379.540 ;
        RECT 1124.310 299.440 1124.630 299.500 ;
        RECT 1125.230 299.440 1125.550 299.500 ;
        RECT 1124.310 299.300 1125.550 299.440 ;
        RECT 1124.310 299.240 1124.630 299.300 ;
        RECT 1125.230 299.240 1125.550 299.300 ;
        RECT 1124.770 241.300 1125.090 241.360 ;
        RECT 1125.230 241.300 1125.550 241.360 ;
        RECT 1124.770 241.160 1125.550 241.300 ;
        RECT 1124.770 241.100 1125.090 241.160 ;
        RECT 1125.230 241.100 1125.550 241.160 ;
        RECT 1124.770 234.500 1125.090 234.560 ;
        RECT 1124.575 234.360 1125.090 234.500 ;
        RECT 1124.770 234.300 1125.090 234.360 ;
        RECT 1124.770 186.560 1125.090 186.620 ;
        RECT 1124.575 186.420 1125.090 186.560 ;
        RECT 1124.770 186.360 1125.090 186.420 ;
        RECT 1124.770 158.820 1125.090 159.080 ;
        RECT 1124.860 158.400 1125.000 158.820 ;
        RECT 1124.770 158.140 1125.090 158.400 ;
        RECT 1124.770 144.740 1125.090 144.800 ;
        RECT 1124.575 144.600 1125.090 144.740 ;
        RECT 1124.770 144.540 1125.090 144.600 ;
        RECT 1124.770 97.140 1125.090 97.200 ;
        RECT 1124.575 97.000 1125.090 97.140 ;
        RECT 1124.770 96.940 1125.090 97.000 ;
        RECT 1124.770 96.460 1125.090 96.520 ;
        RECT 1124.575 96.320 1125.090 96.460 ;
        RECT 1124.770 96.260 1125.090 96.320 ;
        RECT 1124.785 48.520 1125.075 48.565 ;
        RECT 1125.230 48.520 1125.550 48.580 ;
        RECT 1124.785 48.380 1125.550 48.520 ;
        RECT 1124.785 48.335 1125.075 48.380 ;
        RECT 1125.230 48.320 1125.550 48.380 ;
        RECT 1001.950 20.300 1002.270 20.360 ;
        RECT 1125.230 20.300 1125.550 20.360 ;
        RECT 1001.950 20.160 1125.550 20.300 ;
        RECT 1001.950 20.100 1002.270 20.160 ;
        RECT 1125.230 20.100 1125.550 20.160 ;
      LAYER via ;
        RECT 1124.340 434.900 1124.600 435.160 ;
        RECT 1126.640 434.900 1126.900 435.160 ;
        RECT 1124.340 427.420 1124.600 427.680 ;
        RECT 1124.800 379.480 1125.060 379.740 ;
        RECT 1124.340 299.240 1124.600 299.500 ;
        RECT 1125.260 299.240 1125.520 299.500 ;
        RECT 1124.800 241.100 1125.060 241.360 ;
        RECT 1125.260 241.100 1125.520 241.360 ;
        RECT 1124.800 234.300 1125.060 234.560 ;
        RECT 1124.800 186.360 1125.060 186.620 ;
        RECT 1124.800 158.820 1125.060 159.080 ;
        RECT 1124.800 158.140 1125.060 158.400 ;
        RECT 1124.800 144.540 1125.060 144.800 ;
        RECT 1124.800 96.940 1125.060 97.200 ;
        RECT 1124.800 96.260 1125.060 96.520 ;
        RECT 1125.260 48.320 1125.520 48.580 ;
        RECT 1001.980 20.100 1002.240 20.360 ;
        RECT 1125.260 20.100 1125.520 20.360 ;
      LAYER met2 ;
        RECT 1128.610 510.410 1128.890 514.000 ;
        RECT 1126.700 510.270 1128.890 510.410 ;
        RECT 1126.700 435.190 1126.840 510.270 ;
        RECT 1128.610 510.000 1128.890 510.270 ;
        RECT 1124.340 434.870 1124.600 435.190 ;
        RECT 1126.640 434.870 1126.900 435.190 ;
        RECT 1124.400 427.710 1124.540 434.870 ;
        RECT 1124.340 427.390 1124.600 427.710 ;
        RECT 1124.800 379.450 1125.060 379.770 ;
        RECT 1124.860 379.170 1125.000 379.450 ;
        RECT 1124.400 379.030 1125.000 379.170 ;
        RECT 1124.400 337.690 1124.540 379.030 ;
        RECT 1124.400 337.550 1125.460 337.690 ;
        RECT 1125.320 299.530 1125.460 337.550 ;
        RECT 1124.340 299.210 1124.600 299.530 ;
        RECT 1125.260 299.210 1125.520 299.530 ;
        RECT 1124.400 264.930 1124.540 299.210 ;
        RECT 1124.400 264.790 1125.460 264.930 ;
        RECT 1125.320 241.390 1125.460 264.790 ;
        RECT 1124.800 241.070 1125.060 241.390 ;
        RECT 1125.260 241.070 1125.520 241.390 ;
        RECT 1124.860 234.590 1125.000 241.070 ;
        RECT 1124.800 234.270 1125.060 234.590 ;
        RECT 1124.800 186.330 1125.060 186.650 ;
        RECT 1124.860 159.110 1125.000 186.330 ;
        RECT 1124.800 158.790 1125.060 159.110 ;
        RECT 1124.800 158.110 1125.060 158.430 ;
        RECT 1124.860 144.830 1125.000 158.110 ;
        RECT 1124.800 144.510 1125.060 144.830 ;
        RECT 1124.800 96.910 1125.060 97.230 ;
        RECT 1124.860 96.550 1125.000 96.910 ;
        RECT 1124.800 96.230 1125.060 96.550 ;
        RECT 1125.260 48.290 1125.520 48.610 ;
        RECT 1125.320 20.390 1125.460 48.290 ;
        RECT 1001.980 20.070 1002.240 20.390 ;
        RECT 1125.260 20.070 1125.520 20.390 ;
        RECT 1002.040 2.400 1002.180 20.070 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.430 19.960 1019.750 20.020 ;
        RECT 1138.570 19.960 1138.890 20.020 ;
        RECT 1019.430 19.820 1138.890 19.960 ;
        RECT 1019.430 19.760 1019.750 19.820 ;
        RECT 1138.570 19.760 1138.890 19.820 ;
      LAYER via ;
        RECT 1019.460 19.760 1019.720 20.020 ;
        RECT 1138.600 19.760 1138.860 20.020 ;
      LAYER met2 ;
        RECT 1141.490 510.410 1141.770 514.000 ;
        RECT 1138.660 510.270 1141.770 510.410 ;
        RECT 1138.660 20.050 1138.800 510.270 ;
        RECT 1141.490 510.000 1141.770 510.270 ;
        RECT 1019.460 19.730 1019.720 20.050 ;
        RECT 1138.600 19.730 1138.860 20.050 ;
        RECT 1019.520 2.400 1019.660 19.730 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 17.920 1037.690 17.980 ;
        RECT 1152.370 17.920 1152.690 17.980 ;
        RECT 1037.370 17.780 1152.690 17.920 ;
        RECT 1037.370 17.720 1037.690 17.780 ;
        RECT 1152.370 17.720 1152.690 17.780 ;
      LAYER via ;
        RECT 1037.400 17.720 1037.660 17.980 ;
        RECT 1152.400 17.720 1152.660 17.980 ;
      LAYER met2 ;
        RECT 1154.370 510.410 1154.650 514.000 ;
        RECT 1152.460 510.270 1154.650 510.410 ;
        RECT 1152.460 18.010 1152.600 510.270 ;
        RECT 1154.370 510.000 1154.650 510.270 ;
        RECT 1037.400 17.690 1037.660 18.010 ;
        RECT 1152.400 17.690 1152.660 18.010 ;
        RECT 1037.460 2.400 1037.600 17.690 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 17.240 1167.410 17.300 ;
        RECT 1059.080 17.100 1167.410 17.240 ;
        RECT 1059.080 16.900 1059.220 17.100 ;
        RECT 1167.090 17.040 1167.410 17.100 ;
        RECT 1055.400 16.760 1059.220 16.900 ;
        RECT 1055.400 16.620 1055.540 16.760 ;
        RECT 1055.310 16.360 1055.630 16.620 ;
      LAYER via ;
        RECT 1167.120 17.040 1167.380 17.300 ;
        RECT 1055.340 16.360 1055.600 16.620 ;
      LAYER met2 ;
        RECT 1167.250 510.340 1167.530 514.000 ;
        RECT 1167.180 510.000 1167.530 510.340 ;
        RECT 1167.180 17.330 1167.320 510.000 ;
        RECT 1167.120 17.010 1167.380 17.330 ;
        RECT 1055.340 16.330 1055.600 16.650 ;
        RECT 1055.400 2.400 1055.540 16.330 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1124.385 16.405 1124.555 17.595 ;
        RECT 1124.845 16.405 1125.015 17.595 ;
        RECT 1167.625 16.405 1167.795 17.255 ;
      LAYER mcon ;
        RECT 1124.385 17.425 1124.555 17.595 ;
        RECT 1124.845 17.425 1125.015 17.595 ;
        RECT 1167.625 17.085 1167.795 17.255 ;
      LAYER met1 ;
        RECT 1124.325 17.580 1124.615 17.625 ;
        RECT 1124.785 17.580 1125.075 17.625 ;
        RECT 1180.890 17.580 1181.210 17.640 ;
        RECT 1124.325 17.440 1125.075 17.580 ;
        RECT 1124.325 17.395 1124.615 17.440 ;
        RECT 1124.785 17.395 1125.075 17.440 ;
        RECT 1173.620 17.440 1181.210 17.580 ;
        RECT 1167.565 17.240 1167.855 17.285 ;
        RECT 1173.620 17.240 1173.760 17.440 ;
        RECT 1180.890 17.380 1181.210 17.440 ;
        RECT 1167.565 17.100 1173.760 17.240 ;
        RECT 1167.565 17.055 1167.855 17.100 ;
        RECT 1073.250 16.560 1073.570 16.620 ;
        RECT 1124.325 16.560 1124.615 16.605 ;
        RECT 1073.250 16.420 1124.615 16.560 ;
        RECT 1073.250 16.360 1073.570 16.420 ;
        RECT 1124.325 16.375 1124.615 16.420 ;
        RECT 1124.785 16.560 1125.075 16.605 ;
        RECT 1167.565 16.560 1167.855 16.605 ;
        RECT 1124.785 16.420 1167.855 16.560 ;
        RECT 1124.785 16.375 1125.075 16.420 ;
        RECT 1167.565 16.375 1167.855 16.420 ;
      LAYER via ;
        RECT 1180.920 17.380 1181.180 17.640 ;
        RECT 1073.280 16.360 1073.540 16.620 ;
      LAYER met2 ;
        RECT 1180.130 510.410 1180.410 514.000 ;
        RECT 1180.130 510.270 1181.120 510.410 ;
        RECT 1180.130 510.000 1180.410 510.270 ;
        RECT 1180.980 17.670 1181.120 510.270 ;
        RECT 1180.920 17.350 1181.180 17.670 ;
        RECT 1073.280 16.330 1073.540 16.650 ;
        RECT 1073.340 2.400 1073.480 16.330 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.870 472.840 1187.190 472.900 ;
        RECT 1190.550 472.840 1190.870 472.900 ;
        RECT 1186.870 472.700 1190.870 472.840 ;
        RECT 1186.870 472.640 1187.190 472.700 ;
        RECT 1190.550 472.640 1190.870 472.700 ;
        RECT 1090.730 18.600 1091.050 18.660 ;
        RECT 1186.870 18.600 1187.190 18.660 ;
        RECT 1090.730 18.460 1187.190 18.600 ;
        RECT 1090.730 18.400 1091.050 18.460 ;
        RECT 1186.870 18.400 1187.190 18.460 ;
      LAYER via ;
        RECT 1186.900 472.640 1187.160 472.900 ;
        RECT 1190.580 472.640 1190.840 472.900 ;
        RECT 1090.760 18.400 1091.020 18.660 ;
        RECT 1186.900 18.400 1187.160 18.660 ;
      LAYER met2 ;
        RECT 1192.550 510.410 1192.830 514.000 ;
        RECT 1190.640 510.270 1192.830 510.410 ;
        RECT 1190.640 472.930 1190.780 510.270 ;
        RECT 1192.550 510.000 1192.830 510.270 ;
        RECT 1186.900 472.610 1187.160 472.930 ;
        RECT 1190.580 472.610 1190.840 472.930 ;
        RECT 1186.960 18.690 1187.100 472.610 ;
        RECT 1090.760 18.370 1091.020 18.690 ;
        RECT 1186.900 18.370 1187.160 18.690 ;
        RECT 1090.820 2.400 1090.960 18.370 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.670 472.840 1200.990 472.900 ;
        RECT 1203.430 472.840 1203.750 472.900 ;
        RECT 1200.670 472.700 1203.750 472.840 ;
        RECT 1200.670 472.640 1200.990 472.700 ;
        RECT 1203.430 472.640 1203.750 472.700 ;
        RECT 1108.670 18.260 1108.990 18.320 ;
        RECT 1200.670 18.260 1200.990 18.320 ;
        RECT 1108.670 18.120 1200.990 18.260 ;
        RECT 1108.670 18.060 1108.990 18.120 ;
        RECT 1200.670 18.060 1200.990 18.120 ;
      LAYER via ;
        RECT 1200.700 472.640 1200.960 472.900 ;
        RECT 1203.460 472.640 1203.720 472.900 ;
        RECT 1108.700 18.060 1108.960 18.320 ;
        RECT 1200.700 18.060 1200.960 18.320 ;
      LAYER met2 ;
        RECT 1205.430 510.410 1205.710 514.000 ;
        RECT 1203.520 510.270 1205.710 510.410 ;
        RECT 1203.520 472.930 1203.660 510.270 ;
        RECT 1205.430 510.000 1205.710 510.270 ;
        RECT 1200.700 472.610 1200.960 472.930 ;
        RECT 1203.460 472.610 1203.720 472.930 ;
        RECT 1200.760 18.350 1200.900 472.610 ;
        RECT 1108.700 18.030 1108.960 18.350 ;
        RECT 1200.700 18.030 1200.960 18.350 ;
        RECT 1108.760 2.400 1108.900 18.030 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 19.620 1126.930 19.680 ;
        RECT 1214.470 19.620 1214.790 19.680 ;
        RECT 1126.610 19.480 1214.790 19.620 ;
        RECT 1126.610 19.420 1126.930 19.480 ;
        RECT 1214.470 19.420 1214.790 19.480 ;
      LAYER via ;
        RECT 1126.640 19.420 1126.900 19.680 ;
        RECT 1214.500 19.420 1214.760 19.680 ;
      LAYER met2 ;
        RECT 1218.310 511.090 1218.590 514.000 ;
        RECT 1215.020 510.950 1218.590 511.090 ;
        RECT 1215.020 449.210 1215.160 510.950 ;
        RECT 1218.310 510.000 1218.590 510.950 ;
        RECT 1214.560 449.070 1215.160 449.210 ;
        RECT 1214.560 19.710 1214.700 449.070 ;
        RECT 1126.640 19.390 1126.900 19.710 ;
        RECT 1214.500 19.390 1214.760 19.710 ;
        RECT 1126.700 2.400 1126.840 19.390 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.550 19.280 1144.870 19.340 ;
        RECT 1228.270 19.280 1228.590 19.340 ;
        RECT 1144.550 19.140 1228.590 19.280 ;
        RECT 1144.550 19.080 1144.870 19.140 ;
        RECT 1228.270 19.080 1228.590 19.140 ;
      LAYER via ;
        RECT 1144.580 19.080 1144.840 19.340 ;
        RECT 1228.300 19.080 1228.560 19.340 ;
      LAYER met2 ;
        RECT 1231.190 510.410 1231.470 514.000 ;
        RECT 1228.360 510.270 1231.470 510.410 ;
        RECT 1228.360 19.370 1228.500 510.270 ;
        RECT 1231.190 510.000 1231.470 510.270 ;
        RECT 1144.580 19.050 1144.840 19.370 ;
        RECT 1228.300 19.050 1228.560 19.370 ;
        RECT 1144.640 2.400 1144.780 19.050 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 17.920 1162.810 17.980 ;
        RECT 1242.070 17.920 1242.390 17.980 ;
        RECT 1162.490 17.780 1242.390 17.920 ;
        RECT 1162.490 17.720 1162.810 17.780 ;
        RECT 1242.070 17.720 1242.390 17.780 ;
      LAYER via ;
        RECT 1162.520 17.720 1162.780 17.980 ;
        RECT 1242.100 17.720 1242.360 17.980 ;
      LAYER met2 ;
        RECT 1244.070 510.410 1244.350 514.000 ;
        RECT 1242.160 510.270 1244.350 510.410 ;
        RECT 1242.160 18.010 1242.300 510.270 ;
        RECT 1244.070 510.000 1244.350 510.270 ;
        RECT 1162.520 17.690 1162.780 18.010 ;
        RECT 1242.100 17.690 1242.360 18.010 ;
        RECT 1162.580 2.400 1162.720 17.690 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 196.760 683.030 196.820 ;
        RECT 897.530 196.760 897.850 196.820 ;
        RECT 682.710 196.620 897.850 196.760 ;
        RECT 682.710 196.560 683.030 196.620 ;
        RECT 897.530 196.560 897.850 196.620 ;
        RECT 680.410 16.900 680.730 16.960 ;
        RECT 682.710 16.900 683.030 16.960 ;
        RECT 680.410 16.760 683.030 16.900 ;
        RECT 680.410 16.700 680.730 16.760 ;
        RECT 682.710 16.700 683.030 16.760 ;
      LAYER via ;
        RECT 682.740 196.560 683.000 196.820 ;
        RECT 897.560 196.560 897.820 196.820 ;
        RECT 680.440 16.700 680.700 16.960 ;
        RECT 682.740 16.700 683.000 16.960 ;
      LAYER met2 ;
        RECT 898.150 510.410 898.430 514.000 ;
        RECT 897.620 510.270 898.430 510.410 ;
        RECT 897.620 196.850 897.760 510.270 ;
        RECT 898.150 510.000 898.430 510.270 ;
        RECT 682.740 196.530 683.000 196.850 ;
        RECT 897.560 196.530 897.820 196.850 ;
        RECT 682.800 16.990 682.940 196.530 ;
        RECT 680.440 16.670 680.700 16.990 ;
        RECT 682.740 16.670 683.000 16.990 ;
        RECT 680.500 2.400 680.640 16.670 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 20.640 1180.290 20.700 ;
        RECT 1255.870 20.640 1256.190 20.700 ;
        RECT 1179.970 20.500 1256.190 20.640 ;
        RECT 1179.970 20.440 1180.290 20.500 ;
        RECT 1255.870 20.440 1256.190 20.500 ;
      LAYER via ;
        RECT 1180.000 20.440 1180.260 20.700 ;
        RECT 1255.900 20.440 1256.160 20.700 ;
      LAYER met2 ;
        RECT 1256.950 510.410 1257.230 514.000 ;
        RECT 1255.960 510.270 1257.230 510.410 ;
        RECT 1255.960 20.730 1256.100 510.270 ;
        RECT 1256.950 510.000 1257.230 510.270 ;
        RECT 1180.000 20.410 1180.260 20.730 ;
        RECT 1255.900 20.410 1256.160 20.730 ;
        RECT 1180.060 2.400 1180.200 20.410 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1263.305 386.325 1263.475 434.775 ;
        RECT 1262.385 234.685 1262.555 242.335 ;
      LAYER mcon ;
        RECT 1263.305 434.605 1263.475 434.775 ;
        RECT 1262.385 242.165 1262.555 242.335 ;
      LAYER met1 ;
        RECT 1263.245 434.760 1263.535 434.805 ;
        RECT 1263.690 434.760 1264.010 434.820 ;
        RECT 1263.245 434.620 1264.010 434.760 ;
        RECT 1263.245 434.575 1263.535 434.620 ;
        RECT 1263.690 434.560 1264.010 434.620 ;
        RECT 1263.230 386.480 1263.550 386.540 ;
        RECT 1263.035 386.340 1263.550 386.480 ;
        RECT 1263.230 386.280 1263.550 386.340 ;
        RECT 1262.310 357.920 1262.630 357.980 ;
        RECT 1263.230 357.920 1263.550 357.980 ;
        RECT 1262.310 357.780 1263.550 357.920 ;
        RECT 1262.310 357.720 1262.630 357.780 ;
        RECT 1263.230 357.720 1263.550 357.780 ;
        RECT 1262.310 289.920 1262.630 289.980 ;
        RECT 1263.230 289.920 1263.550 289.980 ;
        RECT 1262.310 289.780 1263.550 289.920 ;
        RECT 1262.310 289.720 1262.630 289.780 ;
        RECT 1263.230 289.720 1263.550 289.780 ;
        RECT 1262.325 242.320 1262.615 242.365 ;
        RECT 1263.230 242.320 1263.550 242.380 ;
        RECT 1262.325 242.180 1263.550 242.320 ;
        RECT 1262.325 242.135 1262.615 242.180 ;
        RECT 1263.230 242.120 1263.550 242.180 ;
        RECT 1262.310 234.840 1262.630 234.900 ;
        RECT 1262.115 234.700 1262.630 234.840 ;
        RECT 1262.310 234.640 1262.630 234.700 ;
        RECT 1262.310 193.360 1262.630 193.420 ;
        RECT 1263.230 193.360 1263.550 193.420 ;
        RECT 1262.310 193.220 1263.550 193.360 ;
        RECT 1262.310 193.160 1262.630 193.220 ;
        RECT 1263.230 193.160 1263.550 193.220 ;
        RECT 1197.910 18.600 1198.230 18.660 ;
        RECT 1263.230 18.600 1263.550 18.660 ;
        RECT 1197.910 18.460 1263.550 18.600 ;
        RECT 1197.910 18.400 1198.230 18.460 ;
        RECT 1263.230 18.400 1263.550 18.460 ;
      LAYER via ;
        RECT 1263.720 434.560 1263.980 434.820 ;
        RECT 1263.260 386.280 1263.520 386.540 ;
        RECT 1262.340 357.720 1262.600 357.980 ;
        RECT 1263.260 357.720 1263.520 357.980 ;
        RECT 1262.340 289.720 1262.600 289.980 ;
        RECT 1263.260 289.720 1263.520 289.980 ;
        RECT 1263.260 242.120 1263.520 242.380 ;
        RECT 1262.340 234.640 1262.600 234.900 ;
        RECT 1262.340 193.160 1262.600 193.420 ;
        RECT 1263.260 193.160 1263.520 193.420 ;
        RECT 1197.940 18.400 1198.200 18.660 ;
        RECT 1263.260 18.400 1263.520 18.660 ;
      LAYER met2 ;
        RECT 1269.370 511.090 1269.650 514.000 ;
        RECT 1266.080 510.950 1269.650 511.090 ;
        RECT 1266.080 449.210 1266.220 510.950 ;
        RECT 1269.370 510.000 1269.650 510.950 ;
        RECT 1265.160 449.070 1266.220 449.210 ;
        RECT 1265.160 448.530 1265.300 449.070 ;
        RECT 1263.780 448.390 1265.300 448.530 ;
        RECT 1263.780 434.850 1263.920 448.390 ;
        RECT 1263.720 434.530 1263.980 434.850 ;
        RECT 1263.260 386.250 1263.520 386.570 ;
        RECT 1263.320 358.010 1263.460 386.250 ;
        RECT 1262.340 357.690 1262.600 358.010 ;
        RECT 1263.260 357.690 1263.520 358.010 ;
        RECT 1262.400 290.010 1262.540 357.690 ;
        RECT 1262.340 289.690 1262.600 290.010 ;
        RECT 1263.260 289.690 1263.520 290.010 ;
        RECT 1263.320 242.410 1263.460 289.690 ;
        RECT 1263.260 242.090 1263.520 242.410 ;
        RECT 1262.340 234.610 1262.600 234.930 ;
        RECT 1262.400 193.450 1262.540 234.610 ;
        RECT 1262.340 193.130 1262.600 193.450 ;
        RECT 1263.260 193.130 1263.520 193.450 ;
        RECT 1263.320 18.690 1263.460 193.130 ;
        RECT 1197.940 18.370 1198.200 18.690 ;
        RECT 1263.260 18.370 1263.520 18.690 ;
        RECT 1198.000 2.400 1198.140 18.370 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1277.105 89.845 1277.275 137.955 ;
      LAYER mcon ;
        RECT 1277.105 137.785 1277.275 137.955 ;
      LAYER met1 ;
        RECT 1279.330 476.240 1279.650 476.300 ;
        RECT 1282.090 476.240 1282.410 476.300 ;
        RECT 1279.330 476.100 1282.410 476.240 ;
        RECT 1279.330 476.040 1279.650 476.100 ;
        RECT 1282.090 476.040 1282.410 476.100 ;
        RECT 1277.030 338.200 1277.350 338.260 ;
        RECT 1277.490 338.200 1277.810 338.260 ;
        RECT 1277.030 338.060 1277.810 338.200 ;
        RECT 1277.030 338.000 1277.350 338.060 ;
        RECT 1277.490 338.000 1277.810 338.060 ;
        RECT 1277.030 137.940 1277.350 138.000 ;
        RECT 1276.835 137.800 1277.350 137.940 ;
        RECT 1277.030 137.740 1277.350 137.800 ;
        RECT 1277.030 90.000 1277.350 90.060 ;
        RECT 1276.835 89.860 1277.350 90.000 ;
        RECT 1277.030 89.800 1277.350 89.860 ;
        RECT 1215.850 19.620 1216.170 19.680 ;
        RECT 1277.030 19.620 1277.350 19.680 ;
        RECT 1215.850 19.480 1277.350 19.620 ;
        RECT 1215.850 19.420 1216.170 19.480 ;
        RECT 1277.030 19.420 1277.350 19.480 ;
      LAYER via ;
        RECT 1279.360 476.040 1279.620 476.300 ;
        RECT 1282.120 476.040 1282.380 476.300 ;
        RECT 1277.060 338.000 1277.320 338.260 ;
        RECT 1277.520 338.000 1277.780 338.260 ;
        RECT 1277.060 137.740 1277.320 138.000 ;
        RECT 1277.060 89.800 1277.320 90.060 ;
        RECT 1215.880 19.420 1216.140 19.680 ;
        RECT 1277.060 19.420 1277.320 19.680 ;
      LAYER met2 ;
        RECT 1282.250 510.340 1282.530 514.000 ;
        RECT 1282.180 510.000 1282.530 510.340 ;
        RECT 1282.180 476.330 1282.320 510.000 ;
        RECT 1279.360 476.010 1279.620 476.330 ;
        RECT 1282.120 476.010 1282.380 476.330 ;
        RECT 1279.420 435.725 1279.560 476.010 ;
        RECT 1279.350 435.355 1279.630 435.725 ;
        RECT 1277.050 434.675 1277.330 435.045 ;
        RECT 1277.120 339.050 1277.260 434.675 ;
        RECT 1277.120 338.910 1277.720 339.050 ;
        RECT 1277.580 338.290 1277.720 338.910 ;
        RECT 1277.060 337.970 1277.320 338.290 ;
        RECT 1277.520 337.970 1277.780 338.290 ;
        RECT 1277.120 138.030 1277.260 337.970 ;
        RECT 1277.060 137.710 1277.320 138.030 ;
        RECT 1277.060 89.770 1277.320 90.090 ;
        RECT 1277.120 19.710 1277.260 89.770 ;
        RECT 1215.880 19.390 1216.140 19.710 ;
        RECT 1277.060 19.390 1277.320 19.710 ;
        RECT 1215.940 2.400 1216.080 19.390 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
      LAYER via2 ;
        RECT 1279.350 435.400 1279.630 435.680 ;
        RECT 1277.050 434.720 1277.330 435.000 ;
      LAYER met3 ;
        RECT 1279.325 435.690 1279.655 435.705 ;
        RECT 1276.350 435.390 1279.655 435.690 ;
        RECT 1276.350 435.010 1276.650 435.390 ;
        RECT 1279.325 435.375 1279.655 435.390 ;
        RECT 1277.025 435.010 1277.355 435.025 ;
        RECT 1276.350 434.710 1277.355 435.010 ;
        RECT 1277.025 434.695 1277.355 434.710 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1291.365 421.005 1291.535 469.115 ;
        RECT 1290.905 234.685 1291.075 282.455 ;
      LAYER mcon ;
        RECT 1291.365 468.945 1291.535 469.115 ;
        RECT 1290.905 282.285 1291.075 282.455 ;
      LAYER met1 ;
        RECT 1291.750 476.240 1292.070 476.300 ;
        RECT 1294.970 476.240 1295.290 476.300 ;
        RECT 1291.750 476.100 1295.290 476.240 ;
        RECT 1291.750 476.040 1292.070 476.100 ;
        RECT 1294.970 476.040 1295.290 476.100 ;
        RECT 1291.305 469.100 1291.595 469.145 ;
        RECT 1291.750 469.100 1292.070 469.160 ;
        RECT 1291.305 468.960 1292.070 469.100 ;
        RECT 1291.305 468.915 1291.595 468.960 ;
        RECT 1291.750 468.900 1292.070 468.960 ;
        RECT 1291.290 421.160 1291.610 421.220 ;
        RECT 1291.095 421.020 1291.610 421.160 ;
        RECT 1291.290 420.960 1291.610 421.020 ;
        RECT 1291.290 386.620 1291.610 386.880 ;
        RECT 1291.380 386.200 1291.520 386.620 ;
        RECT 1291.290 385.940 1291.610 386.200 ;
        RECT 1290.830 331.400 1291.150 331.460 ;
        RECT 1291.290 331.400 1291.610 331.460 ;
        RECT 1290.830 331.260 1291.610 331.400 ;
        RECT 1290.830 331.200 1291.150 331.260 ;
        RECT 1291.290 331.200 1291.610 331.260 ;
        RECT 1290.830 282.440 1291.150 282.500 ;
        RECT 1290.635 282.300 1291.150 282.440 ;
        RECT 1290.830 282.240 1291.150 282.300 ;
        RECT 1290.830 234.840 1291.150 234.900 ;
        RECT 1290.635 234.700 1291.150 234.840 ;
        RECT 1290.830 234.640 1291.150 234.700 ;
        RECT 1290.830 193.020 1291.150 193.080 ;
        RECT 1291.290 193.020 1291.610 193.080 ;
        RECT 1290.830 192.880 1291.610 193.020 ;
        RECT 1290.830 192.820 1291.150 192.880 ;
        RECT 1291.290 192.820 1291.610 192.880 ;
        RECT 1233.790 19.280 1234.110 19.340 ;
        RECT 1291.750 19.280 1292.070 19.340 ;
        RECT 1233.790 19.140 1292.070 19.280 ;
        RECT 1233.790 19.080 1234.110 19.140 ;
        RECT 1291.750 19.080 1292.070 19.140 ;
      LAYER via ;
        RECT 1291.780 476.040 1292.040 476.300 ;
        RECT 1295.000 476.040 1295.260 476.300 ;
        RECT 1291.780 468.900 1292.040 469.160 ;
        RECT 1291.320 420.960 1291.580 421.220 ;
        RECT 1291.320 386.620 1291.580 386.880 ;
        RECT 1291.320 385.940 1291.580 386.200 ;
        RECT 1290.860 331.200 1291.120 331.460 ;
        RECT 1291.320 331.200 1291.580 331.460 ;
        RECT 1290.860 282.240 1291.120 282.500 ;
        RECT 1290.860 234.640 1291.120 234.900 ;
        RECT 1290.860 192.820 1291.120 193.080 ;
        RECT 1291.320 192.820 1291.580 193.080 ;
        RECT 1233.820 19.080 1234.080 19.340 ;
        RECT 1291.780 19.080 1292.040 19.340 ;
      LAYER met2 ;
        RECT 1295.130 510.340 1295.410 514.000 ;
        RECT 1295.060 510.000 1295.410 510.340 ;
        RECT 1295.060 476.330 1295.200 510.000 ;
        RECT 1291.780 476.010 1292.040 476.330 ;
        RECT 1295.000 476.010 1295.260 476.330 ;
        RECT 1291.840 469.190 1291.980 476.010 ;
        RECT 1291.780 468.870 1292.040 469.190 ;
        RECT 1291.320 420.930 1291.580 421.250 ;
        RECT 1291.380 386.910 1291.520 420.930 ;
        RECT 1291.320 386.590 1291.580 386.910 ;
        RECT 1291.320 385.910 1291.580 386.230 ;
        RECT 1291.380 331.490 1291.520 385.910 ;
        RECT 1290.860 331.170 1291.120 331.490 ;
        RECT 1291.320 331.170 1291.580 331.490 ;
        RECT 1290.920 282.530 1291.060 331.170 ;
        RECT 1290.860 282.210 1291.120 282.530 ;
        RECT 1290.860 234.610 1291.120 234.930 ;
        RECT 1290.920 193.110 1291.060 234.610 ;
        RECT 1290.860 192.790 1291.120 193.110 ;
        RECT 1291.320 192.790 1291.580 193.110 ;
        RECT 1291.380 62.290 1291.520 192.790 ;
        RECT 1291.380 62.150 1291.980 62.290 ;
        RECT 1291.840 19.370 1291.980 62.150 ;
        RECT 1233.820 19.050 1234.080 19.370 ;
        RECT 1291.780 19.050 1292.040 19.370 ;
        RECT 1233.880 2.400 1234.020 19.050 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1304.245 241.485 1304.415 289.595 ;
        RECT 1304.245 193.545 1304.415 240.975 ;
        RECT 1304.245 48.365 1304.415 96.475 ;
      LAYER mcon ;
        RECT 1304.245 289.425 1304.415 289.595 ;
        RECT 1304.245 240.805 1304.415 240.975 ;
        RECT 1304.245 96.305 1304.415 96.475 ;
      LAYER met1 ;
        RECT 1304.170 289.580 1304.490 289.640 ;
        RECT 1304.170 289.440 1304.685 289.580 ;
        RECT 1304.170 289.380 1304.490 289.440 ;
        RECT 1304.170 241.640 1304.490 241.700 ;
        RECT 1304.170 241.500 1304.685 241.640 ;
        RECT 1304.170 241.440 1304.490 241.500 ;
        RECT 1304.170 240.960 1304.490 241.020 ;
        RECT 1304.170 240.820 1304.685 240.960 ;
        RECT 1304.170 240.760 1304.490 240.820 ;
        RECT 1304.170 193.700 1304.490 193.760 ;
        RECT 1304.170 193.560 1304.685 193.700 ;
        RECT 1304.170 193.500 1304.490 193.560 ;
        RECT 1304.170 96.460 1304.490 96.520 ;
        RECT 1304.170 96.320 1304.685 96.460 ;
        RECT 1304.170 96.260 1304.490 96.320 ;
        RECT 1304.185 48.520 1304.475 48.565 ;
        RECT 1305.090 48.520 1305.410 48.580 ;
        RECT 1304.185 48.380 1305.410 48.520 ;
        RECT 1304.185 48.335 1304.475 48.380 ;
        RECT 1305.090 48.320 1305.410 48.380 ;
        RECT 1251.730 16.900 1252.050 16.960 ;
        RECT 1305.090 16.900 1305.410 16.960 ;
        RECT 1251.730 16.760 1305.410 16.900 ;
        RECT 1251.730 16.700 1252.050 16.760 ;
        RECT 1305.090 16.700 1305.410 16.760 ;
      LAYER via ;
        RECT 1304.200 289.380 1304.460 289.640 ;
        RECT 1304.200 241.440 1304.460 241.700 ;
        RECT 1304.200 240.760 1304.460 241.020 ;
        RECT 1304.200 193.500 1304.460 193.760 ;
        RECT 1304.200 96.260 1304.460 96.520 ;
        RECT 1305.120 48.320 1305.380 48.580 ;
        RECT 1251.760 16.700 1252.020 16.960 ;
        RECT 1305.120 16.700 1305.380 16.960 ;
      LAYER met2 ;
        RECT 1308.010 510.410 1308.290 514.000 ;
        RECT 1306.100 510.270 1308.290 510.410 ;
        RECT 1306.100 386.765 1306.240 510.270 ;
        RECT 1308.010 510.000 1308.290 510.270 ;
        RECT 1306.030 386.395 1306.310 386.765 ;
        RECT 1304.190 385.715 1304.470 386.085 ;
        RECT 1304.260 289.670 1304.400 385.715 ;
        RECT 1304.200 289.350 1304.460 289.670 ;
        RECT 1304.200 241.410 1304.460 241.730 ;
        RECT 1304.260 241.050 1304.400 241.410 ;
        RECT 1304.200 240.730 1304.460 241.050 ;
        RECT 1304.200 193.470 1304.460 193.790 ;
        RECT 1304.260 96.550 1304.400 193.470 ;
        RECT 1304.200 96.230 1304.460 96.550 ;
        RECT 1305.120 48.290 1305.380 48.610 ;
        RECT 1305.180 16.990 1305.320 48.290 ;
        RECT 1251.760 16.670 1252.020 16.990 ;
        RECT 1305.120 16.670 1305.380 16.990 ;
        RECT 1251.820 2.400 1251.960 16.670 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
      LAYER via2 ;
        RECT 1306.030 386.440 1306.310 386.720 ;
        RECT 1304.190 385.760 1304.470 386.040 ;
      LAYER met3 ;
        RECT 1306.005 386.730 1306.335 386.745 ;
        RECT 1304.870 386.430 1306.335 386.730 ;
        RECT 1304.165 386.050 1304.495 386.065 ;
        RECT 1304.870 386.050 1305.170 386.430 ;
        RECT 1306.005 386.415 1306.335 386.430 ;
        RECT 1304.165 385.750 1305.170 386.050 ;
        RECT 1304.165 385.735 1304.495 385.750 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 17.580 1269.530 17.640 ;
        RECT 1317.970 17.580 1318.290 17.640 ;
        RECT 1269.210 17.440 1318.290 17.580 ;
        RECT 1269.210 17.380 1269.530 17.440 ;
        RECT 1317.970 17.380 1318.290 17.440 ;
      LAYER via ;
        RECT 1269.240 17.380 1269.500 17.640 ;
        RECT 1318.000 17.380 1318.260 17.640 ;
      LAYER met2 ;
        RECT 1320.890 510.410 1321.170 514.000 ;
        RECT 1318.060 510.270 1321.170 510.410 ;
        RECT 1318.060 17.670 1318.200 510.270 ;
        RECT 1320.890 510.000 1321.170 510.270 ;
        RECT 1269.240 17.350 1269.500 17.670 ;
        RECT 1318.000 17.350 1318.260 17.670 ;
        RECT 1269.300 2.400 1269.440 17.350 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 18.600 1287.470 18.660 ;
        RECT 1331.770 18.600 1332.090 18.660 ;
        RECT 1287.150 18.460 1332.090 18.600 ;
        RECT 1287.150 18.400 1287.470 18.460 ;
        RECT 1331.770 18.400 1332.090 18.460 ;
      LAYER via ;
        RECT 1287.180 18.400 1287.440 18.660 ;
        RECT 1331.800 18.400 1332.060 18.660 ;
      LAYER met2 ;
        RECT 1333.770 510.410 1334.050 514.000 ;
        RECT 1331.860 510.270 1334.050 510.410 ;
        RECT 1331.860 18.690 1332.000 510.270 ;
        RECT 1333.770 510.000 1334.050 510.270 ;
        RECT 1287.180 18.370 1287.440 18.690 ;
        RECT 1331.800 18.370 1332.060 18.690 ;
        RECT 1287.240 2.400 1287.380 18.370 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1305.090 15.200 1305.410 15.260 ;
        RECT 1345.570 15.200 1345.890 15.260 ;
        RECT 1305.090 15.060 1345.890 15.200 ;
        RECT 1305.090 15.000 1305.410 15.060 ;
        RECT 1345.570 15.000 1345.890 15.060 ;
      LAYER via ;
        RECT 1305.120 15.000 1305.380 15.260 ;
        RECT 1345.600 15.000 1345.860 15.260 ;
      LAYER met2 ;
        RECT 1346.190 510.410 1346.470 514.000 ;
        RECT 1345.660 510.270 1346.470 510.410 ;
        RECT 1345.660 15.290 1345.800 510.270 ;
        RECT 1346.190 510.000 1346.470 510.270 ;
        RECT 1305.120 14.970 1305.380 15.290 ;
        RECT 1345.600 14.970 1345.860 15.290 ;
        RECT 1305.180 2.400 1305.320 14.970 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.470 457.880 1352.790 457.940 ;
        RECT 1357.070 457.880 1357.390 457.940 ;
        RECT 1352.470 457.740 1357.390 457.880 ;
        RECT 1352.470 457.680 1352.790 457.740 ;
        RECT 1357.070 457.680 1357.390 457.740 ;
        RECT 1323.030 17.920 1323.350 17.980 ;
        RECT 1352.470 17.920 1352.790 17.980 ;
        RECT 1323.030 17.780 1352.790 17.920 ;
        RECT 1323.030 17.720 1323.350 17.780 ;
        RECT 1352.470 17.720 1352.790 17.780 ;
      LAYER via ;
        RECT 1352.500 457.680 1352.760 457.940 ;
        RECT 1357.100 457.680 1357.360 457.940 ;
        RECT 1323.060 17.720 1323.320 17.980 ;
        RECT 1352.500 17.720 1352.760 17.980 ;
      LAYER met2 ;
        RECT 1359.070 510.410 1359.350 514.000 ;
        RECT 1357.160 510.270 1359.350 510.410 ;
        RECT 1357.160 457.970 1357.300 510.270 ;
        RECT 1359.070 510.000 1359.350 510.270 ;
        RECT 1352.500 457.650 1352.760 457.970 ;
        RECT 1357.100 457.650 1357.360 457.970 ;
        RECT 1352.560 18.010 1352.700 457.650 ;
        RECT 1323.060 17.690 1323.320 18.010 ;
        RECT 1352.500 17.690 1352.760 18.010 ;
        RECT 1323.120 2.400 1323.260 17.690 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.270 461.960 1366.590 462.020 ;
        RECT 1369.950 461.960 1370.270 462.020 ;
        RECT 1366.270 461.820 1370.270 461.960 ;
        RECT 1366.270 461.760 1366.590 461.820 ;
        RECT 1369.950 461.760 1370.270 461.820 ;
        RECT 1340.510 18.260 1340.830 18.320 ;
        RECT 1366.270 18.260 1366.590 18.320 ;
        RECT 1340.510 18.120 1366.590 18.260 ;
        RECT 1340.510 18.060 1340.830 18.120 ;
        RECT 1366.270 18.060 1366.590 18.120 ;
      LAYER via ;
        RECT 1366.300 461.760 1366.560 462.020 ;
        RECT 1369.980 461.760 1370.240 462.020 ;
        RECT 1340.540 18.060 1340.800 18.320 ;
        RECT 1366.300 18.060 1366.560 18.320 ;
      LAYER met2 ;
        RECT 1371.950 510.410 1372.230 514.000 ;
        RECT 1370.040 510.270 1372.230 510.410 ;
        RECT 1370.040 462.050 1370.180 510.270 ;
        RECT 1371.950 510.000 1372.230 510.270 ;
        RECT 1366.300 461.730 1366.560 462.050 ;
        RECT 1369.980 461.730 1370.240 462.050 ;
        RECT 1366.360 18.350 1366.500 461.730 ;
        RECT 1340.540 18.030 1340.800 18.350 ;
        RECT 1366.300 18.030 1366.560 18.350 ;
        RECT 1340.600 2.400 1340.740 18.030 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 203.560 703.730 203.620 ;
        RECT 911.330 203.560 911.650 203.620 ;
        RECT 703.410 203.420 911.650 203.560 ;
        RECT 703.410 203.360 703.730 203.420 ;
        RECT 911.330 203.360 911.650 203.420 ;
        RECT 698.350 16.900 698.670 16.960 ;
        RECT 703.410 16.900 703.730 16.960 ;
        RECT 698.350 16.760 703.730 16.900 ;
        RECT 698.350 16.700 698.670 16.760 ;
        RECT 703.410 16.700 703.730 16.760 ;
      LAYER via ;
        RECT 703.440 203.360 703.700 203.620 ;
        RECT 911.360 203.360 911.620 203.620 ;
        RECT 698.380 16.700 698.640 16.960 ;
        RECT 703.440 16.700 703.700 16.960 ;
      LAYER met2 ;
        RECT 911.030 510.340 911.310 514.000 ;
        RECT 910.960 510.000 911.310 510.340 ;
        RECT 910.960 473.690 911.100 510.000 ;
        RECT 910.960 473.550 911.560 473.690 ;
        RECT 911.420 203.650 911.560 473.550 ;
        RECT 703.440 203.330 703.700 203.650 ;
        RECT 911.360 203.330 911.620 203.650 ;
        RECT 703.500 16.990 703.640 203.330 ;
        RECT 698.380 16.670 698.640 16.990 ;
        RECT 703.440 16.670 703.700 16.990 ;
        RECT 698.440 2.400 698.580 16.670 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.070 472.840 1380.390 472.900 ;
        RECT 1382.830 472.840 1383.150 472.900 ;
        RECT 1380.070 472.700 1383.150 472.840 ;
        RECT 1380.070 472.640 1380.390 472.700 ;
        RECT 1382.830 472.640 1383.150 472.700 ;
        RECT 1358.450 20.640 1358.770 20.700 ;
        RECT 1380.070 20.640 1380.390 20.700 ;
        RECT 1358.450 20.500 1380.390 20.640 ;
        RECT 1358.450 20.440 1358.770 20.500 ;
        RECT 1380.070 20.440 1380.390 20.500 ;
      LAYER via ;
        RECT 1380.100 472.640 1380.360 472.900 ;
        RECT 1382.860 472.640 1383.120 472.900 ;
        RECT 1358.480 20.440 1358.740 20.700 ;
        RECT 1380.100 20.440 1380.360 20.700 ;
      LAYER met2 ;
        RECT 1384.830 510.410 1385.110 514.000 ;
        RECT 1382.920 510.270 1385.110 510.410 ;
        RECT 1382.920 472.930 1383.060 510.270 ;
        RECT 1384.830 510.000 1385.110 510.270 ;
        RECT 1380.100 472.610 1380.360 472.930 ;
        RECT 1382.860 472.610 1383.120 472.930 ;
        RECT 1380.160 20.730 1380.300 472.610 ;
        RECT 1358.480 20.410 1358.740 20.730 ;
        RECT 1380.100 20.410 1380.360 20.730 ;
        RECT 1358.540 2.400 1358.680 20.410 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.330 386.480 1394.650 386.540 ;
        RECT 1394.790 386.480 1395.110 386.540 ;
        RECT 1394.330 386.340 1395.110 386.480 ;
        RECT 1394.330 386.280 1394.650 386.340 ;
        RECT 1394.790 386.280 1395.110 386.340 ;
        RECT 1376.390 20.300 1376.710 20.360 ;
        RECT 1393.410 20.300 1393.730 20.360 ;
        RECT 1376.390 20.160 1393.730 20.300 ;
        RECT 1376.390 20.100 1376.710 20.160 ;
        RECT 1393.410 20.100 1393.730 20.160 ;
      LAYER via ;
        RECT 1394.360 386.280 1394.620 386.540 ;
        RECT 1394.820 386.280 1395.080 386.540 ;
        RECT 1376.420 20.100 1376.680 20.360 ;
        RECT 1393.440 20.100 1393.700 20.360 ;
      LAYER met2 ;
        RECT 1397.710 510.410 1397.990 514.000 ;
        RECT 1395.800 510.270 1397.990 510.410 ;
        RECT 1395.800 449.210 1395.940 510.270 ;
        RECT 1397.710 510.000 1397.990 510.270 ;
        RECT 1394.880 449.070 1395.940 449.210 ;
        RECT 1394.880 386.570 1395.020 449.070 ;
        RECT 1394.360 386.250 1394.620 386.570 ;
        RECT 1394.820 386.250 1395.080 386.570 ;
        RECT 1394.420 207.130 1394.560 386.250 ;
        RECT 1393.960 206.990 1394.560 207.130 ;
        RECT 1393.960 206.450 1394.100 206.990 ;
        RECT 1393.960 206.310 1394.560 206.450 ;
        RECT 1394.420 110.570 1394.560 206.310 ;
        RECT 1393.960 110.430 1394.560 110.570 ;
        RECT 1393.960 109.890 1394.100 110.430 ;
        RECT 1393.960 109.750 1394.560 109.890 ;
        RECT 1394.420 20.810 1394.560 109.750 ;
        RECT 1393.500 20.670 1394.560 20.810 ;
        RECT 1393.500 20.390 1393.640 20.670 ;
        RECT 1376.420 20.070 1376.680 20.390 ;
        RECT 1393.440 20.070 1393.700 20.390 ;
        RECT 1376.480 2.400 1376.620 20.070 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.330 20.300 1394.650 20.360 ;
        RECT 1407.670 20.300 1407.990 20.360 ;
        RECT 1394.330 20.160 1407.990 20.300 ;
        RECT 1394.330 20.100 1394.650 20.160 ;
        RECT 1407.670 20.100 1407.990 20.160 ;
      LAYER via ;
        RECT 1394.360 20.100 1394.620 20.360 ;
        RECT 1407.700 20.100 1407.960 20.360 ;
      LAYER met2 ;
        RECT 1410.590 510.410 1410.870 514.000 ;
        RECT 1407.760 510.270 1410.870 510.410 ;
        RECT 1407.760 20.390 1407.900 510.270 ;
        RECT 1410.590 510.000 1410.870 510.270 ;
        RECT 1394.360 20.070 1394.620 20.390 ;
        RECT 1407.700 20.070 1407.960 20.390 ;
        RECT 1394.420 2.400 1394.560 20.070 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1412.270 20.300 1412.590 20.360 ;
        RECT 1421.470 20.300 1421.790 20.360 ;
        RECT 1412.270 20.160 1421.790 20.300 ;
        RECT 1412.270 20.100 1412.590 20.160 ;
        RECT 1421.470 20.100 1421.790 20.160 ;
      LAYER via ;
        RECT 1412.300 20.100 1412.560 20.360 ;
        RECT 1421.500 20.100 1421.760 20.360 ;
      LAYER met2 ;
        RECT 1423.010 510.410 1423.290 514.000 ;
        RECT 1421.560 510.270 1423.290 510.410 ;
        RECT 1421.560 20.390 1421.700 510.270 ;
        RECT 1423.010 510.000 1423.290 510.270 ;
        RECT 1412.300 20.070 1412.560 20.390 ;
        RECT 1421.500 20.070 1421.760 20.390 ;
        RECT 1412.360 2.400 1412.500 20.070 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.750 17.920 1430.070 17.980 ;
        RECT 1435.270 17.920 1435.590 17.980 ;
        RECT 1429.750 17.780 1435.590 17.920 ;
        RECT 1429.750 17.720 1430.070 17.780 ;
        RECT 1435.270 17.720 1435.590 17.780 ;
      LAYER via ;
        RECT 1429.780 17.720 1430.040 17.980 ;
        RECT 1435.300 17.720 1435.560 17.980 ;
      LAYER met2 ;
        RECT 1435.890 510.410 1436.170 514.000 ;
        RECT 1435.360 510.270 1436.170 510.410 ;
        RECT 1435.360 18.010 1435.500 510.270 ;
        RECT 1435.890 510.000 1436.170 510.270 ;
        RECT 1429.780 17.690 1430.040 18.010 ;
        RECT 1435.300 17.690 1435.560 18.010 ;
        RECT 1429.840 2.400 1429.980 17.690 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.630 20.640 1442.950 20.700 ;
        RECT 1447.690 20.640 1448.010 20.700 ;
        RECT 1442.630 20.500 1448.010 20.640 ;
        RECT 1442.630 20.440 1442.950 20.500 ;
        RECT 1447.690 20.440 1448.010 20.500 ;
      LAYER via ;
        RECT 1442.660 20.440 1442.920 20.700 ;
        RECT 1447.720 20.440 1447.980 20.700 ;
      LAYER met2 ;
        RECT 1448.770 511.090 1449.050 514.000 ;
        RECT 1445.480 510.950 1449.050 511.090 ;
        RECT 1445.480 449.210 1445.620 510.950 ;
        RECT 1448.770 510.000 1449.050 510.950 ;
        RECT 1443.180 449.070 1445.620 449.210 ;
        RECT 1443.180 400.930 1443.320 449.070 ;
        RECT 1442.720 400.790 1443.320 400.930 ;
        RECT 1442.720 20.730 1442.860 400.790 ;
        RECT 1442.660 20.410 1442.920 20.730 ;
        RECT 1447.720 20.410 1447.980 20.730 ;
        RECT 1447.780 2.400 1447.920 20.410 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 17.240 1462.730 17.300 ;
        RECT 1465.630 17.240 1465.950 17.300 ;
        RECT 1462.410 17.100 1465.950 17.240 ;
        RECT 1462.410 17.040 1462.730 17.100 ;
        RECT 1465.630 17.040 1465.950 17.100 ;
      LAYER via ;
        RECT 1462.440 17.040 1462.700 17.300 ;
        RECT 1465.660 17.040 1465.920 17.300 ;
      LAYER met2 ;
        RECT 1461.650 510.410 1461.930 514.000 ;
        RECT 1461.650 510.270 1462.640 510.410 ;
        RECT 1461.650 510.000 1461.930 510.270 ;
        RECT 1462.500 17.330 1462.640 510.270 ;
        RECT 1462.440 17.010 1462.700 17.330 ;
        RECT 1465.660 17.010 1465.920 17.330 ;
        RECT 1465.720 2.400 1465.860 17.010 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1476.210 20.640 1476.530 20.700 ;
        RECT 1483.570 20.640 1483.890 20.700 ;
        RECT 1476.210 20.500 1483.890 20.640 ;
        RECT 1476.210 20.440 1476.530 20.500 ;
        RECT 1483.570 20.440 1483.890 20.500 ;
      LAYER via ;
        RECT 1476.240 20.440 1476.500 20.700 ;
        RECT 1483.600 20.440 1483.860 20.700 ;
      LAYER met2 ;
        RECT 1474.530 510.410 1474.810 514.000 ;
        RECT 1474.530 510.270 1476.440 510.410 ;
        RECT 1474.530 510.000 1474.810 510.270 ;
        RECT 1476.300 20.730 1476.440 510.270 ;
        RECT 1476.240 20.410 1476.500 20.730 ;
        RECT 1483.600 20.410 1483.860 20.730 ;
        RECT 1483.660 2.400 1483.800 20.410 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 15.540 1490.330 15.600 ;
        RECT 1501.510 15.540 1501.830 15.600 ;
        RECT 1490.010 15.400 1501.830 15.540 ;
        RECT 1490.010 15.340 1490.330 15.400 ;
        RECT 1501.510 15.340 1501.830 15.400 ;
      LAYER via ;
        RECT 1490.040 15.340 1490.300 15.600 ;
        RECT 1501.540 15.340 1501.800 15.600 ;
      LAYER met2 ;
        RECT 1487.410 510.410 1487.690 514.000 ;
        RECT 1487.410 510.270 1490.240 510.410 ;
        RECT 1487.410 510.000 1487.690 510.270 ;
        RECT 1490.100 15.630 1490.240 510.270 ;
        RECT 1490.040 15.310 1490.300 15.630 ;
        RECT 1501.540 15.310 1501.800 15.630 ;
        RECT 1501.600 2.400 1501.740 15.310 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1503.810 17.580 1504.130 17.640 ;
        RECT 1518.990 17.580 1519.310 17.640 ;
        RECT 1503.810 17.440 1519.310 17.580 ;
        RECT 1503.810 17.380 1504.130 17.440 ;
        RECT 1518.990 17.380 1519.310 17.440 ;
      LAYER via ;
        RECT 1503.840 17.380 1504.100 17.640 ;
        RECT 1519.020 17.380 1519.280 17.640 ;
      LAYER met2 ;
        RECT 1500.290 510.410 1500.570 514.000 ;
        RECT 1500.290 510.270 1504.040 510.410 ;
        RECT 1500.290 510.000 1500.570 510.270 ;
        RECT 1503.900 17.670 1504.040 510.270 ;
        RECT 1503.840 17.350 1504.100 17.670 ;
        RECT 1519.020 17.350 1519.280 17.670 ;
        RECT 1519.080 2.400 1519.220 17.350 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 920.145 399.925 920.315 434.775 ;
        RECT 918.765 331.245 918.935 386.155 ;
      LAYER mcon ;
        RECT 920.145 434.605 920.315 434.775 ;
        RECT 918.765 385.985 918.935 386.155 ;
      LAYER met1 ;
        RECT 920.070 434.760 920.390 434.820 ;
        RECT 919.875 434.620 920.390 434.760 ;
        RECT 920.070 434.560 920.390 434.620 ;
        RECT 918.690 400.080 919.010 400.140 ;
        RECT 920.085 400.080 920.375 400.125 ;
        RECT 918.690 399.940 920.375 400.080 ;
        RECT 918.690 399.880 919.010 399.940 ;
        RECT 920.085 399.895 920.375 399.940 ;
        RECT 918.690 386.140 919.010 386.200 ;
        RECT 918.495 386.000 919.010 386.140 ;
        RECT 918.690 385.940 919.010 386.000 ;
        RECT 918.690 331.400 919.010 331.460 ;
        RECT 918.495 331.260 919.010 331.400 ;
        RECT 918.690 331.200 919.010 331.260 ;
        RECT 918.690 289.720 919.010 289.980 ;
        RECT 918.780 289.300 918.920 289.720 ;
        RECT 918.690 289.040 919.010 289.300 ;
        RECT 918.690 255.380 919.010 255.640 ;
        RECT 918.780 254.960 918.920 255.380 ;
        RECT 918.690 254.700 919.010 254.960 ;
        RECT 717.210 210.360 717.530 210.420 ;
        RECT 918.690 210.360 919.010 210.420 ;
        RECT 717.210 210.220 919.010 210.360 ;
        RECT 717.210 210.160 717.530 210.220 ;
        RECT 918.690 210.160 919.010 210.220 ;
      LAYER via ;
        RECT 920.100 434.560 920.360 434.820 ;
        RECT 918.720 399.880 918.980 400.140 ;
        RECT 918.720 385.940 918.980 386.200 ;
        RECT 918.720 331.200 918.980 331.460 ;
        RECT 918.720 289.720 918.980 289.980 ;
        RECT 918.720 289.040 918.980 289.300 ;
        RECT 918.720 255.380 918.980 255.640 ;
        RECT 918.720 254.700 918.980 254.960 ;
        RECT 717.240 210.160 717.500 210.420 ;
        RECT 918.720 210.160 918.980 210.420 ;
      LAYER met2 ;
        RECT 923.910 511.090 924.190 514.000 ;
        RECT 920.620 510.950 924.190 511.090 ;
        RECT 920.620 449.210 920.760 510.950 ;
        RECT 923.910 510.000 924.190 510.950 ;
        RECT 920.160 449.070 920.760 449.210 ;
        RECT 920.160 434.850 920.300 449.070 ;
        RECT 920.100 434.530 920.360 434.850 ;
        RECT 918.720 399.850 918.980 400.170 ;
        RECT 918.780 386.230 918.920 399.850 ;
        RECT 918.720 385.910 918.980 386.230 ;
        RECT 918.720 331.170 918.980 331.490 ;
        RECT 918.780 290.010 918.920 331.170 ;
        RECT 918.720 289.690 918.980 290.010 ;
        RECT 918.720 289.010 918.980 289.330 ;
        RECT 918.780 255.670 918.920 289.010 ;
        RECT 918.720 255.350 918.980 255.670 ;
        RECT 918.720 254.670 918.980 254.990 ;
        RECT 918.780 210.450 918.920 254.670 ;
        RECT 717.240 210.130 717.500 210.450 ;
        RECT 918.720 210.130 918.980 210.450 ;
        RECT 717.300 16.900 717.440 210.130 ;
        RECT 716.380 16.760 717.440 16.900 ;
        RECT 716.380 2.400 716.520 16.760 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1512.550 503.440 1512.870 503.500 ;
        RECT 1517.610 503.440 1517.930 503.500 ;
        RECT 1512.550 503.300 1517.930 503.440 ;
        RECT 1512.550 503.240 1512.870 503.300 ;
        RECT 1517.610 503.240 1517.930 503.300 ;
        RECT 1517.610 20.640 1517.930 20.700 ;
        RECT 1536.930 20.640 1537.250 20.700 ;
        RECT 1517.610 20.500 1537.250 20.640 ;
        RECT 1517.610 20.440 1517.930 20.500 ;
        RECT 1536.930 20.440 1537.250 20.500 ;
      LAYER via ;
        RECT 1512.580 503.240 1512.840 503.500 ;
        RECT 1517.640 503.240 1517.900 503.500 ;
        RECT 1517.640 20.440 1517.900 20.700 ;
        RECT 1536.960 20.440 1537.220 20.700 ;
      LAYER met2 ;
        RECT 1512.710 510.340 1512.990 514.000 ;
        RECT 1512.640 510.000 1512.990 510.340 ;
        RECT 1512.640 503.530 1512.780 510.000 ;
        RECT 1512.580 503.210 1512.840 503.530 ;
        RECT 1517.640 503.210 1517.900 503.530 ;
        RECT 1517.700 20.730 1517.840 503.210 ;
        RECT 1517.640 20.410 1517.900 20.730 ;
        RECT 1536.960 20.410 1537.220 20.730 ;
        RECT 1537.020 2.400 1537.160 20.410 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1525.430 503.100 1525.750 503.160 ;
        RECT 1531.410 503.100 1531.730 503.160 ;
        RECT 1525.430 502.960 1531.730 503.100 ;
        RECT 1525.430 502.900 1525.750 502.960 ;
        RECT 1531.410 502.900 1531.730 502.960 ;
        RECT 1531.410 20.300 1531.730 20.360 ;
        RECT 1554.870 20.300 1555.190 20.360 ;
        RECT 1531.410 20.160 1555.190 20.300 ;
        RECT 1531.410 20.100 1531.730 20.160 ;
        RECT 1554.870 20.100 1555.190 20.160 ;
      LAYER via ;
        RECT 1525.460 502.900 1525.720 503.160 ;
        RECT 1531.440 502.900 1531.700 503.160 ;
        RECT 1531.440 20.100 1531.700 20.360 ;
        RECT 1554.900 20.100 1555.160 20.360 ;
      LAYER met2 ;
        RECT 1525.590 510.340 1525.870 514.000 ;
        RECT 1525.520 510.000 1525.870 510.340 ;
        RECT 1525.520 503.190 1525.660 510.000 ;
        RECT 1525.460 502.870 1525.720 503.190 ;
        RECT 1531.440 502.870 1531.700 503.190 ;
        RECT 1531.500 20.390 1531.640 502.870 ;
        RECT 1531.440 20.070 1531.700 20.390 ;
        RECT 1554.900 20.070 1555.160 20.390 ;
        RECT 1554.960 2.400 1555.100 20.070 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 16.560 1538.630 16.620 ;
        RECT 1572.810 16.560 1573.130 16.620 ;
        RECT 1538.310 16.420 1573.130 16.560 ;
        RECT 1538.310 16.360 1538.630 16.420 ;
        RECT 1572.810 16.360 1573.130 16.420 ;
      LAYER via ;
        RECT 1538.340 16.360 1538.600 16.620 ;
        RECT 1572.840 16.360 1573.100 16.620 ;
      LAYER met2 ;
        RECT 1538.470 510.340 1538.750 514.000 ;
        RECT 1538.400 510.000 1538.750 510.340 ;
        RECT 1538.400 16.650 1538.540 510.000 ;
        RECT 1538.340 16.330 1538.600 16.650 ;
        RECT 1572.840 16.330 1573.100 16.650 ;
        RECT 1572.900 2.400 1573.040 16.330 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1550.805 399.925 1550.975 434.775 ;
        RECT 1551.265 295.885 1551.435 317.475 ;
        RECT 1551.265 203.405 1551.435 227.715 ;
        RECT 1551.265 61.625 1551.435 137.615 ;
      LAYER mcon ;
        RECT 1550.805 434.605 1550.975 434.775 ;
        RECT 1551.265 317.305 1551.435 317.475 ;
        RECT 1551.265 227.545 1551.435 227.715 ;
        RECT 1551.265 137.445 1551.435 137.615 ;
      LAYER met1 ;
        RECT 1550.730 434.760 1551.050 434.820 ;
        RECT 1550.535 434.620 1551.050 434.760 ;
        RECT 1550.730 434.560 1551.050 434.620 ;
        RECT 1550.745 400.080 1551.035 400.125 ;
        RECT 1551.190 400.080 1551.510 400.140 ;
        RECT 1550.745 399.940 1551.510 400.080 ;
        RECT 1550.745 399.895 1551.035 399.940 ;
        RECT 1551.190 399.880 1551.510 399.940 ;
        RECT 1550.270 332.080 1550.590 332.140 ;
        RECT 1551.190 332.080 1551.510 332.140 ;
        RECT 1550.270 331.940 1551.510 332.080 ;
        RECT 1550.270 331.880 1550.590 331.940 ;
        RECT 1551.190 331.880 1551.510 331.940 ;
        RECT 1550.270 317.460 1550.590 317.520 ;
        RECT 1551.205 317.460 1551.495 317.505 ;
        RECT 1550.270 317.320 1551.495 317.460 ;
        RECT 1550.270 317.260 1550.590 317.320 ;
        RECT 1551.205 317.275 1551.495 317.320 ;
        RECT 1551.190 296.040 1551.510 296.100 ;
        RECT 1550.995 295.900 1551.510 296.040 ;
        RECT 1551.190 295.840 1551.510 295.900 ;
        RECT 1550.270 227.700 1550.590 227.760 ;
        RECT 1551.205 227.700 1551.495 227.745 ;
        RECT 1550.270 227.560 1551.495 227.700 ;
        RECT 1550.270 227.500 1550.590 227.560 ;
        RECT 1551.205 227.515 1551.495 227.560 ;
        RECT 1551.190 203.560 1551.510 203.620 ;
        RECT 1550.995 203.420 1551.510 203.560 ;
        RECT 1551.190 203.360 1551.510 203.420 ;
        RECT 1551.190 159.020 1551.510 159.080 ;
        RECT 1550.820 158.880 1551.510 159.020 ;
        RECT 1550.820 158.740 1550.960 158.880 ;
        RECT 1551.190 158.820 1551.510 158.880 ;
        RECT 1550.730 158.480 1551.050 158.740 ;
        RECT 1550.270 137.600 1550.590 137.660 ;
        RECT 1551.205 137.600 1551.495 137.645 ;
        RECT 1550.270 137.460 1551.495 137.600 ;
        RECT 1550.270 137.400 1550.590 137.460 ;
        RECT 1551.205 137.415 1551.495 137.460 ;
        RECT 1551.205 61.780 1551.495 61.825 ;
        RECT 1551.650 61.780 1551.970 61.840 ;
        RECT 1551.205 61.640 1551.970 61.780 ;
        RECT 1551.205 61.595 1551.495 61.640 ;
        RECT 1551.650 61.580 1551.970 61.640 ;
        RECT 1551.190 24.380 1551.510 24.440 ;
        RECT 1590.290 24.380 1590.610 24.440 ;
        RECT 1551.190 24.240 1590.610 24.380 ;
        RECT 1551.190 24.180 1551.510 24.240 ;
        RECT 1590.290 24.180 1590.610 24.240 ;
      LAYER via ;
        RECT 1550.760 434.560 1551.020 434.820 ;
        RECT 1551.220 399.880 1551.480 400.140 ;
        RECT 1550.300 331.880 1550.560 332.140 ;
        RECT 1551.220 331.880 1551.480 332.140 ;
        RECT 1550.300 317.260 1550.560 317.520 ;
        RECT 1551.220 295.840 1551.480 296.100 ;
        RECT 1550.300 227.500 1550.560 227.760 ;
        RECT 1551.220 203.360 1551.480 203.620 ;
        RECT 1551.220 158.820 1551.480 159.080 ;
        RECT 1550.760 158.480 1551.020 158.740 ;
        RECT 1550.300 137.400 1550.560 137.660 ;
        RECT 1551.680 61.580 1551.940 61.840 ;
        RECT 1551.220 24.180 1551.480 24.440 ;
        RECT 1590.320 24.180 1590.580 24.440 ;
      LAYER met2 ;
        RECT 1551.350 510.410 1551.630 514.000 ;
        RECT 1550.820 510.270 1551.630 510.410 ;
        RECT 1550.820 483.325 1550.960 510.270 ;
        RECT 1551.350 510.000 1551.630 510.270 ;
        RECT 1550.750 482.955 1551.030 483.325 ;
        RECT 1551.670 482.955 1551.950 483.325 ;
        RECT 1551.740 448.530 1551.880 482.955 ;
        RECT 1550.820 448.390 1551.880 448.530 ;
        RECT 1550.820 434.850 1550.960 448.390 ;
        RECT 1550.760 434.530 1551.020 434.850 ;
        RECT 1551.220 399.850 1551.480 400.170 ;
        RECT 1551.280 332.170 1551.420 399.850 ;
        RECT 1550.300 331.850 1550.560 332.170 ;
        RECT 1551.220 331.850 1551.480 332.170 ;
        RECT 1550.360 317.550 1550.500 331.850 ;
        RECT 1550.300 317.230 1550.560 317.550 ;
        RECT 1551.220 295.810 1551.480 296.130 ;
        RECT 1551.280 228.210 1551.420 295.810 ;
        RECT 1550.360 228.070 1551.420 228.210 ;
        RECT 1550.360 227.790 1550.500 228.070 ;
        RECT 1550.300 227.470 1550.560 227.790 ;
        RECT 1551.220 203.330 1551.480 203.650 ;
        RECT 1551.280 159.110 1551.420 203.330 ;
        RECT 1551.220 158.790 1551.480 159.110 ;
        RECT 1550.760 158.450 1551.020 158.770 ;
        RECT 1550.820 137.770 1550.960 158.450 ;
        RECT 1550.360 137.690 1550.960 137.770 ;
        RECT 1550.300 137.630 1550.960 137.690 ;
        RECT 1550.300 137.370 1550.560 137.630 ;
        RECT 1551.680 61.550 1551.940 61.870 ;
        RECT 1551.740 48.010 1551.880 61.550 ;
        RECT 1551.280 47.870 1551.880 48.010 ;
        RECT 1551.280 24.470 1551.420 47.870 ;
        RECT 1551.220 24.150 1551.480 24.470 ;
        RECT 1590.320 24.150 1590.580 24.470 ;
        RECT 1590.380 2.400 1590.520 24.150 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
      LAYER via2 ;
        RECT 1550.750 483.000 1551.030 483.280 ;
        RECT 1551.670 483.000 1551.950 483.280 ;
      LAYER met3 ;
        RECT 1550.725 483.290 1551.055 483.305 ;
        RECT 1551.645 483.290 1551.975 483.305 ;
        RECT 1550.725 482.990 1551.975 483.290 ;
        RECT 1550.725 482.975 1551.055 482.990 ;
        RECT 1551.645 482.975 1551.975 482.990 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 17.920 1566.230 17.980 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1565.910 17.780 1608.550 17.920 ;
        RECT 1565.910 17.720 1566.230 17.780 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
      LAYER via ;
        RECT 1565.940 17.720 1566.200 17.980 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
      LAYER met2 ;
        RECT 1564.230 510.410 1564.510 514.000 ;
        RECT 1564.230 510.270 1566.140 510.410 ;
        RECT 1564.230 510.000 1564.510 510.270 ;
        RECT 1566.000 18.010 1566.140 510.270 ;
        RECT 1565.940 17.690 1566.200 18.010 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1608.320 2.400 1608.460 17.690 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 17.580 1580.030 17.640 ;
        RECT 1626.170 17.580 1626.490 17.640 ;
        RECT 1579.710 17.440 1626.490 17.580 ;
        RECT 1579.710 17.380 1580.030 17.440 ;
        RECT 1626.170 17.380 1626.490 17.440 ;
      LAYER via ;
        RECT 1579.740 17.380 1580.000 17.640 ;
        RECT 1626.200 17.380 1626.460 17.640 ;
      LAYER met2 ;
        RECT 1577.110 510.410 1577.390 514.000 ;
        RECT 1577.110 510.270 1579.940 510.410 ;
        RECT 1577.110 510.000 1577.390 510.270 ;
        RECT 1579.800 17.670 1579.940 510.270 ;
        RECT 1579.740 17.350 1580.000 17.670 ;
        RECT 1626.200 17.350 1626.460 17.670 ;
        RECT 1626.260 2.400 1626.400 17.350 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1589.370 503.440 1589.690 503.500 ;
        RECT 1593.510 503.440 1593.830 503.500 ;
        RECT 1589.370 503.300 1593.830 503.440 ;
        RECT 1589.370 503.240 1589.690 503.300 ;
        RECT 1593.510 503.240 1593.830 503.300 ;
        RECT 1593.510 18.600 1593.830 18.660 ;
        RECT 1644.110 18.600 1644.430 18.660 ;
        RECT 1593.510 18.460 1644.430 18.600 ;
        RECT 1593.510 18.400 1593.830 18.460 ;
        RECT 1644.110 18.400 1644.430 18.460 ;
      LAYER via ;
        RECT 1589.400 503.240 1589.660 503.500 ;
        RECT 1593.540 503.240 1593.800 503.500 ;
        RECT 1593.540 18.400 1593.800 18.660 ;
        RECT 1644.140 18.400 1644.400 18.660 ;
      LAYER met2 ;
        RECT 1589.530 510.340 1589.810 514.000 ;
        RECT 1589.460 510.000 1589.810 510.340 ;
        RECT 1589.460 503.530 1589.600 510.000 ;
        RECT 1589.400 503.210 1589.660 503.530 ;
        RECT 1593.540 503.210 1593.800 503.530 ;
        RECT 1593.600 18.690 1593.740 503.210 ;
        RECT 1593.540 18.370 1593.800 18.690 ;
        RECT 1644.140 18.370 1644.400 18.690 ;
        RECT 1644.200 2.400 1644.340 18.370 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1602.250 476.580 1602.570 476.640 ;
        RECT 1607.310 476.580 1607.630 476.640 ;
        RECT 1602.250 476.440 1607.630 476.580 ;
        RECT 1602.250 476.380 1602.570 476.440 ;
        RECT 1607.310 476.380 1607.630 476.440 ;
        RECT 1607.310 19.960 1607.630 20.020 ;
        RECT 1662.050 19.960 1662.370 20.020 ;
        RECT 1607.310 19.820 1662.370 19.960 ;
        RECT 1607.310 19.760 1607.630 19.820 ;
        RECT 1662.050 19.760 1662.370 19.820 ;
      LAYER via ;
        RECT 1602.280 476.380 1602.540 476.640 ;
        RECT 1607.340 476.380 1607.600 476.640 ;
        RECT 1607.340 19.760 1607.600 20.020 ;
        RECT 1662.080 19.760 1662.340 20.020 ;
      LAYER met2 ;
        RECT 1602.410 510.340 1602.690 514.000 ;
        RECT 1602.340 510.000 1602.690 510.340 ;
        RECT 1602.340 476.670 1602.480 510.000 ;
        RECT 1602.280 476.350 1602.540 476.670 ;
        RECT 1607.340 476.350 1607.600 476.670 ;
        RECT 1607.400 20.050 1607.540 476.350 ;
        RECT 1607.340 19.730 1607.600 20.050 ;
        RECT 1662.080 19.730 1662.340 20.050 ;
        RECT 1662.140 2.400 1662.280 19.730 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.130 503.440 1615.450 503.500 ;
        RECT 1621.110 503.440 1621.430 503.500 ;
        RECT 1615.130 503.300 1621.430 503.440 ;
        RECT 1615.130 503.240 1615.450 503.300 ;
        RECT 1621.110 503.240 1621.430 503.300 ;
        RECT 1621.110 19.620 1621.430 19.680 ;
        RECT 1679.530 19.620 1679.850 19.680 ;
        RECT 1621.110 19.480 1679.850 19.620 ;
        RECT 1621.110 19.420 1621.430 19.480 ;
        RECT 1679.530 19.420 1679.850 19.480 ;
      LAYER via ;
        RECT 1615.160 503.240 1615.420 503.500 ;
        RECT 1621.140 503.240 1621.400 503.500 ;
        RECT 1621.140 19.420 1621.400 19.680 ;
        RECT 1679.560 19.420 1679.820 19.680 ;
      LAYER met2 ;
        RECT 1615.290 510.340 1615.570 514.000 ;
        RECT 1615.220 510.000 1615.570 510.340 ;
        RECT 1615.220 503.530 1615.360 510.000 ;
        RECT 1615.160 503.210 1615.420 503.530 ;
        RECT 1621.140 503.210 1621.400 503.530 ;
        RECT 1621.200 19.710 1621.340 503.210 ;
        RECT 1621.140 19.390 1621.400 19.710 ;
        RECT 1679.560 19.390 1679.820 19.710 ;
        RECT 1679.620 2.400 1679.760 19.390 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 17.240 1628.330 17.300 ;
        RECT 1697.470 17.240 1697.790 17.300 ;
        RECT 1628.010 17.100 1697.790 17.240 ;
        RECT 1628.010 17.040 1628.330 17.100 ;
        RECT 1697.470 17.040 1697.790 17.100 ;
      LAYER via ;
        RECT 1628.040 17.040 1628.300 17.300 ;
        RECT 1697.500 17.040 1697.760 17.300 ;
      LAYER met2 ;
        RECT 1628.170 510.340 1628.450 514.000 ;
        RECT 1628.100 510.000 1628.450 510.340 ;
        RECT 1628.100 17.330 1628.240 510.000 ;
        RECT 1628.040 17.010 1628.300 17.330 ;
        RECT 1697.500 17.010 1697.760 17.330 ;
        RECT 1697.560 2.400 1697.700 17.010 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 217.160 738.230 217.220 ;
        RECT 932.030 217.160 932.350 217.220 ;
        RECT 737.910 217.020 932.350 217.160 ;
        RECT 737.910 216.960 738.230 217.020 ;
        RECT 932.030 216.960 932.350 217.020 ;
        RECT 734.230 17.580 734.550 17.640 ;
        RECT 737.910 17.580 738.230 17.640 ;
        RECT 734.230 17.440 738.230 17.580 ;
        RECT 734.230 17.380 734.550 17.440 ;
        RECT 737.910 17.380 738.230 17.440 ;
      LAYER via ;
        RECT 737.940 216.960 738.200 217.220 ;
        RECT 932.060 216.960 932.320 217.220 ;
        RECT 734.260 17.380 734.520 17.640 ;
        RECT 737.940 17.380 738.200 17.640 ;
      LAYER met2 ;
        RECT 936.790 511.090 937.070 514.000 ;
        RECT 933.040 510.950 937.070 511.090 ;
        RECT 933.040 490.010 933.180 510.950 ;
        RECT 936.790 510.000 937.070 510.950 ;
        RECT 932.120 489.870 933.180 490.010 ;
        RECT 932.120 217.250 932.260 489.870 ;
        RECT 737.940 216.930 738.200 217.250 ;
        RECT 932.060 216.930 932.320 217.250 ;
        RECT 738.000 17.670 738.140 216.930 ;
        RECT 734.260 17.350 734.520 17.670 ;
        RECT 737.940 17.350 738.200 17.670 ;
        RECT 734.320 2.400 734.460 17.350 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1640.045 331.245 1640.215 379.355 ;
        RECT 1640.045 282.965 1640.215 330.735 ;
        RECT 1639.585 131.665 1639.755 158.695 ;
        RECT 1640.505 109.565 1640.675 131.155 ;
      LAYER mcon ;
        RECT 1640.045 379.185 1640.215 379.355 ;
        RECT 1640.045 330.565 1640.215 330.735 ;
        RECT 1639.585 158.525 1639.755 158.695 ;
        RECT 1640.505 130.985 1640.675 131.155 ;
      LAYER met1 ;
        RECT 1640.890 483.040 1641.210 483.100 ;
        RECT 1641.350 483.040 1641.670 483.100 ;
        RECT 1640.890 482.900 1641.670 483.040 ;
        RECT 1640.890 482.840 1641.210 482.900 ;
        RECT 1641.350 482.840 1641.670 482.900 ;
        RECT 1639.970 400.220 1640.290 400.480 ;
        RECT 1640.060 399.740 1640.200 400.220 ;
        RECT 1640.430 399.740 1640.750 399.800 ;
        RECT 1640.060 399.600 1640.750 399.740 ;
        RECT 1640.430 399.540 1640.750 399.600 ;
        RECT 1639.985 379.340 1640.275 379.385 ;
        RECT 1640.430 379.340 1640.750 379.400 ;
        RECT 1639.985 379.200 1640.750 379.340 ;
        RECT 1639.985 379.155 1640.275 379.200 ;
        RECT 1640.430 379.140 1640.750 379.200 ;
        RECT 1639.970 331.400 1640.290 331.460 ;
        RECT 1639.775 331.260 1640.290 331.400 ;
        RECT 1639.970 331.200 1640.290 331.260 ;
        RECT 1639.970 330.720 1640.290 330.780 ;
        RECT 1639.775 330.580 1640.290 330.720 ;
        RECT 1639.970 330.520 1640.290 330.580 ;
        RECT 1639.970 283.120 1640.290 283.180 ;
        RECT 1639.775 282.980 1640.290 283.120 ;
        RECT 1639.970 282.920 1640.290 282.980 ;
        RECT 1639.510 235.180 1639.830 235.240 ;
        RECT 1639.970 235.180 1640.290 235.240 ;
        RECT 1639.510 235.040 1640.290 235.180 ;
        RECT 1639.510 234.980 1639.830 235.040 ;
        RECT 1639.970 234.980 1640.290 235.040 ;
        RECT 1639.970 227.700 1640.290 227.760 ;
        RECT 1640.430 227.700 1640.750 227.760 ;
        RECT 1639.970 227.560 1640.750 227.700 ;
        RECT 1639.970 227.500 1640.290 227.560 ;
        RECT 1640.430 227.500 1640.750 227.560 ;
        RECT 1639.525 158.680 1639.815 158.725 ;
        RECT 1640.430 158.680 1640.750 158.740 ;
        RECT 1639.525 158.540 1640.750 158.680 ;
        RECT 1639.525 158.495 1639.815 158.540 ;
        RECT 1640.430 158.480 1640.750 158.540 ;
        RECT 1639.510 131.820 1639.830 131.880 ;
        RECT 1639.315 131.680 1639.830 131.820 ;
        RECT 1639.510 131.620 1639.830 131.680 ;
        RECT 1639.510 131.140 1639.830 131.200 ;
        RECT 1640.445 131.140 1640.735 131.185 ;
        RECT 1639.510 131.000 1640.735 131.140 ;
        RECT 1639.510 130.940 1639.830 131.000 ;
        RECT 1640.445 130.955 1640.735 131.000 ;
        RECT 1640.430 109.720 1640.750 109.780 ;
        RECT 1640.235 109.580 1640.750 109.720 ;
        RECT 1640.430 109.520 1640.750 109.580 ;
        RECT 1640.430 48.660 1640.750 48.920 ;
        RECT 1640.520 48.240 1640.660 48.660 ;
        RECT 1640.430 47.980 1640.750 48.240 ;
        RECT 1640.430 18.940 1640.750 19.000 ;
        RECT 1715.410 18.940 1715.730 19.000 ;
        RECT 1640.430 18.800 1715.730 18.940 ;
        RECT 1640.430 18.740 1640.750 18.800 ;
        RECT 1715.410 18.740 1715.730 18.800 ;
      LAYER via ;
        RECT 1640.920 482.840 1641.180 483.100 ;
        RECT 1641.380 482.840 1641.640 483.100 ;
        RECT 1640.000 400.220 1640.260 400.480 ;
        RECT 1640.460 399.540 1640.720 399.800 ;
        RECT 1640.460 379.140 1640.720 379.400 ;
        RECT 1640.000 331.200 1640.260 331.460 ;
        RECT 1640.000 330.520 1640.260 330.780 ;
        RECT 1640.000 282.920 1640.260 283.180 ;
        RECT 1639.540 234.980 1639.800 235.240 ;
        RECT 1640.000 234.980 1640.260 235.240 ;
        RECT 1640.000 227.500 1640.260 227.760 ;
        RECT 1640.460 227.500 1640.720 227.760 ;
        RECT 1640.460 158.480 1640.720 158.740 ;
        RECT 1639.540 131.620 1639.800 131.880 ;
        RECT 1639.540 130.940 1639.800 131.200 ;
        RECT 1640.460 109.520 1640.720 109.780 ;
        RECT 1640.460 48.660 1640.720 48.920 ;
        RECT 1640.460 47.980 1640.720 48.240 ;
        RECT 1640.460 18.740 1640.720 19.000 ;
        RECT 1715.440 18.740 1715.700 19.000 ;
      LAYER met2 ;
        RECT 1641.050 510.410 1641.330 514.000 ;
        RECT 1640.520 510.270 1641.330 510.410 ;
        RECT 1640.520 483.325 1640.660 510.270 ;
        RECT 1641.050 510.000 1641.330 510.270 ;
        RECT 1640.450 482.955 1640.730 483.325 ;
        RECT 1640.920 482.810 1641.180 483.130 ;
        RECT 1641.370 482.955 1641.650 483.325 ;
        RECT 1641.380 482.810 1641.640 482.955 ;
        RECT 1640.980 435.045 1641.120 482.810 ;
        RECT 1639.990 434.675 1640.270 435.045 ;
        RECT 1640.910 434.675 1641.190 435.045 ;
        RECT 1640.060 400.510 1640.200 434.675 ;
        RECT 1640.000 400.190 1640.260 400.510 ;
        RECT 1640.460 399.510 1640.720 399.830 ;
        RECT 1640.520 379.430 1640.660 399.510 ;
        RECT 1640.460 379.110 1640.720 379.430 ;
        RECT 1640.000 331.170 1640.260 331.490 ;
        RECT 1640.060 330.810 1640.200 331.170 ;
        RECT 1640.000 330.490 1640.260 330.810 ;
        RECT 1640.000 282.890 1640.260 283.210 ;
        RECT 1640.060 255.410 1640.200 282.890 ;
        RECT 1639.600 255.270 1640.200 255.410 ;
        RECT 1639.600 235.270 1639.740 255.270 ;
        RECT 1639.540 234.950 1639.800 235.270 ;
        RECT 1640.000 234.950 1640.260 235.270 ;
        RECT 1640.060 227.790 1640.200 234.950 ;
        RECT 1640.000 227.470 1640.260 227.790 ;
        RECT 1640.460 227.470 1640.720 227.790 ;
        RECT 1640.520 158.770 1640.660 227.470 ;
        RECT 1640.460 158.450 1640.720 158.770 ;
        RECT 1639.540 131.590 1639.800 131.910 ;
        RECT 1639.600 131.230 1639.740 131.590 ;
        RECT 1639.540 130.910 1639.800 131.230 ;
        RECT 1640.460 109.490 1640.720 109.810 ;
        RECT 1640.520 48.950 1640.660 109.490 ;
        RECT 1640.460 48.630 1640.720 48.950 ;
        RECT 1640.460 47.950 1640.720 48.270 ;
        RECT 1640.520 19.030 1640.660 47.950 ;
        RECT 1640.460 18.710 1640.720 19.030 ;
        RECT 1715.440 18.710 1715.700 19.030 ;
        RECT 1715.500 2.400 1715.640 18.710 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
      LAYER via2 ;
        RECT 1640.450 483.000 1640.730 483.280 ;
        RECT 1641.370 483.000 1641.650 483.280 ;
        RECT 1639.990 434.720 1640.270 435.000 ;
        RECT 1640.910 434.720 1641.190 435.000 ;
      LAYER met3 ;
        RECT 1640.425 483.290 1640.755 483.305 ;
        RECT 1641.345 483.290 1641.675 483.305 ;
        RECT 1640.425 482.990 1641.675 483.290 ;
        RECT 1640.425 482.975 1640.755 482.990 ;
        RECT 1641.345 482.975 1641.675 482.990 ;
        RECT 1639.965 435.010 1640.295 435.025 ;
        RECT 1640.885 435.010 1641.215 435.025 ;
        RECT 1639.965 434.710 1641.215 435.010 ;
        RECT 1639.965 434.695 1640.295 434.710 ;
        RECT 1640.885 434.695 1641.215 434.710 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.610 18.600 1655.930 18.660 ;
        RECT 1733.350 18.600 1733.670 18.660 ;
        RECT 1655.610 18.460 1733.670 18.600 ;
        RECT 1655.610 18.400 1655.930 18.460 ;
        RECT 1733.350 18.400 1733.670 18.460 ;
      LAYER via ;
        RECT 1655.640 18.400 1655.900 18.660 ;
        RECT 1733.380 18.400 1733.640 18.660 ;
      LAYER met2 ;
        RECT 1653.930 510.410 1654.210 514.000 ;
        RECT 1653.930 510.270 1655.840 510.410 ;
        RECT 1653.930 510.000 1654.210 510.270 ;
        RECT 1655.700 18.690 1655.840 510.270 ;
        RECT 1655.640 18.370 1655.900 18.690 ;
        RECT 1733.380 18.370 1733.640 18.690 ;
        RECT 1733.440 2.400 1733.580 18.370 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.410 18.260 1669.730 18.320 ;
        RECT 1751.290 18.260 1751.610 18.320 ;
        RECT 1669.410 18.120 1751.610 18.260 ;
        RECT 1669.410 18.060 1669.730 18.120 ;
        RECT 1751.290 18.060 1751.610 18.120 ;
      LAYER via ;
        RECT 1669.440 18.060 1669.700 18.320 ;
        RECT 1751.320 18.060 1751.580 18.320 ;
      LAYER met2 ;
        RECT 1666.350 510.410 1666.630 514.000 ;
        RECT 1666.350 510.270 1669.640 510.410 ;
        RECT 1666.350 510.000 1666.630 510.270 ;
        RECT 1669.500 18.350 1669.640 510.270 ;
        RECT 1669.440 18.030 1669.700 18.350 ;
        RECT 1751.320 18.030 1751.580 18.350 ;
        RECT 1751.380 2.400 1751.520 18.030 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1738.485 16.745 1738.655 17.935 ;
      LAYER mcon ;
        RECT 1738.485 17.765 1738.655 17.935 ;
      LAYER met1 ;
        RECT 1679.070 503.440 1679.390 503.500 ;
        RECT 1682.750 503.440 1683.070 503.500 ;
        RECT 1679.070 503.300 1683.070 503.440 ;
        RECT 1679.070 503.240 1679.390 503.300 ;
        RECT 1682.750 503.240 1683.070 503.300 ;
        RECT 1682.750 17.920 1683.070 17.980 ;
        RECT 1738.425 17.920 1738.715 17.965 ;
        RECT 1682.750 17.780 1738.715 17.920 ;
        RECT 1682.750 17.720 1683.070 17.780 ;
        RECT 1738.425 17.735 1738.715 17.780 ;
        RECT 1738.425 16.900 1738.715 16.945 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1738.425 16.760 1769.090 16.900 ;
        RECT 1738.425 16.715 1738.715 16.760 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
      LAYER via ;
        RECT 1679.100 503.240 1679.360 503.500 ;
        RECT 1682.780 503.240 1683.040 503.500 ;
        RECT 1682.780 17.720 1683.040 17.980 ;
        RECT 1768.800 16.700 1769.060 16.960 ;
      LAYER met2 ;
        RECT 1679.230 510.340 1679.510 514.000 ;
        RECT 1679.160 510.000 1679.510 510.340 ;
        RECT 1679.160 503.530 1679.300 510.000 ;
        RECT 1679.100 503.210 1679.360 503.530 ;
        RECT 1682.780 503.210 1683.040 503.530 ;
        RECT 1682.840 18.010 1682.980 503.210 ;
        RECT 1682.780 17.690 1683.040 18.010 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1691.950 503.440 1692.270 503.500 ;
        RECT 1697.010 503.440 1697.330 503.500 ;
        RECT 1691.950 503.300 1697.330 503.440 ;
        RECT 1691.950 503.240 1692.270 503.300 ;
        RECT 1697.010 503.240 1697.330 503.300 ;
        RECT 1697.010 17.580 1697.330 17.640 ;
        RECT 1786.710 17.580 1787.030 17.640 ;
        RECT 1697.010 17.440 1787.030 17.580 ;
        RECT 1697.010 17.380 1697.330 17.440 ;
        RECT 1786.710 17.380 1787.030 17.440 ;
      LAYER via ;
        RECT 1691.980 503.240 1692.240 503.500 ;
        RECT 1697.040 503.240 1697.300 503.500 ;
        RECT 1697.040 17.380 1697.300 17.640 ;
        RECT 1786.740 17.380 1787.000 17.640 ;
      LAYER met2 ;
        RECT 1692.110 510.340 1692.390 514.000 ;
        RECT 1692.040 510.000 1692.390 510.340 ;
        RECT 1692.040 503.530 1692.180 510.000 ;
        RECT 1691.980 503.210 1692.240 503.530 ;
        RECT 1697.040 503.210 1697.300 503.530 ;
        RECT 1697.100 17.670 1697.240 503.210 ;
        RECT 1697.040 17.350 1697.300 17.670 ;
        RECT 1786.740 17.350 1787.000 17.670 ;
        RECT 1786.800 2.400 1786.940 17.350 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1704.830 503.100 1705.150 503.160 ;
        RECT 1710.810 503.100 1711.130 503.160 ;
        RECT 1704.830 502.960 1711.130 503.100 ;
        RECT 1704.830 502.900 1705.150 502.960 ;
        RECT 1710.810 502.900 1711.130 502.960 ;
        RECT 1710.810 17.240 1711.130 17.300 ;
        RECT 1804.650 17.240 1804.970 17.300 ;
        RECT 1710.810 17.100 1804.970 17.240 ;
        RECT 1710.810 17.040 1711.130 17.100 ;
        RECT 1804.650 17.040 1804.970 17.100 ;
      LAYER via ;
        RECT 1704.860 502.900 1705.120 503.160 ;
        RECT 1710.840 502.900 1711.100 503.160 ;
        RECT 1710.840 17.040 1711.100 17.300 ;
        RECT 1804.680 17.040 1804.940 17.300 ;
      LAYER met2 ;
        RECT 1704.990 510.340 1705.270 514.000 ;
        RECT 1704.920 510.000 1705.270 510.340 ;
        RECT 1704.920 503.190 1705.060 510.000 ;
        RECT 1704.860 502.870 1705.120 503.190 ;
        RECT 1710.840 502.870 1711.100 503.190 ;
        RECT 1710.900 17.330 1711.040 502.870 ;
        RECT 1710.840 17.010 1711.100 17.330 ;
        RECT 1804.680 17.010 1804.940 17.330 ;
        RECT 1804.740 2.400 1804.880 17.010 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 19.620 1718.030 19.680 ;
        RECT 1822.590 19.620 1822.910 19.680 ;
        RECT 1717.710 19.480 1822.910 19.620 ;
        RECT 1717.710 19.420 1718.030 19.480 ;
        RECT 1822.590 19.420 1822.910 19.480 ;
      LAYER via ;
        RECT 1717.740 19.420 1718.000 19.680 ;
        RECT 1822.620 19.420 1822.880 19.680 ;
      LAYER met2 ;
        RECT 1717.870 510.340 1718.150 514.000 ;
        RECT 1717.800 510.000 1718.150 510.340 ;
        RECT 1717.800 19.710 1717.940 510.000 ;
        RECT 1717.740 19.390 1718.000 19.710 ;
        RECT 1822.620 19.390 1822.880 19.710 ;
        RECT 1822.680 2.400 1822.820 19.390 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.510 19.960 1731.830 20.020 ;
        RECT 1840.070 19.960 1840.390 20.020 ;
        RECT 1731.510 19.820 1840.390 19.960 ;
        RECT 1731.510 19.760 1731.830 19.820 ;
        RECT 1840.070 19.760 1840.390 19.820 ;
      LAYER via ;
        RECT 1731.540 19.760 1731.800 20.020 ;
        RECT 1840.100 19.760 1840.360 20.020 ;
      LAYER met2 ;
        RECT 1730.750 510.410 1731.030 514.000 ;
        RECT 1730.750 510.270 1731.740 510.410 ;
        RECT 1730.750 510.000 1731.030 510.270 ;
        RECT 1731.600 20.050 1731.740 510.270 ;
        RECT 1731.540 19.730 1731.800 20.050 ;
        RECT 1840.100 19.730 1840.360 20.050 ;
        RECT 1840.160 2.400 1840.300 19.730 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1858.010 19.620 1858.330 19.680 ;
        RECT 1828.200 19.480 1858.330 19.620 ;
        RECT 1745.310 19.280 1745.630 19.340 ;
        RECT 1828.200 19.280 1828.340 19.480 ;
        RECT 1858.010 19.420 1858.330 19.480 ;
        RECT 1745.310 19.140 1828.340 19.280 ;
        RECT 1745.310 19.080 1745.630 19.140 ;
      LAYER via ;
        RECT 1745.340 19.080 1745.600 19.340 ;
        RECT 1858.040 19.420 1858.300 19.680 ;
      LAYER met2 ;
        RECT 1743.170 510.410 1743.450 514.000 ;
        RECT 1743.170 510.270 1745.540 510.410 ;
        RECT 1743.170 510.000 1743.450 510.270 ;
        RECT 1745.400 19.370 1745.540 510.270 ;
        RECT 1858.040 19.390 1858.300 19.710 ;
        RECT 1745.340 19.050 1745.600 19.370 ;
        RECT 1858.100 2.400 1858.240 19.390 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 18.940 1759.430 19.000 ;
        RECT 1875.950 18.940 1876.270 19.000 ;
        RECT 1759.110 18.800 1876.270 18.940 ;
        RECT 1759.110 18.740 1759.430 18.800 ;
        RECT 1875.950 18.740 1876.270 18.800 ;
      LAYER via ;
        RECT 1759.140 18.740 1759.400 19.000 ;
        RECT 1875.980 18.740 1876.240 19.000 ;
      LAYER met2 ;
        RECT 1756.050 510.410 1756.330 514.000 ;
        RECT 1756.050 510.270 1759.340 510.410 ;
        RECT 1756.050 510.000 1756.330 510.270 ;
        RECT 1759.200 19.030 1759.340 510.270 ;
        RECT 1759.140 18.710 1759.400 19.030 ;
        RECT 1875.980 18.710 1876.240 19.030 ;
        RECT 1876.040 2.400 1876.180 18.710 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 224.300 758.930 224.360 ;
        RECT 945.370 224.300 945.690 224.360 ;
        RECT 758.610 224.160 945.690 224.300 ;
        RECT 758.610 224.100 758.930 224.160 ;
        RECT 945.370 224.100 945.690 224.160 ;
        RECT 752.170 17.580 752.490 17.640 ;
        RECT 758.610 17.580 758.930 17.640 ;
        RECT 752.170 17.440 758.930 17.580 ;
        RECT 752.170 17.380 752.490 17.440 ;
        RECT 758.610 17.380 758.930 17.440 ;
      LAYER via ;
        RECT 758.640 224.100 758.900 224.360 ;
        RECT 945.400 224.100 945.660 224.360 ;
        RECT 752.200 17.380 752.460 17.640 ;
        RECT 758.640 17.380 758.900 17.640 ;
      LAYER met2 ;
        RECT 949.670 511.090 949.950 514.000 ;
        RECT 945.920 510.950 949.950 511.090 ;
        RECT 945.920 490.010 946.060 510.950 ;
        RECT 949.670 510.000 949.950 510.950 ;
        RECT 945.460 489.870 946.060 490.010 ;
        RECT 945.460 224.390 945.600 489.870 ;
        RECT 758.640 224.070 758.900 224.390 ;
        RECT 945.400 224.070 945.660 224.390 ;
        RECT 758.700 17.670 758.840 224.070 ;
        RECT 752.200 17.350 752.460 17.670 ;
        RECT 758.640 17.350 758.900 17.670 ;
        RECT 752.260 2.400 752.400 17.350 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 503.440 1769.090 503.500 ;
        RECT 1772.910 503.440 1773.230 503.500 ;
        RECT 1768.770 503.300 1773.230 503.440 ;
        RECT 1768.770 503.240 1769.090 503.300 ;
        RECT 1772.910 503.240 1773.230 503.300 ;
        RECT 1772.910 18.600 1773.230 18.660 ;
        RECT 1893.890 18.600 1894.210 18.660 ;
        RECT 1772.910 18.460 1894.210 18.600 ;
        RECT 1772.910 18.400 1773.230 18.460 ;
        RECT 1893.890 18.400 1894.210 18.460 ;
      LAYER via ;
        RECT 1768.800 503.240 1769.060 503.500 ;
        RECT 1772.940 503.240 1773.200 503.500 ;
        RECT 1772.940 18.400 1773.200 18.660 ;
        RECT 1893.920 18.400 1894.180 18.660 ;
      LAYER met2 ;
        RECT 1768.930 510.340 1769.210 514.000 ;
        RECT 1768.860 510.000 1769.210 510.340 ;
        RECT 1768.860 503.530 1769.000 510.000 ;
        RECT 1768.800 503.210 1769.060 503.530 ;
        RECT 1772.940 503.210 1773.200 503.530 ;
        RECT 1773.000 18.690 1773.140 503.210 ;
        RECT 1772.940 18.370 1773.200 18.690 ;
        RECT 1893.920 18.370 1894.180 18.690 ;
        RECT 1893.980 2.400 1894.120 18.370 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1781.650 503.440 1781.970 503.500 ;
        RECT 1786.710 503.440 1787.030 503.500 ;
        RECT 1781.650 503.300 1787.030 503.440 ;
        RECT 1781.650 503.240 1781.970 503.300 ;
        RECT 1786.710 503.240 1787.030 503.300 ;
        RECT 1786.710 18.060 1787.030 18.320 ;
        RECT 1786.800 17.920 1786.940 18.060 ;
        RECT 1911.830 17.920 1912.150 17.980 ;
        RECT 1786.800 17.780 1912.150 17.920 ;
        RECT 1911.830 17.720 1912.150 17.780 ;
      LAYER via ;
        RECT 1781.680 503.240 1781.940 503.500 ;
        RECT 1786.740 503.240 1787.000 503.500 ;
        RECT 1786.740 18.060 1787.000 18.320 ;
        RECT 1911.860 17.720 1912.120 17.980 ;
      LAYER met2 ;
        RECT 1781.810 510.340 1782.090 514.000 ;
        RECT 1781.740 510.000 1782.090 510.340 ;
        RECT 1781.740 503.530 1781.880 510.000 ;
        RECT 1781.680 503.210 1781.940 503.530 ;
        RECT 1786.740 503.210 1787.000 503.530 ;
        RECT 1786.800 18.350 1786.940 503.210 ;
        RECT 1786.740 18.030 1787.000 18.350 ;
        RECT 1911.860 17.690 1912.120 18.010 ;
        RECT 1911.920 2.400 1912.060 17.690 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1794.530 499.360 1794.850 499.420 ;
        RECT 1800.510 499.360 1800.830 499.420 ;
        RECT 1794.530 499.220 1800.830 499.360 ;
        RECT 1794.530 499.160 1794.850 499.220 ;
        RECT 1800.510 499.160 1800.830 499.220 ;
        RECT 1800.510 18.260 1800.830 18.320 ;
        RECT 1929.310 18.260 1929.630 18.320 ;
        RECT 1800.510 18.120 1929.630 18.260 ;
        RECT 1800.510 18.060 1800.830 18.120 ;
        RECT 1929.310 18.060 1929.630 18.120 ;
      LAYER via ;
        RECT 1794.560 499.160 1794.820 499.420 ;
        RECT 1800.540 499.160 1800.800 499.420 ;
        RECT 1800.540 18.060 1800.800 18.320 ;
        RECT 1929.340 18.060 1929.600 18.320 ;
      LAYER met2 ;
        RECT 1794.690 510.340 1794.970 514.000 ;
        RECT 1794.620 510.000 1794.970 510.340 ;
        RECT 1794.620 499.450 1794.760 510.000 ;
        RECT 1794.560 499.130 1794.820 499.450 ;
        RECT 1800.540 499.130 1800.800 499.450 ;
        RECT 1800.600 18.350 1800.740 499.130 ;
        RECT 1800.540 18.030 1800.800 18.350 ;
        RECT 1929.340 18.030 1929.600 18.350 ;
        RECT 1929.400 2.400 1929.540 18.030 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.410 17.240 1807.730 17.300 ;
        RECT 1947.250 17.240 1947.570 17.300 ;
        RECT 1807.410 17.100 1947.570 17.240 ;
        RECT 1807.410 17.040 1807.730 17.100 ;
        RECT 1947.250 17.040 1947.570 17.100 ;
      LAYER via ;
        RECT 1807.440 17.040 1807.700 17.300 ;
        RECT 1947.280 17.040 1947.540 17.300 ;
      LAYER met2 ;
        RECT 1807.570 510.340 1807.850 514.000 ;
        RECT 1807.500 510.000 1807.850 510.340 ;
        RECT 1807.500 17.330 1807.640 510.000 ;
        RECT 1807.440 17.010 1807.700 17.330 ;
        RECT 1947.280 17.010 1947.540 17.330 ;
        RECT 1947.340 2.400 1947.480 17.010 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 17.580 1821.530 17.640 ;
        RECT 1965.190 17.580 1965.510 17.640 ;
        RECT 1821.210 17.440 1965.510 17.580 ;
        RECT 1821.210 17.380 1821.530 17.440 ;
        RECT 1965.190 17.380 1965.510 17.440 ;
      LAYER via ;
        RECT 1821.240 17.380 1821.500 17.640 ;
        RECT 1965.220 17.380 1965.480 17.640 ;
      LAYER met2 ;
        RECT 1819.990 510.410 1820.270 514.000 ;
        RECT 1819.990 510.270 1821.440 510.410 ;
        RECT 1819.990 510.000 1820.270 510.270 ;
        RECT 1821.300 17.670 1821.440 510.270 ;
        RECT 1821.240 17.350 1821.500 17.670 ;
        RECT 1965.220 17.350 1965.480 17.670 ;
        RECT 1965.280 2.400 1965.420 17.350 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1834.550 162.420 1834.870 162.480 ;
        RECT 1980.370 162.420 1980.690 162.480 ;
        RECT 1834.550 162.280 1980.690 162.420 ;
        RECT 1834.550 162.220 1834.870 162.280 ;
        RECT 1980.370 162.220 1980.690 162.280 ;
        RECT 1980.370 62.120 1980.690 62.180 ;
        RECT 1983.130 62.120 1983.450 62.180 ;
        RECT 1980.370 61.980 1983.450 62.120 ;
        RECT 1980.370 61.920 1980.690 61.980 ;
        RECT 1983.130 61.920 1983.450 61.980 ;
      LAYER via ;
        RECT 1834.580 162.220 1834.840 162.480 ;
        RECT 1980.400 162.220 1980.660 162.480 ;
        RECT 1980.400 61.920 1980.660 62.180 ;
        RECT 1983.160 61.920 1983.420 62.180 ;
      LAYER met2 ;
        RECT 1832.870 510.410 1833.150 514.000 ;
        RECT 1832.870 510.270 1834.780 510.410 ;
        RECT 1832.870 510.000 1833.150 510.270 ;
        RECT 1834.640 162.510 1834.780 510.270 ;
        RECT 1834.580 162.190 1834.840 162.510 ;
        RECT 1980.400 162.190 1980.660 162.510 ;
        RECT 1980.460 62.210 1980.600 162.190 ;
        RECT 1980.400 61.890 1980.660 62.210 ;
        RECT 1983.160 61.890 1983.420 62.210 ;
        RECT 1983.220 2.400 1983.360 61.890 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.810 183.160 1849.130 183.220 ;
        RECT 2001.070 183.160 2001.390 183.220 ;
        RECT 1848.810 183.020 2001.390 183.160 ;
        RECT 1848.810 182.960 1849.130 183.020 ;
        RECT 2001.070 182.960 2001.390 183.020 ;
      LAYER via ;
        RECT 1848.840 182.960 1849.100 183.220 ;
        RECT 2001.100 182.960 2001.360 183.220 ;
      LAYER met2 ;
        RECT 1845.750 510.410 1846.030 514.000 ;
        RECT 1845.750 510.270 1849.040 510.410 ;
        RECT 1845.750 510.000 1846.030 510.270 ;
        RECT 1848.900 183.250 1849.040 510.270 ;
        RECT 1848.840 182.930 1849.100 183.250 ;
        RECT 2001.100 182.930 2001.360 183.250 ;
        RECT 2001.160 2.400 2001.300 182.930 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1858.470 503.100 1858.790 503.160 ;
        RECT 1862.610 503.100 1862.930 503.160 ;
        RECT 1858.470 502.960 1862.930 503.100 ;
        RECT 1858.470 502.900 1858.790 502.960 ;
        RECT 1862.610 502.900 1862.930 502.960 ;
        RECT 1862.610 189.620 1862.930 189.680 ;
        RECT 2014.870 189.620 2015.190 189.680 ;
        RECT 1862.610 189.480 2015.190 189.620 ;
        RECT 1862.610 189.420 1862.930 189.480 ;
        RECT 2014.870 189.420 2015.190 189.480 ;
        RECT 2014.870 62.260 2015.190 62.520 ;
        RECT 2014.960 61.780 2015.100 62.260 ;
        RECT 2018.550 61.780 2018.870 61.840 ;
        RECT 2014.960 61.640 2018.870 61.780 ;
        RECT 2018.550 61.580 2018.870 61.640 ;
        RECT 2018.550 47.980 2018.870 48.240 ;
        RECT 2018.640 47.560 2018.780 47.980 ;
        RECT 2018.550 47.300 2018.870 47.560 ;
      LAYER via ;
        RECT 1858.500 502.900 1858.760 503.160 ;
        RECT 1862.640 502.900 1862.900 503.160 ;
        RECT 1862.640 189.420 1862.900 189.680 ;
        RECT 2014.900 189.420 2015.160 189.680 ;
        RECT 2014.900 62.260 2015.160 62.520 ;
        RECT 2018.580 61.580 2018.840 61.840 ;
        RECT 2018.580 47.980 2018.840 48.240 ;
        RECT 2018.580 47.300 2018.840 47.560 ;
      LAYER met2 ;
        RECT 1858.630 510.340 1858.910 514.000 ;
        RECT 1858.560 510.000 1858.910 510.340 ;
        RECT 1858.560 503.190 1858.700 510.000 ;
        RECT 1858.500 502.870 1858.760 503.190 ;
        RECT 1862.640 502.870 1862.900 503.190 ;
        RECT 1862.700 189.710 1862.840 502.870 ;
        RECT 1862.640 189.390 1862.900 189.710 ;
        RECT 2014.900 189.390 2015.160 189.710 ;
        RECT 2014.960 62.550 2015.100 189.390 ;
        RECT 2014.900 62.230 2015.160 62.550 ;
        RECT 2018.580 61.550 2018.840 61.870 ;
        RECT 2018.640 48.270 2018.780 61.550 ;
        RECT 2018.580 47.950 2018.840 48.270 ;
        RECT 2018.580 47.270 2018.840 47.590 ;
        RECT 2018.640 2.400 2018.780 47.270 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2036.565 2.805 2036.735 48.195 ;
      LAYER mcon ;
        RECT 2036.565 48.025 2036.735 48.195 ;
      LAYER met1 ;
        RECT 1871.350 503.440 1871.670 503.500 ;
        RECT 1875.950 503.440 1876.270 503.500 ;
        RECT 1871.350 503.300 1876.270 503.440 ;
        RECT 1871.350 503.240 1871.670 503.300 ;
        RECT 1875.950 503.240 1876.270 503.300 ;
        RECT 1875.950 210.360 1876.270 210.420 ;
        RECT 2035.570 210.360 2035.890 210.420 ;
        RECT 1875.950 210.220 2035.890 210.360 ;
        RECT 1875.950 210.160 1876.270 210.220 ;
        RECT 2035.570 210.160 2035.890 210.220 ;
        RECT 2036.490 48.180 2036.810 48.240 ;
        RECT 2036.295 48.040 2036.810 48.180 ;
        RECT 2036.490 47.980 2036.810 48.040 ;
        RECT 2036.490 2.960 2036.810 3.020 ;
        RECT 2036.295 2.820 2036.810 2.960 ;
        RECT 2036.490 2.760 2036.810 2.820 ;
      LAYER via ;
        RECT 1871.380 503.240 1871.640 503.500 ;
        RECT 1875.980 503.240 1876.240 503.500 ;
        RECT 1875.980 210.160 1876.240 210.420 ;
        RECT 2035.600 210.160 2035.860 210.420 ;
        RECT 2036.520 47.980 2036.780 48.240 ;
        RECT 2036.520 2.760 2036.780 3.020 ;
      LAYER met2 ;
        RECT 1871.510 510.340 1871.790 514.000 ;
        RECT 1871.440 510.000 1871.790 510.340 ;
        RECT 1871.440 503.530 1871.580 510.000 ;
        RECT 1871.380 503.210 1871.640 503.530 ;
        RECT 1875.980 503.210 1876.240 503.530 ;
        RECT 1876.040 210.450 1876.180 503.210 ;
        RECT 1875.980 210.130 1876.240 210.450 ;
        RECT 2035.600 210.130 2035.860 210.450 ;
        RECT 2035.660 62.120 2035.800 210.130 ;
        RECT 2035.660 61.980 2036.720 62.120 ;
        RECT 2036.580 48.270 2036.720 61.980 ;
        RECT 2036.520 47.950 2036.780 48.270 ;
        RECT 2036.520 2.730 2036.780 3.050 ;
        RECT 2036.580 2.400 2036.720 2.730 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1884.230 498.340 1884.550 498.400 ;
        RECT 1890.210 498.340 1890.530 498.400 ;
        RECT 1884.230 498.200 1890.530 498.340 ;
        RECT 1884.230 498.140 1884.550 498.200 ;
        RECT 1890.210 498.140 1890.530 498.200 ;
        RECT 1890.210 224.300 1890.530 224.360 ;
        RECT 2049.370 224.300 2049.690 224.360 ;
        RECT 1890.210 224.160 2049.690 224.300 ;
        RECT 1890.210 224.100 1890.530 224.160 ;
        RECT 2049.370 224.100 2049.690 224.160 ;
        RECT 2049.370 62.120 2049.690 62.180 ;
        RECT 2054.430 62.120 2054.750 62.180 ;
        RECT 2049.370 61.980 2054.750 62.120 ;
        RECT 2049.370 61.920 2049.690 61.980 ;
        RECT 2054.430 61.920 2054.750 61.980 ;
      LAYER via ;
        RECT 1884.260 498.140 1884.520 498.400 ;
        RECT 1890.240 498.140 1890.500 498.400 ;
        RECT 1890.240 224.100 1890.500 224.360 ;
        RECT 2049.400 224.100 2049.660 224.360 ;
        RECT 2049.400 61.920 2049.660 62.180 ;
        RECT 2054.460 61.920 2054.720 62.180 ;
      LAYER met2 ;
        RECT 1884.390 510.340 1884.670 514.000 ;
        RECT 1884.320 510.000 1884.670 510.340 ;
        RECT 1884.320 498.430 1884.460 510.000 ;
        RECT 1884.260 498.110 1884.520 498.430 ;
        RECT 1890.240 498.110 1890.500 498.430 ;
        RECT 1890.300 224.390 1890.440 498.110 ;
        RECT 1890.240 224.070 1890.500 224.390 ;
        RECT 2049.400 224.070 2049.660 224.390 ;
        RECT 2049.460 62.210 2049.600 224.070 ;
        RECT 2049.400 61.890 2049.660 62.210 ;
        RECT 2054.460 61.890 2054.720 62.210 ;
        RECT 2054.520 2.400 2054.660 61.890 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 231.100 772.730 231.160 ;
        RECT 959.170 231.100 959.490 231.160 ;
        RECT 772.410 230.960 959.490 231.100 ;
        RECT 772.410 230.900 772.730 230.960 ;
        RECT 959.170 230.900 959.490 230.960 ;
        RECT 769.650 20.640 769.970 20.700 ;
        RECT 772.410 20.640 772.730 20.700 ;
        RECT 769.650 20.500 772.730 20.640 ;
        RECT 769.650 20.440 769.970 20.500 ;
        RECT 772.410 20.440 772.730 20.500 ;
      LAYER via ;
        RECT 772.440 230.900 772.700 231.160 ;
        RECT 959.200 230.900 959.460 231.160 ;
        RECT 769.680 20.440 769.940 20.700 ;
        RECT 772.440 20.440 772.700 20.700 ;
      LAYER met2 ;
        RECT 962.090 510.410 962.370 514.000 ;
        RECT 959.260 510.270 962.370 510.410 ;
        RECT 959.260 231.190 959.400 510.270 ;
        RECT 962.090 510.000 962.370 510.270 ;
        RECT 772.440 230.870 772.700 231.190 ;
        RECT 959.200 230.870 959.460 231.190 ;
        RECT 772.500 20.730 772.640 230.870 ;
        RECT 769.680 20.410 769.940 20.730 ;
        RECT 772.440 20.410 772.700 20.730 ;
        RECT 769.740 2.400 769.880 20.410 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2072.445 2.805 2072.615 48.195 ;
      LAYER mcon ;
        RECT 2072.445 48.025 2072.615 48.195 ;
      LAYER met1 ;
        RECT 1896.190 448.700 1896.510 448.760 ;
        RECT 1897.110 448.700 1897.430 448.760 ;
        RECT 1896.190 448.560 1897.430 448.700 ;
        RECT 1896.190 448.500 1896.510 448.560 ;
        RECT 1897.110 448.500 1897.430 448.560 ;
        RECT 1896.650 400.560 1896.970 400.820 ;
        RECT 1896.740 400.140 1896.880 400.560 ;
        RECT 1896.650 399.880 1896.970 400.140 ;
        RECT 1896.190 237.900 1896.510 237.960 ;
        RECT 2070.070 237.900 2070.390 237.960 ;
        RECT 1896.190 237.760 2070.390 237.900 ;
        RECT 1896.190 237.700 1896.510 237.760 ;
        RECT 2070.070 237.700 2070.390 237.760 ;
        RECT 2070.070 62.120 2070.390 62.180 ;
        RECT 2072.370 62.120 2072.690 62.180 ;
        RECT 2070.070 61.980 2072.690 62.120 ;
        RECT 2070.070 61.920 2070.390 61.980 ;
        RECT 2072.370 61.920 2072.690 61.980 ;
        RECT 2072.370 48.180 2072.690 48.240 ;
        RECT 2072.175 48.040 2072.690 48.180 ;
        RECT 2072.370 47.980 2072.690 48.040 ;
        RECT 2072.370 2.960 2072.690 3.020 ;
        RECT 2072.175 2.820 2072.690 2.960 ;
        RECT 2072.370 2.760 2072.690 2.820 ;
      LAYER via ;
        RECT 1896.220 448.500 1896.480 448.760 ;
        RECT 1897.140 448.500 1897.400 448.760 ;
        RECT 1896.680 400.560 1896.940 400.820 ;
        RECT 1896.680 399.880 1896.940 400.140 ;
        RECT 1896.220 237.700 1896.480 237.960 ;
        RECT 2070.100 237.700 2070.360 237.960 ;
        RECT 2070.100 61.920 2070.360 62.180 ;
        RECT 2072.400 61.920 2072.660 62.180 ;
        RECT 2072.400 47.980 2072.660 48.240 ;
        RECT 2072.400 2.760 2072.660 3.020 ;
      LAYER met2 ;
        RECT 1896.810 510.410 1897.090 514.000 ;
        RECT 1896.280 510.270 1897.090 510.410 ;
        RECT 1896.280 483.325 1896.420 510.270 ;
        RECT 1896.810 510.000 1897.090 510.270 ;
        RECT 1896.210 482.955 1896.490 483.325 ;
        RECT 1897.130 482.955 1897.410 483.325 ;
        RECT 1897.200 448.790 1897.340 482.955 ;
        RECT 1896.220 448.530 1896.480 448.790 ;
        RECT 1896.220 448.470 1896.880 448.530 ;
        RECT 1897.140 448.470 1897.400 448.790 ;
        RECT 1896.280 448.390 1896.880 448.470 ;
        RECT 1896.740 400.850 1896.880 448.390 ;
        RECT 1896.680 400.530 1896.940 400.850 ;
        RECT 1896.680 399.850 1896.940 400.170 ;
        RECT 1896.740 351.970 1896.880 399.850 ;
        RECT 1896.280 351.830 1896.880 351.970 ;
        RECT 1896.280 351.290 1896.420 351.830 ;
        RECT 1896.280 351.150 1896.880 351.290 ;
        RECT 1896.740 255.410 1896.880 351.150 ;
        RECT 1896.280 255.270 1896.880 255.410 ;
        RECT 1896.280 237.990 1896.420 255.270 ;
        RECT 1896.220 237.670 1896.480 237.990 ;
        RECT 2070.100 237.670 2070.360 237.990 ;
        RECT 2070.160 62.210 2070.300 237.670 ;
        RECT 2070.100 61.890 2070.360 62.210 ;
        RECT 2072.400 61.890 2072.660 62.210 ;
        RECT 2072.460 48.270 2072.600 61.890 ;
        RECT 2072.400 47.950 2072.660 48.270 ;
        RECT 2072.400 2.730 2072.660 3.050 ;
        RECT 2072.460 2.400 2072.600 2.730 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 1896.210 483.000 1896.490 483.280 ;
        RECT 1897.130 483.000 1897.410 483.280 ;
      LAYER met3 ;
        RECT 1896.185 483.290 1896.515 483.305 ;
        RECT 1897.105 483.290 1897.435 483.305 ;
        RECT 1896.185 482.990 1897.435 483.290 ;
        RECT 1896.185 482.975 1896.515 482.990 ;
        RECT 1897.105 482.975 1897.435 482.990 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.450 245.040 1910.770 245.100 ;
        RECT 2083.870 245.040 2084.190 245.100 ;
        RECT 1910.450 244.900 2084.190 245.040 ;
        RECT 1910.450 244.840 1910.770 244.900 ;
        RECT 2083.870 244.840 2084.190 244.900 ;
        RECT 2083.870 37.980 2084.190 38.040 ;
        RECT 2089.850 37.980 2090.170 38.040 ;
        RECT 2083.870 37.840 2090.170 37.980 ;
        RECT 2083.870 37.780 2084.190 37.840 ;
        RECT 2089.850 37.780 2090.170 37.840 ;
      LAYER via ;
        RECT 1910.480 244.840 1910.740 245.100 ;
        RECT 2083.900 244.840 2084.160 245.100 ;
        RECT 2083.900 37.780 2084.160 38.040 ;
        RECT 2089.880 37.780 2090.140 38.040 ;
      LAYER met2 ;
        RECT 1909.690 510.410 1909.970 514.000 ;
        RECT 1909.690 510.270 1910.680 510.410 ;
        RECT 1909.690 510.000 1909.970 510.270 ;
        RECT 1910.540 245.130 1910.680 510.270 ;
        RECT 1910.480 244.810 1910.740 245.130 ;
        RECT 2083.900 244.810 2084.160 245.130 ;
        RECT 2083.960 38.070 2084.100 244.810 ;
        RECT 2083.900 37.750 2084.160 38.070 ;
        RECT 2089.880 37.750 2090.140 38.070 ;
        RECT 2089.940 2.400 2090.080 37.750 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.250 258.640 1924.570 258.700 ;
        RECT 2104.570 258.640 2104.890 258.700 ;
        RECT 1924.250 258.500 2104.890 258.640 ;
        RECT 1924.250 258.440 1924.570 258.500 ;
        RECT 2104.570 258.440 2104.890 258.500 ;
        RECT 2104.570 62.120 2104.890 62.180 ;
        RECT 2107.790 62.120 2108.110 62.180 ;
        RECT 2104.570 61.980 2108.110 62.120 ;
        RECT 2104.570 61.920 2104.890 61.980 ;
        RECT 2107.790 61.920 2108.110 61.980 ;
      LAYER via ;
        RECT 1924.280 258.440 1924.540 258.700 ;
        RECT 2104.600 258.440 2104.860 258.700 ;
        RECT 2104.600 61.920 2104.860 62.180 ;
        RECT 2107.820 61.920 2108.080 62.180 ;
      LAYER met2 ;
        RECT 1922.570 510.410 1922.850 514.000 ;
        RECT 1922.570 510.270 1924.480 510.410 ;
        RECT 1922.570 510.000 1922.850 510.270 ;
        RECT 1924.340 258.730 1924.480 510.270 ;
        RECT 1924.280 258.410 1924.540 258.730 ;
        RECT 2104.600 258.410 2104.860 258.730 ;
        RECT 2104.660 62.210 2104.800 258.410 ;
        RECT 2104.600 61.890 2104.860 62.210 ;
        RECT 2107.820 61.890 2108.080 62.210 ;
        RECT 2107.880 2.400 2108.020 61.890 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 24.040 1938.830 24.100 ;
        RECT 2125.730 24.040 2126.050 24.100 ;
        RECT 1938.510 23.900 2126.050 24.040 ;
        RECT 1938.510 23.840 1938.830 23.900 ;
        RECT 2125.730 23.840 2126.050 23.900 ;
      LAYER via ;
        RECT 1938.540 23.840 1938.800 24.100 ;
        RECT 2125.760 23.840 2126.020 24.100 ;
      LAYER met2 ;
        RECT 1935.450 510.410 1935.730 514.000 ;
        RECT 1935.450 510.270 1938.740 510.410 ;
        RECT 1935.450 510.000 1935.730 510.270 ;
        RECT 1938.600 24.130 1938.740 510.270 ;
        RECT 1938.540 23.810 1938.800 24.130 ;
        RECT 2125.760 23.810 2126.020 24.130 ;
        RECT 2125.820 2.400 2125.960 23.810 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1951.005 193.205 1951.175 241.315 ;
      LAYER mcon ;
        RECT 1951.005 241.145 1951.175 241.315 ;
      LAYER met1 ;
        RECT 1948.170 496.980 1948.490 497.040 ;
        RECT 1948.170 496.840 1952.080 496.980 ;
        RECT 1948.170 496.780 1948.490 496.840 ;
        RECT 1951.940 496.300 1952.080 496.840 ;
        RECT 1952.310 496.300 1952.630 496.360 ;
        RECT 1951.940 496.160 1952.630 496.300 ;
        RECT 1952.310 496.100 1952.630 496.160 ;
        RECT 1950.930 410.620 1951.250 410.680 ;
        RECT 1951.850 410.620 1952.170 410.680 ;
        RECT 1950.930 410.480 1952.170 410.620 ;
        RECT 1950.930 410.420 1951.250 410.480 ;
        RECT 1951.850 410.420 1952.170 410.480 ;
        RECT 1950.010 310.660 1950.330 310.720 ;
        RECT 1950.470 310.660 1950.790 310.720 ;
        RECT 1950.010 310.520 1950.790 310.660 ;
        RECT 1950.010 310.460 1950.330 310.520 ;
        RECT 1950.470 310.460 1950.790 310.520 ;
        RECT 1950.930 262.380 1951.250 262.440 ;
        RECT 1951.390 262.380 1951.710 262.440 ;
        RECT 1950.930 262.240 1951.710 262.380 ;
        RECT 1950.930 262.180 1951.250 262.240 ;
        RECT 1951.390 262.180 1951.710 262.240 ;
        RECT 1950.945 241.300 1951.235 241.345 ;
        RECT 1951.390 241.300 1951.710 241.360 ;
        RECT 1950.945 241.160 1951.710 241.300 ;
        RECT 1950.945 241.115 1951.235 241.160 ;
        RECT 1951.390 241.100 1951.710 241.160 ;
        RECT 1950.930 193.360 1951.250 193.420 ;
        RECT 1950.735 193.220 1951.250 193.360 ;
        RECT 1950.930 193.160 1951.250 193.220 ;
        RECT 1950.930 162.080 1951.250 162.140 ;
        RECT 2139.070 162.080 2139.390 162.140 ;
        RECT 1950.930 161.940 2139.390 162.080 ;
        RECT 1950.930 161.880 1951.250 161.940 ;
        RECT 2139.070 161.880 2139.390 161.940 ;
        RECT 2139.070 62.120 2139.390 62.180 ;
        RECT 2143.670 62.120 2143.990 62.180 ;
        RECT 2139.070 61.980 2143.990 62.120 ;
        RECT 2139.070 61.920 2139.390 61.980 ;
        RECT 2143.670 61.920 2143.990 61.980 ;
      LAYER via ;
        RECT 1948.200 496.780 1948.460 497.040 ;
        RECT 1952.340 496.100 1952.600 496.360 ;
        RECT 1950.960 410.420 1951.220 410.680 ;
        RECT 1951.880 410.420 1952.140 410.680 ;
        RECT 1950.040 310.460 1950.300 310.720 ;
        RECT 1950.500 310.460 1950.760 310.720 ;
        RECT 1950.960 262.180 1951.220 262.440 ;
        RECT 1951.420 262.180 1951.680 262.440 ;
        RECT 1951.420 241.100 1951.680 241.360 ;
        RECT 1950.960 193.160 1951.220 193.420 ;
        RECT 1950.960 161.880 1951.220 162.140 ;
        RECT 2139.100 161.880 2139.360 162.140 ;
        RECT 2139.100 61.920 2139.360 62.180 ;
        RECT 2143.700 61.920 2143.960 62.180 ;
      LAYER met2 ;
        RECT 1948.330 510.340 1948.610 514.000 ;
        RECT 1948.260 510.000 1948.610 510.340 ;
        RECT 1948.260 497.070 1948.400 510.000 ;
        RECT 1948.200 496.750 1948.460 497.070 ;
        RECT 1952.340 496.070 1952.600 496.390 ;
        RECT 1952.400 468.930 1952.540 496.070 ;
        RECT 1951.940 468.790 1952.540 468.930 ;
        RECT 1951.940 448.530 1952.080 468.790 ;
        RECT 1951.020 448.390 1952.080 448.530 ;
        RECT 1951.020 410.710 1951.160 448.390 ;
        RECT 1950.960 410.390 1951.220 410.710 ;
        RECT 1951.880 410.390 1952.140 410.710 ;
        RECT 1951.940 386.765 1952.080 410.390 ;
        RECT 1950.950 386.650 1951.230 386.765 ;
        RECT 1950.560 386.510 1951.230 386.650 ;
        RECT 1950.560 310.750 1950.700 386.510 ;
        RECT 1950.950 386.395 1951.230 386.510 ;
        RECT 1951.870 386.395 1952.150 386.765 ;
        RECT 1950.040 310.430 1950.300 310.750 ;
        RECT 1950.500 310.430 1950.760 310.750 ;
        RECT 1950.100 304.370 1950.240 310.430 ;
        RECT 1950.100 304.230 1951.160 304.370 ;
        RECT 1951.020 262.470 1951.160 304.230 ;
        RECT 1950.960 262.150 1951.220 262.470 ;
        RECT 1951.420 262.150 1951.680 262.470 ;
        RECT 1951.480 241.390 1951.620 262.150 ;
        RECT 1951.420 241.070 1951.680 241.390 ;
        RECT 1950.960 193.130 1951.220 193.450 ;
        RECT 1951.020 162.170 1951.160 193.130 ;
        RECT 1950.960 161.850 1951.220 162.170 ;
        RECT 2139.100 161.850 2139.360 162.170 ;
        RECT 2139.160 62.210 2139.300 161.850 ;
        RECT 2139.100 61.890 2139.360 62.210 ;
        RECT 2143.700 61.890 2143.960 62.210 ;
        RECT 2143.760 2.400 2143.900 61.890 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
      LAYER via2 ;
        RECT 1950.950 386.440 1951.230 386.720 ;
        RECT 1951.870 386.440 1952.150 386.720 ;
      LAYER met3 ;
        RECT 1950.925 386.730 1951.255 386.745 ;
        RECT 1951.845 386.730 1952.175 386.745 ;
        RECT 1950.925 386.430 1952.175 386.730 ;
        RECT 1950.925 386.415 1951.255 386.430 ;
        RECT 1951.845 386.415 1952.175 386.430 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2139.145 282.965 2139.315 286.195 ;
        RECT 2159.845 186.405 2160.015 234.515 ;
        RECT 2159.845 89.845 2160.015 137.955 ;
        RECT 2161.685 2.805 2161.855 48.195 ;
      LAYER mcon ;
        RECT 2139.145 286.025 2139.315 286.195 ;
        RECT 2159.845 234.345 2160.015 234.515 ;
        RECT 2159.845 137.785 2160.015 137.955 ;
        RECT 2161.685 48.025 2161.855 48.195 ;
      LAYER met1 ;
        RECT 1961.050 496.980 1961.370 497.040 ;
        RECT 1965.650 496.980 1965.970 497.040 ;
        RECT 1961.050 496.840 1965.970 496.980 ;
        RECT 1961.050 496.780 1961.370 496.840 ;
        RECT 1965.650 496.780 1965.970 496.840 ;
        RECT 1965.650 286.180 1965.970 286.240 ;
        RECT 2139.085 286.180 2139.375 286.225 ;
        RECT 1965.650 286.040 2139.375 286.180 ;
        RECT 1965.650 285.980 1965.970 286.040 ;
        RECT 2139.085 285.995 2139.375 286.040 ;
        RECT 2139.085 283.120 2139.375 283.165 ;
        RECT 2159.770 283.120 2160.090 283.180 ;
        RECT 2139.085 282.980 2160.090 283.120 ;
        RECT 2139.085 282.935 2139.375 282.980 ;
        RECT 2159.770 282.920 2160.090 282.980 ;
        RECT 2159.770 234.500 2160.090 234.560 ;
        RECT 2159.575 234.360 2160.090 234.500 ;
        RECT 2159.770 234.300 2160.090 234.360 ;
        RECT 2159.770 186.560 2160.090 186.620 ;
        RECT 2159.575 186.420 2160.090 186.560 ;
        RECT 2159.770 186.360 2160.090 186.420 ;
        RECT 2159.770 137.940 2160.090 138.000 ;
        RECT 2159.575 137.800 2160.090 137.940 ;
        RECT 2159.770 137.740 2160.090 137.800 ;
        RECT 2159.770 90.000 2160.090 90.060 ;
        RECT 2159.575 89.860 2160.090 90.000 ;
        RECT 2159.770 89.800 2160.090 89.860 ;
        RECT 2161.610 48.180 2161.930 48.240 ;
        RECT 2161.415 48.040 2161.930 48.180 ;
        RECT 2161.610 47.980 2161.930 48.040 ;
        RECT 2161.610 2.960 2161.930 3.020 ;
        RECT 2161.415 2.820 2161.930 2.960 ;
        RECT 2161.610 2.760 2161.930 2.820 ;
      LAYER via ;
        RECT 1961.080 496.780 1961.340 497.040 ;
        RECT 1965.680 496.780 1965.940 497.040 ;
        RECT 1965.680 285.980 1965.940 286.240 ;
        RECT 2159.800 282.920 2160.060 283.180 ;
        RECT 2159.800 234.300 2160.060 234.560 ;
        RECT 2159.800 186.360 2160.060 186.620 ;
        RECT 2159.800 137.740 2160.060 138.000 ;
        RECT 2159.800 89.800 2160.060 90.060 ;
        RECT 2161.640 47.980 2161.900 48.240 ;
        RECT 2161.640 2.760 2161.900 3.020 ;
      LAYER met2 ;
        RECT 1961.210 510.340 1961.490 514.000 ;
        RECT 1961.140 510.000 1961.490 510.340 ;
        RECT 1961.140 497.070 1961.280 510.000 ;
        RECT 1961.080 496.750 1961.340 497.070 ;
        RECT 1965.680 496.750 1965.940 497.070 ;
        RECT 1965.740 286.270 1965.880 496.750 ;
        RECT 1965.680 285.950 1965.940 286.270 ;
        RECT 2159.800 282.890 2160.060 283.210 ;
        RECT 2159.860 234.590 2160.000 282.890 ;
        RECT 2159.800 234.270 2160.060 234.590 ;
        RECT 2159.800 186.330 2160.060 186.650 ;
        RECT 2159.860 138.030 2160.000 186.330 ;
        RECT 2159.800 137.710 2160.060 138.030 ;
        RECT 2159.800 89.770 2160.060 90.090 ;
        RECT 2159.860 74.530 2160.000 89.770 ;
        RECT 2159.860 74.390 2160.460 74.530 ;
        RECT 2160.320 61.610 2160.460 74.390 ;
        RECT 2160.320 61.470 2161.840 61.610 ;
        RECT 2161.700 48.270 2161.840 61.470 ;
        RECT 2161.640 47.950 2161.900 48.270 ;
        RECT 2161.640 2.730 2161.900 3.050 ;
        RECT 2161.700 2.400 2161.840 2.730 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.470 496.980 1973.790 497.040 ;
        RECT 1979.450 496.980 1979.770 497.040 ;
        RECT 1973.470 496.840 1979.770 496.980 ;
        RECT 1973.470 496.780 1973.790 496.840 ;
        RECT 1979.450 496.780 1979.770 496.840 ;
        RECT 1979.450 293.320 1979.770 293.380 ;
        RECT 2173.570 293.320 2173.890 293.380 ;
        RECT 1979.450 293.180 2173.890 293.320 ;
        RECT 1979.450 293.120 1979.770 293.180 ;
        RECT 2173.570 293.120 2173.890 293.180 ;
        RECT 2173.570 62.120 2173.890 62.180 ;
        RECT 2179.090 62.120 2179.410 62.180 ;
        RECT 2173.570 61.980 2179.410 62.120 ;
        RECT 2173.570 61.920 2173.890 61.980 ;
        RECT 2179.090 61.920 2179.410 61.980 ;
      LAYER via ;
        RECT 1973.500 496.780 1973.760 497.040 ;
        RECT 1979.480 496.780 1979.740 497.040 ;
        RECT 1979.480 293.120 1979.740 293.380 ;
        RECT 2173.600 293.120 2173.860 293.380 ;
        RECT 2173.600 61.920 2173.860 62.180 ;
        RECT 2179.120 61.920 2179.380 62.180 ;
      LAYER met2 ;
        RECT 1973.630 510.340 1973.910 514.000 ;
        RECT 1973.560 510.000 1973.910 510.340 ;
        RECT 1973.560 497.070 1973.700 510.000 ;
        RECT 1973.500 496.750 1973.760 497.070 ;
        RECT 1979.480 496.750 1979.740 497.070 ;
        RECT 1979.540 293.410 1979.680 496.750 ;
        RECT 1979.480 293.090 1979.740 293.410 ;
        RECT 2173.600 293.090 2173.860 293.410 ;
        RECT 2173.660 62.210 2173.800 293.090 ;
        RECT 2173.600 61.890 2173.860 62.210 ;
        RECT 2179.120 61.890 2179.380 62.210 ;
        RECT 2179.180 2.400 2179.320 61.890 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.350 497.320 1986.670 497.380 ;
        RECT 1997.390 497.320 1997.710 497.380 ;
        RECT 1986.350 497.180 1997.710 497.320 ;
        RECT 1986.350 497.120 1986.670 497.180 ;
        RECT 1997.390 497.120 1997.710 497.180 ;
        RECT 1997.390 182.820 1997.710 182.880 ;
        RECT 2194.270 182.820 2194.590 182.880 ;
        RECT 1997.390 182.680 2194.590 182.820 ;
        RECT 1997.390 182.620 1997.710 182.680 ;
        RECT 2194.270 182.620 2194.590 182.680 ;
      LAYER via ;
        RECT 1986.380 497.120 1986.640 497.380 ;
        RECT 1997.420 497.120 1997.680 497.380 ;
        RECT 1997.420 182.620 1997.680 182.880 ;
        RECT 2194.300 182.620 2194.560 182.880 ;
      LAYER met2 ;
        RECT 1986.510 510.340 1986.790 514.000 ;
        RECT 1986.440 510.000 1986.790 510.340 ;
        RECT 1986.440 497.410 1986.580 510.000 ;
        RECT 1986.380 497.090 1986.640 497.410 ;
        RECT 1997.420 497.090 1997.680 497.410 ;
        RECT 1997.480 182.910 1997.620 497.090 ;
        RECT 1997.420 182.590 1997.680 182.910 ;
        RECT 2194.300 182.590 2194.560 182.910 ;
        RECT 2194.360 17.410 2194.500 182.590 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1999.230 493.580 1999.550 493.640 ;
        RECT 2214.970 493.580 2215.290 493.640 ;
        RECT 1999.230 493.440 2215.290 493.580 ;
        RECT 1999.230 493.380 1999.550 493.440 ;
        RECT 2214.970 493.380 2215.290 493.440 ;
      LAYER via ;
        RECT 1999.260 493.380 1999.520 493.640 ;
        RECT 2215.000 493.380 2215.260 493.640 ;
      LAYER met2 ;
        RECT 1999.390 510.340 1999.670 514.000 ;
        RECT 1999.320 510.000 1999.670 510.340 ;
        RECT 1999.320 493.670 1999.460 510.000 ;
        RECT 1999.260 493.350 1999.520 493.670 ;
        RECT 2215.000 493.350 2215.260 493.670 ;
        RECT 2215.060 2.400 2215.200 493.350 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2014.410 20.640 2014.730 20.700 ;
        RECT 2232.910 20.640 2233.230 20.700 ;
        RECT 2014.410 20.500 2233.230 20.640 ;
        RECT 2014.410 20.440 2014.730 20.500 ;
        RECT 2232.910 20.440 2233.230 20.500 ;
      LAYER via ;
        RECT 2014.440 20.440 2014.700 20.700 ;
        RECT 2232.940 20.440 2233.200 20.700 ;
      LAYER met2 ;
        RECT 2012.270 510.410 2012.550 514.000 ;
        RECT 2012.270 510.270 2014.640 510.410 ;
        RECT 2012.270 510.000 2012.550 510.270 ;
        RECT 2014.500 20.730 2014.640 510.270 ;
        RECT 2014.440 20.410 2014.700 20.730 ;
        RECT 2232.940 20.410 2233.200 20.730 ;
        RECT 2233.000 2.400 2233.140 20.410 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 237.900 793.430 237.960 ;
        RECT 973.430 237.900 973.750 237.960 ;
        RECT 793.110 237.760 973.750 237.900 ;
        RECT 793.110 237.700 793.430 237.760 ;
        RECT 973.430 237.700 973.750 237.760 ;
        RECT 787.590 19.280 787.910 19.340 ;
        RECT 793.110 19.280 793.430 19.340 ;
        RECT 787.590 19.140 793.430 19.280 ;
        RECT 787.590 19.080 787.910 19.140 ;
        RECT 793.110 19.080 793.430 19.140 ;
      LAYER via ;
        RECT 793.140 237.700 793.400 237.960 ;
        RECT 973.460 237.700 973.720 237.960 ;
        RECT 787.620 19.080 787.880 19.340 ;
        RECT 793.140 19.080 793.400 19.340 ;
      LAYER met2 ;
        RECT 974.970 510.410 975.250 514.000 ;
        RECT 973.520 510.270 975.250 510.410 ;
        RECT 973.520 237.990 973.660 510.270 ;
        RECT 974.970 510.000 975.250 510.270 ;
        RECT 793.140 237.670 793.400 237.990 ;
        RECT 973.460 237.670 973.720 237.990 ;
        RECT 793.200 19.370 793.340 237.670 ;
        RECT 787.620 19.050 787.880 19.370 ;
        RECT 793.140 19.050 793.400 19.370 ;
        RECT 787.680 2.400 787.820 19.050 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.210 19.960 2028.530 20.020 ;
        RECT 2250.850 19.960 2251.170 20.020 ;
        RECT 2028.210 19.820 2251.170 19.960 ;
        RECT 2028.210 19.760 2028.530 19.820 ;
        RECT 2250.850 19.760 2251.170 19.820 ;
      LAYER via ;
        RECT 2028.240 19.760 2028.500 20.020 ;
        RECT 2250.880 19.760 2251.140 20.020 ;
      LAYER met2 ;
        RECT 2025.150 510.410 2025.430 514.000 ;
        RECT 2025.150 510.270 2028.440 510.410 ;
        RECT 2025.150 510.000 2025.430 510.270 ;
        RECT 2028.300 20.050 2028.440 510.270 ;
        RECT 2028.240 19.730 2028.500 20.050 ;
        RECT 2250.880 19.730 2251.140 20.050 ;
        RECT 2250.940 2.400 2251.080 19.730 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2041.165 427.805 2041.335 475.575 ;
        RECT 2040.705 331.245 2040.875 379.355 ;
        RECT 2041.165 89.845 2041.335 137.955 ;
        RECT 2042.085 48.365 2042.255 84.235 ;
      LAYER mcon ;
        RECT 2041.165 475.405 2041.335 475.575 ;
        RECT 2040.705 379.185 2040.875 379.355 ;
        RECT 2041.165 137.785 2041.335 137.955 ;
        RECT 2042.085 84.065 2042.255 84.235 ;
      LAYER met1 ;
        RECT 2037.870 476.240 2038.190 476.300 ;
        RECT 2041.090 476.240 2041.410 476.300 ;
        RECT 2037.870 476.100 2041.410 476.240 ;
        RECT 2037.870 476.040 2038.190 476.100 ;
        RECT 2041.090 476.040 2041.410 476.100 ;
        RECT 2041.090 475.560 2041.410 475.620 ;
        RECT 2040.895 475.420 2041.410 475.560 ;
        RECT 2041.090 475.360 2041.410 475.420 ;
        RECT 2041.090 427.960 2041.410 428.020 ;
        RECT 2040.895 427.820 2041.410 427.960 ;
        RECT 2041.090 427.760 2041.410 427.820 ;
        RECT 2040.630 380.020 2040.950 380.080 ;
        RECT 2041.090 380.020 2041.410 380.080 ;
        RECT 2040.630 379.880 2041.410 380.020 ;
        RECT 2040.630 379.820 2040.950 379.880 ;
        RECT 2041.090 379.820 2041.410 379.880 ;
        RECT 2040.630 379.340 2040.950 379.400 ;
        RECT 2040.435 379.200 2040.950 379.340 ;
        RECT 2040.630 379.140 2040.950 379.200 ;
        RECT 2040.645 331.400 2040.935 331.445 ;
        RECT 2041.090 331.400 2041.410 331.460 ;
        RECT 2040.645 331.260 2041.410 331.400 ;
        RECT 2040.645 331.215 2040.935 331.260 ;
        RECT 2041.090 331.200 2041.410 331.260 ;
        RECT 2040.630 228.040 2040.950 228.100 ;
        RECT 2041.550 228.040 2041.870 228.100 ;
        RECT 2040.630 227.900 2041.870 228.040 ;
        RECT 2040.630 227.840 2040.950 227.900 ;
        RECT 2041.550 227.840 2041.870 227.900 ;
        RECT 2041.090 137.940 2041.410 138.000 ;
        RECT 2040.895 137.800 2041.410 137.940 ;
        RECT 2041.090 137.740 2041.410 137.800 ;
        RECT 2041.105 90.000 2041.395 90.045 ;
        RECT 2042.010 90.000 2042.330 90.060 ;
        RECT 2041.105 89.860 2042.330 90.000 ;
        RECT 2041.105 89.815 2041.395 89.860 ;
        RECT 2042.010 89.800 2042.330 89.860 ;
        RECT 2042.010 84.220 2042.330 84.280 ;
        RECT 2041.815 84.080 2042.330 84.220 ;
        RECT 2042.010 84.020 2042.330 84.080 ;
        RECT 2042.010 48.520 2042.330 48.580 ;
        RECT 2041.815 48.380 2042.330 48.520 ;
        RECT 2042.010 48.320 2042.330 48.380 ;
        RECT 2042.010 20.300 2042.330 20.360 ;
        RECT 2268.330 20.300 2268.650 20.360 ;
        RECT 2042.010 20.160 2268.650 20.300 ;
        RECT 2042.010 20.100 2042.330 20.160 ;
        RECT 2268.330 20.100 2268.650 20.160 ;
      LAYER via ;
        RECT 2037.900 476.040 2038.160 476.300 ;
        RECT 2041.120 476.040 2041.380 476.300 ;
        RECT 2041.120 475.360 2041.380 475.620 ;
        RECT 2041.120 427.760 2041.380 428.020 ;
        RECT 2040.660 379.820 2040.920 380.080 ;
        RECT 2041.120 379.820 2041.380 380.080 ;
        RECT 2040.660 379.140 2040.920 379.400 ;
        RECT 2041.120 331.200 2041.380 331.460 ;
        RECT 2040.660 227.840 2040.920 228.100 ;
        RECT 2041.580 227.840 2041.840 228.100 ;
        RECT 2041.120 137.740 2041.380 138.000 ;
        RECT 2042.040 89.800 2042.300 90.060 ;
        RECT 2042.040 84.020 2042.300 84.280 ;
        RECT 2042.040 48.320 2042.300 48.580 ;
        RECT 2042.040 20.100 2042.300 20.360 ;
        RECT 2268.360 20.100 2268.620 20.360 ;
      LAYER met2 ;
        RECT 2038.030 510.340 2038.310 514.000 ;
        RECT 2037.960 510.000 2038.310 510.340 ;
        RECT 2037.960 476.330 2038.100 510.000 ;
        RECT 2037.900 476.010 2038.160 476.330 ;
        RECT 2041.120 476.010 2041.380 476.330 ;
        RECT 2041.180 475.650 2041.320 476.010 ;
        RECT 2041.120 475.330 2041.380 475.650 ;
        RECT 2041.120 427.730 2041.380 428.050 ;
        RECT 2041.180 380.110 2041.320 427.730 ;
        RECT 2040.660 379.790 2040.920 380.110 ;
        RECT 2041.120 379.790 2041.380 380.110 ;
        RECT 2040.720 379.430 2040.860 379.790 ;
        RECT 2040.660 379.110 2040.920 379.430 ;
        RECT 2041.120 331.170 2041.380 331.490 ;
        RECT 2041.180 303.690 2041.320 331.170 ;
        RECT 2041.180 303.550 2041.780 303.690 ;
        RECT 2041.640 228.130 2041.780 303.550 ;
        RECT 2040.660 227.810 2040.920 228.130 ;
        RECT 2041.580 227.810 2041.840 228.130 ;
        RECT 2040.720 161.570 2040.860 227.810 ;
        RECT 2040.720 161.430 2041.320 161.570 ;
        RECT 2041.180 138.030 2041.320 161.430 ;
        RECT 2041.120 137.710 2041.380 138.030 ;
        RECT 2042.040 89.770 2042.300 90.090 ;
        RECT 2042.100 84.310 2042.240 89.770 ;
        RECT 2042.040 83.990 2042.300 84.310 ;
        RECT 2042.040 48.290 2042.300 48.610 ;
        RECT 2042.100 20.390 2042.240 48.290 ;
        RECT 2042.040 20.070 2042.300 20.390 ;
        RECT 2268.360 20.070 2268.620 20.390 ;
        RECT 2268.420 2.400 2268.560 20.070 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2050.290 496.980 2050.610 497.040 ;
        RECT 2055.810 496.980 2056.130 497.040 ;
        RECT 2050.290 496.840 2056.130 496.980 ;
        RECT 2050.290 496.780 2050.610 496.840 ;
        RECT 2055.810 496.780 2056.130 496.840 ;
        RECT 2055.810 19.620 2056.130 19.680 ;
        RECT 2286.270 19.620 2286.590 19.680 ;
        RECT 2055.810 19.480 2286.590 19.620 ;
        RECT 2055.810 19.420 2056.130 19.480 ;
        RECT 2286.270 19.420 2286.590 19.480 ;
      LAYER via ;
        RECT 2050.320 496.780 2050.580 497.040 ;
        RECT 2055.840 496.780 2056.100 497.040 ;
        RECT 2055.840 19.420 2056.100 19.680 ;
        RECT 2286.300 19.420 2286.560 19.680 ;
      LAYER met2 ;
        RECT 2050.450 510.340 2050.730 514.000 ;
        RECT 2050.380 510.000 2050.730 510.340 ;
        RECT 2050.380 497.070 2050.520 510.000 ;
        RECT 2050.320 496.750 2050.580 497.070 ;
        RECT 2055.840 496.750 2056.100 497.070 ;
        RECT 2055.900 19.710 2056.040 496.750 ;
        RECT 2055.840 19.390 2056.100 19.710 ;
        RECT 2286.300 19.390 2286.560 19.710 ;
        RECT 2286.360 2.400 2286.500 19.390 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2063.170 496.980 2063.490 497.040 ;
        RECT 2069.610 496.980 2069.930 497.040 ;
        RECT 2063.170 496.840 2069.930 496.980 ;
        RECT 2063.170 496.780 2063.490 496.840 ;
        RECT 2069.610 496.780 2069.930 496.840 ;
        RECT 2069.610 19.280 2069.930 19.340 ;
        RECT 2304.210 19.280 2304.530 19.340 ;
        RECT 2069.610 19.140 2304.530 19.280 ;
        RECT 2069.610 19.080 2069.930 19.140 ;
        RECT 2304.210 19.080 2304.530 19.140 ;
      LAYER via ;
        RECT 2063.200 496.780 2063.460 497.040 ;
        RECT 2069.640 496.780 2069.900 497.040 ;
        RECT 2069.640 19.080 2069.900 19.340 ;
        RECT 2304.240 19.080 2304.500 19.340 ;
      LAYER met2 ;
        RECT 2063.330 510.340 2063.610 514.000 ;
        RECT 2063.260 510.000 2063.610 510.340 ;
        RECT 2063.260 497.070 2063.400 510.000 ;
        RECT 2063.200 496.750 2063.460 497.070 ;
        RECT 2069.640 496.750 2069.900 497.070 ;
        RECT 2069.700 19.370 2069.840 496.750 ;
        RECT 2069.640 19.050 2069.900 19.370 ;
        RECT 2304.240 19.050 2304.500 19.370 ;
        RECT 2304.300 2.400 2304.440 19.050 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2075.205 414.205 2075.375 462.315 ;
        RECT 2076.585 179.605 2076.755 244.715 ;
      LAYER mcon ;
        RECT 2075.205 462.145 2075.375 462.315 ;
        RECT 2076.585 244.545 2076.755 244.715 ;
      LAYER met1 ;
        RECT 2075.130 462.300 2075.450 462.360 ;
        RECT 2074.935 462.160 2075.450 462.300 ;
        RECT 2075.130 462.100 2075.450 462.160 ;
        RECT 2075.130 414.360 2075.450 414.420 ;
        RECT 2074.935 414.220 2075.450 414.360 ;
        RECT 2075.130 414.160 2075.450 414.220 ;
        RECT 2075.130 400.220 2075.450 400.480 ;
        RECT 2075.220 399.740 2075.360 400.220 ;
        RECT 2075.590 399.740 2075.910 399.800 ;
        RECT 2075.220 399.600 2075.910 399.740 ;
        RECT 2075.590 399.540 2075.910 399.600 ;
        RECT 2075.590 365.740 2075.910 365.800 ;
        RECT 2076.970 365.740 2077.290 365.800 ;
        RECT 2075.590 365.600 2077.290 365.740 ;
        RECT 2075.590 365.540 2075.910 365.600 ;
        RECT 2076.970 365.540 2077.290 365.600 ;
        RECT 2076.525 244.700 2076.815 244.745 ;
        RECT 2076.970 244.700 2077.290 244.760 ;
        RECT 2076.525 244.560 2077.290 244.700 ;
        RECT 2076.525 244.515 2076.815 244.560 ;
        RECT 2076.970 244.500 2077.290 244.560 ;
        RECT 2076.510 179.760 2076.830 179.820 ;
        RECT 2076.315 179.620 2076.830 179.760 ;
        RECT 2076.510 179.560 2076.830 179.620 ;
        RECT 2075.590 18.940 2075.910 19.000 ;
        RECT 2322.150 18.940 2322.470 19.000 ;
        RECT 2075.590 18.800 2322.470 18.940 ;
        RECT 2075.590 18.740 2075.910 18.800 ;
        RECT 2322.150 18.740 2322.470 18.800 ;
      LAYER via ;
        RECT 2075.160 462.100 2075.420 462.360 ;
        RECT 2075.160 414.160 2075.420 414.420 ;
        RECT 2075.160 400.220 2075.420 400.480 ;
        RECT 2075.620 399.540 2075.880 399.800 ;
        RECT 2075.620 365.540 2075.880 365.800 ;
        RECT 2077.000 365.540 2077.260 365.800 ;
        RECT 2077.000 244.500 2077.260 244.760 ;
        RECT 2076.540 179.560 2076.800 179.820 ;
        RECT 2075.620 18.740 2075.880 19.000 ;
        RECT 2322.180 18.740 2322.440 19.000 ;
      LAYER met2 ;
        RECT 2076.210 510.410 2076.490 514.000 ;
        RECT 2075.220 510.270 2076.490 510.410 ;
        RECT 2075.220 462.390 2075.360 510.270 ;
        RECT 2076.210 510.000 2076.490 510.270 ;
        RECT 2075.160 462.070 2075.420 462.390 ;
        RECT 2075.160 414.130 2075.420 414.450 ;
        RECT 2075.220 400.510 2075.360 414.130 ;
        RECT 2075.160 400.190 2075.420 400.510 ;
        RECT 2075.620 399.510 2075.880 399.830 ;
        RECT 2075.680 365.830 2075.820 399.510 ;
        RECT 2075.620 365.510 2075.880 365.830 ;
        RECT 2077.000 365.510 2077.260 365.830 ;
        RECT 2077.060 244.790 2077.200 365.510 ;
        RECT 2077.000 244.470 2077.260 244.790 ;
        RECT 2076.540 179.530 2076.800 179.850 ;
        RECT 2076.600 62.970 2076.740 179.530 ;
        RECT 2076.140 62.830 2076.740 62.970 ;
        RECT 2076.140 62.290 2076.280 62.830 ;
        RECT 2075.680 62.150 2076.280 62.290 ;
        RECT 2075.680 19.030 2075.820 62.150 ;
        RECT 2075.620 18.710 2075.880 19.030 ;
        RECT 2322.180 18.710 2322.440 19.030 ;
        RECT 2322.240 2.400 2322.380 18.710 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 18.260 2090.630 18.320 ;
        RECT 2339.170 18.260 2339.490 18.320 ;
        RECT 2090.310 18.120 2339.490 18.260 ;
        RECT 2090.310 18.060 2090.630 18.120 ;
        RECT 2339.170 18.060 2339.490 18.120 ;
      LAYER via ;
        RECT 2090.340 18.060 2090.600 18.320 ;
        RECT 2339.200 18.060 2339.460 18.320 ;
      LAYER met2 ;
        RECT 2089.090 510.410 2089.370 514.000 ;
        RECT 2089.090 510.270 2090.540 510.410 ;
        RECT 2089.090 510.000 2089.370 510.270 ;
        RECT 2090.400 18.350 2090.540 510.270 ;
        RECT 2090.340 18.030 2090.600 18.350 ;
        RECT 2339.200 18.030 2339.460 18.350 ;
        RECT 2339.260 16.050 2339.400 18.030 ;
        RECT 2339.260 15.910 2339.860 16.050 ;
        RECT 2339.720 2.400 2339.860 15.910 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 18.600 2104.430 18.660 ;
        RECT 2357.570 18.600 2357.890 18.660 ;
        RECT 2104.110 18.460 2357.890 18.600 ;
        RECT 2104.110 18.400 2104.430 18.460 ;
        RECT 2357.570 18.400 2357.890 18.460 ;
      LAYER via ;
        RECT 2104.140 18.400 2104.400 18.660 ;
        RECT 2357.600 18.400 2357.860 18.660 ;
      LAYER met2 ;
        RECT 2101.970 510.410 2102.250 514.000 ;
        RECT 2101.970 510.270 2104.340 510.410 ;
        RECT 2101.970 510.000 2102.250 510.270 ;
        RECT 2104.200 18.690 2104.340 510.270 ;
        RECT 2104.140 18.370 2104.400 18.690 ;
        RECT 2357.600 18.370 2357.860 18.690 ;
        RECT 2357.660 2.400 2357.800 18.370 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 17.580 2118.230 17.640 ;
        RECT 2375.510 17.580 2375.830 17.640 ;
        RECT 2117.910 17.440 2375.830 17.580 ;
        RECT 2117.910 17.380 2118.230 17.440 ;
        RECT 2375.510 17.380 2375.830 17.440 ;
      LAYER via ;
        RECT 2117.940 17.380 2118.200 17.640 ;
        RECT 2375.540 17.380 2375.800 17.640 ;
      LAYER met2 ;
        RECT 2114.850 510.410 2115.130 514.000 ;
        RECT 2114.850 510.270 2118.140 510.410 ;
        RECT 2114.850 510.000 2115.130 510.270 ;
        RECT 2118.000 17.670 2118.140 510.270 ;
        RECT 2117.940 17.350 2118.200 17.670 ;
        RECT 2375.540 17.350 2375.800 17.670 ;
        RECT 2375.600 2.400 2375.740 17.350 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2131.325 241.485 2131.495 289.595 ;
      LAYER mcon ;
        RECT 2131.325 289.425 2131.495 289.595 ;
      LAYER met1 ;
        RECT 2127.110 503.440 2127.430 503.500 ;
        RECT 2131.250 503.440 2131.570 503.500 ;
        RECT 2127.110 503.300 2131.570 503.440 ;
        RECT 2127.110 503.240 2127.430 503.300 ;
        RECT 2131.250 503.240 2131.570 503.300 ;
        RECT 2130.330 427.620 2130.650 427.680 ;
        RECT 2130.790 427.620 2131.110 427.680 ;
        RECT 2130.330 427.480 2131.110 427.620 ;
        RECT 2130.330 427.420 2130.650 427.480 ;
        RECT 2130.790 427.420 2131.110 427.480 ;
        RECT 2131.250 289.580 2131.570 289.640 ;
        RECT 2131.055 289.440 2131.570 289.580 ;
        RECT 2131.250 289.380 2131.570 289.440 ;
        RECT 2131.265 241.640 2131.555 241.685 ;
        RECT 2131.710 241.640 2132.030 241.700 ;
        RECT 2131.265 241.500 2132.030 241.640 ;
        RECT 2131.265 241.455 2131.555 241.500 ;
        RECT 2131.710 241.440 2132.030 241.500 ;
        RECT 2130.790 206.960 2131.110 207.020 ;
        RECT 2131.710 206.960 2132.030 207.020 ;
        RECT 2130.790 206.820 2132.030 206.960 ;
        RECT 2130.790 206.760 2131.110 206.820 ;
        RECT 2131.710 206.760 2132.030 206.820 ;
        RECT 2130.330 17.920 2130.650 17.980 ;
        RECT 2393.450 17.920 2393.770 17.980 ;
        RECT 2130.330 17.780 2393.770 17.920 ;
        RECT 2130.330 17.720 2130.650 17.780 ;
        RECT 2393.450 17.720 2393.770 17.780 ;
      LAYER via ;
        RECT 2127.140 503.240 2127.400 503.500 ;
        RECT 2131.280 503.240 2131.540 503.500 ;
        RECT 2130.360 427.420 2130.620 427.680 ;
        RECT 2130.820 427.420 2131.080 427.680 ;
        RECT 2131.280 289.380 2131.540 289.640 ;
        RECT 2131.740 241.440 2132.000 241.700 ;
        RECT 2130.820 206.760 2131.080 207.020 ;
        RECT 2131.740 206.760 2132.000 207.020 ;
        RECT 2130.360 17.720 2130.620 17.980 ;
        RECT 2393.480 17.720 2393.740 17.980 ;
      LAYER met2 ;
        RECT 2127.270 510.340 2127.550 514.000 ;
        RECT 2127.200 510.000 2127.550 510.340 ;
        RECT 2127.200 503.530 2127.340 510.000 ;
        RECT 2127.140 503.210 2127.400 503.530 ;
        RECT 2131.280 503.210 2131.540 503.530 ;
        RECT 2131.340 448.530 2131.480 503.210 ;
        RECT 2130.420 448.390 2131.480 448.530 ;
        RECT 2130.420 427.710 2130.560 448.390 ;
        RECT 2130.360 427.390 2130.620 427.710 ;
        RECT 2130.820 427.390 2131.080 427.710 ;
        RECT 2130.880 351.290 2131.020 427.390 ;
        RECT 2130.420 351.150 2131.020 351.290 ;
        RECT 2130.420 303.690 2130.560 351.150 ;
        RECT 2130.420 303.550 2131.020 303.690 ;
        RECT 2130.880 303.010 2131.020 303.550 ;
        RECT 2130.880 302.870 2131.480 303.010 ;
        RECT 2131.340 289.670 2131.480 302.870 ;
        RECT 2131.280 289.350 2131.540 289.670 ;
        RECT 2131.740 241.410 2132.000 241.730 ;
        RECT 2131.800 207.130 2131.940 241.410 ;
        RECT 2130.880 207.050 2131.940 207.130 ;
        RECT 2130.820 206.990 2132.000 207.050 ;
        RECT 2130.820 206.730 2131.080 206.990 ;
        RECT 2131.740 206.730 2132.000 206.990 ;
        RECT 2131.800 111.250 2131.940 206.730 ;
        RECT 2130.420 111.110 2131.940 111.250 ;
        RECT 2130.420 110.570 2130.560 111.110 ;
        RECT 2129.960 110.430 2130.560 110.570 ;
        RECT 2129.960 90.850 2130.100 110.430 ;
        RECT 2129.960 90.710 2130.560 90.850 ;
        RECT 2130.420 18.010 2130.560 90.710 ;
        RECT 2130.360 17.690 2130.620 18.010 ;
        RECT 2393.480 17.690 2393.740 18.010 ;
        RECT 2393.540 2.400 2393.680 17.690 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2139.990 493.240 2140.310 493.300 ;
        RECT 2145.510 493.240 2145.830 493.300 ;
        RECT 2139.990 493.100 2145.830 493.240 ;
        RECT 2139.990 493.040 2140.310 493.100 ;
        RECT 2145.510 493.040 2145.830 493.100 ;
        RECT 2145.510 17.240 2145.830 17.300 ;
        RECT 2411.390 17.240 2411.710 17.300 ;
        RECT 2145.510 17.100 2411.710 17.240 ;
        RECT 2145.510 17.040 2145.830 17.100 ;
        RECT 2411.390 17.040 2411.710 17.100 ;
      LAYER via ;
        RECT 2140.020 493.040 2140.280 493.300 ;
        RECT 2145.540 493.040 2145.800 493.300 ;
        RECT 2145.540 17.040 2145.800 17.300 ;
        RECT 2411.420 17.040 2411.680 17.300 ;
      LAYER met2 ;
        RECT 2140.150 510.340 2140.430 514.000 ;
        RECT 2140.080 510.000 2140.430 510.340 ;
        RECT 2140.080 493.330 2140.220 510.000 ;
        RECT 2140.020 493.010 2140.280 493.330 ;
        RECT 2145.540 493.010 2145.800 493.330 ;
        RECT 2145.600 17.330 2145.740 493.010 ;
        RECT 2145.540 17.010 2145.800 17.330 ;
        RECT 2411.420 17.010 2411.680 17.330 ;
        RECT 2411.480 2.400 2411.620 17.010 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 286.180 807.230 286.240 ;
        RECT 987.230 286.180 987.550 286.240 ;
        RECT 806.910 286.040 987.550 286.180 ;
        RECT 806.910 285.980 807.230 286.040 ;
        RECT 987.230 285.980 987.550 286.040 ;
        RECT 805.530 2.960 805.850 3.020 ;
        RECT 806.910 2.960 807.230 3.020 ;
        RECT 805.530 2.820 807.230 2.960 ;
        RECT 805.530 2.760 805.850 2.820 ;
        RECT 806.910 2.760 807.230 2.820 ;
      LAYER via ;
        RECT 806.940 285.980 807.200 286.240 ;
        RECT 987.260 285.980 987.520 286.240 ;
        RECT 805.560 2.760 805.820 3.020 ;
        RECT 806.940 2.760 807.200 3.020 ;
      LAYER met2 ;
        RECT 987.850 510.410 988.130 514.000 ;
        RECT 987.320 510.270 988.130 510.410 ;
        RECT 987.320 286.270 987.460 510.270 ;
        RECT 987.850 510.000 988.130 510.270 ;
        RECT 806.940 285.950 807.200 286.270 ;
        RECT 987.260 285.950 987.520 286.270 ;
        RECT 807.000 3.050 807.140 285.950 ;
        RECT 805.560 2.730 805.820 3.050 ;
        RECT 806.940 2.730 807.200 3.050 ;
        RECT 805.620 2.400 805.760 2.730 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 6.970 24.040 7.290 24.100 ;
        RECT 407.170 24.040 407.490 24.100 ;
        RECT 6.970 23.900 407.490 24.040 ;
        RECT 6.970 23.840 7.290 23.900 ;
        RECT 407.170 23.840 407.490 23.900 ;
        RECT 2.830 14.180 3.150 14.240 ;
        RECT 6.970 14.180 7.290 14.240 ;
        RECT 2.830 14.040 7.290 14.180 ;
        RECT 2.830 13.980 3.150 14.040 ;
        RECT 6.970 13.980 7.290 14.040 ;
      LAYER via ;
        RECT 7.000 23.840 7.260 24.100 ;
        RECT 407.200 23.840 407.460 24.100 ;
        RECT 2.860 13.980 3.120 14.240 ;
        RECT 7.000 13.980 7.260 14.240 ;
      LAYER met2 ;
        RECT 411.930 510.410 412.210 514.000 ;
        RECT 407.260 510.270 412.210 510.410 ;
        RECT 407.260 24.130 407.400 510.270 ;
        RECT 411.930 510.000 412.210 510.270 ;
        RECT 7.000 23.810 7.260 24.130 ;
        RECT 407.200 23.810 407.460 24.130 ;
        RECT 7.060 14.270 7.200 23.810 ;
        RECT 2.860 13.950 3.120 14.270 ;
        RECT 7.000 13.950 7.260 14.270 ;
        RECT 2.920 2.400 3.060 13.950 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 500.040 45.010 500.100 ;
        RECT 415.910 500.040 416.230 500.100 ;
        RECT 44.690 499.900 416.230 500.040 ;
        RECT 44.690 499.840 45.010 499.900 ;
        RECT 415.910 499.840 416.230 499.900 ;
        RECT 8.350 27.780 8.670 27.840 ;
        RECT 44.690 27.780 45.010 27.840 ;
        RECT 8.350 27.640 45.010 27.780 ;
        RECT 8.350 27.580 8.670 27.640 ;
        RECT 44.690 27.580 45.010 27.640 ;
      LAYER via ;
        RECT 44.720 499.840 44.980 500.100 ;
        RECT 415.940 499.840 416.200 500.100 ;
        RECT 8.380 27.580 8.640 27.840 ;
        RECT 44.720 27.580 44.980 27.840 ;
      LAYER met2 ;
        RECT 416.070 510.340 416.350 514.000 ;
        RECT 416.000 510.000 416.350 510.340 ;
        RECT 416.000 500.130 416.140 510.000 ;
        RECT 44.720 499.810 44.980 500.130 ;
        RECT 415.940 499.810 416.200 500.130 ;
        RECT 44.780 27.870 44.920 499.810 ;
        RECT 8.380 27.550 8.640 27.870 ;
        RECT 44.720 27.550 44.980 27.870 ;
        RECT 8.440 2.400 8.580 27.550 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 389.690 496.980 390.010 497.040 ;
        RECT 420.050 496.980 420.370 497.040 ;
        RECT 389.690 496.840 420.370 496.980 ;
        RECT 389.690 496.780 390.010 496.840 ;
        RECT 420.050 496.780 420.370 496.840 ;
        RECT 14.330 44.780 14.650 44.840 ;
        RECT 389.690 44.780 390.010 44.840 ;
        RECT 14.330 44.640 390.010 44.780 ;
        RECT 14.330 44.580 14.650 44.640 ;
        RECT 389.690 44.580 390.010 44.640 ;
      LAYER via ;
        RECT 389.720 496.780 389.980 497.040 ;
        RECT 420.080 496.780 420.340 497.040 ;
        RECT 14.360 44.580 14.620 44.840 ;
        RECT 389.720 44.580 389.980 44.840 ;
      LAYER met2 ;
        RECT 420.210 510.340 420.490 514.000 ;
        RECT 420.140 510.000 420.490 510.340 ;
        RECT 420.140 497.070 420.280 510.000 ;
        RECT 389.720 496.750 389.980 497.070 ;
        RECT 420.080 496.750 420.340 497.070 ;
        RECT 389.780 44.870 389.920 496.750 ;
        RECT 14.360 44.550 14.620 44.870 ;
        RECT 389.720 44.550 389.980 44.870 ;
        RECT 14.420 2.400 14.560 44.550 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 375.890 500.380 376.210 500.440 ;
        RECT 437.070 500.380 437.390 500.440 ;
        RECT 375.890 500.240 437.390 500.380 ;
        RECT 375.890 500.180 376.210 500.240 ;
        RECT 437.070 500.180 437.390 500.240 ;
        RECT 38.250 30.840 38.570 30.900 ;
        RECT 375.890 30.840 376.210 30.900 ;
        RECT 38.250 30.700 376.210 30.840 ;
        RECT 38.250 30.640 38.570 30.700 ;
        RECT 375.890 30.640 376.210 30.700 ;
      LAYER via ;
        RECT 375.920 500.180 376.180 500.440 ;
        RECT 437.100 500.180 437.360 500.440 ;
        RECT 38.280 30.640 38.540 30.900 ;
        RECT 375.920 30.640 376.180 30.900 ;
      LAYER met2 ;
        RECT 437.230 510.340 437.510 514.000 ;
        RECT 437.160 510.000 437.510 510.340 ;
        RECT 437.160 500.470 437.300 510.000 ;
        RECT 375.920 500.150 376.180 500.470 ;
        RECT 437.100 500.150 437.360 500.470 ;
        RECT 375.980 30.930 376.120 500.150 ;
        RECT 38.280 30.610 38.540 30.930 ;
        RECT 375.920 30.610 376.180 30.930 ;
        RECT 38.340 2.400 38.480 30.610 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 51.580 241.430 51.640 ;
        RECT 579.670 51.580 579.990 51.640 ;
        RECT 241.110 51.440 579.990 51.580 ;
        RECT 241.110 51.380 241.430 51.440 ;
        RECT 579.670 51.380 579.990 51.440 ;
      LAYER via ;
        RECT 241.140 51.380 241.400 51.640 ;
        RECT 579.700 51.380 579.960 51.640 ;
      LAYER met2 ;
        RECT 582.590 510.410 582.870 514.000 ;
        RECT 579.760 510.270 582.870 510.410 ;
        RECT 579.760 51.670 579.900 510.270 ;
        RECT 582.590 510.000 582.870 510.270 ;
        RECT 241.140 51.350 241.400 51.670 ;
        RECT 579.700 51.350 579.960 51.670 ;
        RECT 241.200 17.410 241.340 51.350 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 500.040 441.530 500.100 ;
        RECT 594.850 500.040 595.170 500.100 ;
        RECT 441.210 499.900 595.170 500.040 ;
        RECT 441.210 499.840 441.530 499.900 ;
        RECT 594.850 499.840 595.170 499.900 ;
        RECT 261.810 493.240 262.130 493.300 ;
        RECT 441.210 493.240 441.530 493.300 ;
        RECT 261.810 493.100 441.530 493.240 ;
        RECT 261.810 493.040 262.130 493.100 ;
        RECT 441.210 493.040 441.530 493.100 ;
        RECT 258.130 17.240 258.450 17.300 ;
        RECT 261.810 17.240 262.130 17.300 ;
        RECT 258.130 17.100 262.130 17.240 ;
        RECT 258.130 17.040 258.450 17.100 ;
        RECT 261.810 17.040 262.130 17.100 ;
      LAYER via ;
        RECT 441.240 499.840 441.500 500.100 ;
        RECT 594.880 499.840 595.140 500.100 ;
        RECT 261.840 493.040 262.100 493.300 ;
        RECT 441.240 493.040 441.500 493.300 ;
        RECT 258.160 17.040 258.420 17.300 ;
        RECT 261.840 17.040 262.100 17.300 ;
      LAYER met2 ;
        RECT 595.010 510.340 595.290 514.000 ;
        RECT 594.940 510.000 595.290 510.340 ;
        RECT 594.940 500.130 595.080 510.000 ;
        RECT 441.240 499.810 441.500 500.130 ;
        RECT 594.880 499.810 595.140 500.130 ;
        RECT 441.300 493.330 441.440 499.810 ;
        RECT 261.840 493.010 262.100 493.330 ;
        RECT 441.240 493.010 441.500 493.330 ;
        RECT 261.900 17.330 262.040 493.010 ;
        RECT 258.160 17.010 258.420 17.330 ;
        RECT 261.840 17.010 262.100 17.330 ;
        RECT 258.220 2.400 258.360 17.010 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 486.440 282.830 486.500 ;
        RECT 607.730 486.440 608.050 486.500 ;
        RECT 282.510 486.300 608.050 486.440 ;
        RECT 282.510 486.240 282.830 486.300 ;
        RECT 607.730 486.240 608.050 486.300 ;
        RECT 276.070 16.220 276.390 16.280 ;
        RECT 282.510 16.220 282.830 16.280 ;
        RECT 276.070 16.080 282.830 16.220 ;
        RECT 276.070 16.020 276.390 16.080 ;
        RECT 282.510 16.020 282.830 16.080 ;
      LAYER via ;
        RECT 282.540 486.240 282.800 486.500 ;
        RECT 607.760 486.240 608.020 486.500 ;
        RECT 276.100 16.020 276.360 16.280 ;
        RECT 282.540 16.020 282.800 16.280 ;
      LAYER met2 ;
        RECT 607.890 510.340 608.170 514.000 ;
        RECT 607.820 510.000 608.170 510.340 ;
        RECT 607.820 486.530 607.960 510.000 ;
        RECT 282.540 486.210 282.800 486.530 ;
        RECT 607.760 486.210 608.020 486.530 ;
        RECT 282.600 16.310 282.740 486.210 ;
        RECT 276.100 15.990 276.360 16.310 ;
        RECT 282.540 15.990 282.800 16.310 ;
        RECT 276.160 2.400 276.300 15.990 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 614.170 472.840 614.490 472.900 ;
        RECT 619.230 472.840 619.550 472.900 ;
        RECT 614.170 472.700 619.550 472.840 ;
        RECT 614.170 472.640 614.490 472.700 ;
        RECT 619.230 472.640 619.550 472.700 ;
        RECT 296.310 58.720 296.630 58.780 ;
        RECT 614.170 58.720 614.490 58.780 ;
        RECT 296.310 58.580 614.490 58.720 ;
        RECT 296.310 58.520 296.630 58.580 ;
        RECT 614.170 58.520 614.490 58.580 ;
        RECT 294.010 16.900 294.330 16.960 ;
        RECT 296.310 16.900 296.630 16.960 ;
        RECT 294.010 16.760 296.630 16.900 ;
        RECT 294.010 16.700 294.330 16.760 ;
        RECT 296.310 16.700 296.630 16.760 ;
      LAYER via ;
        RECT 614.200 472.640 614.460 472.900 ;
        RECT 619.260 472.640 619.520 472.900 ;
        RECT 296.340 58.520 296.600 58.780 ;
        RECT 614.200 58.520 614.460 58.780 ;
        RECT 294.040 16.700 294.300 16.960 ;
        RECT 296.340 16.700 296.600 16.960 ;
      LAYER met2 ;
        RECT 620.770 510.410 621.050 514.000 ;
        RECT 619.320 510.270 621.050 510.410 ;
        RECT 619.320 472.930 619.460 510.270 ;
        RECT 620.770 510.000 621.050 510.270 ;
        RECT 614.200 472.610 614.460 472.930 ;
        RECT 619.260 472.610 619.520 472.930 ;
        RECT 614.260 58.810 614.400 472.610 ;
        RECT 296.340 58.490 296.600 58.810 ;
        RECT 614.200 58.490 614.460 58.810 ;
        RECT 296.400 16.990 296.540 58.490 ;
        RECT 294.040 16.670 294.300 16.990 ;
        RECT 296.340 16.670 296.600 16.990 ;
        RECT 294.100 2.400 294.240 16.670 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.970 472.840 628.290 472.900 ;
        RECT 632.110 472.840 632.430 472.900 ;
        RECT 627.970 472.700 632.430 472.840 ;
        RECT 627.970 472.640 628.290 472.700 ;
        RECT 632.110 472.640 632.430 472.700 ;
        RECT 317.010 65.520 317.330 65.580 ;
        RECT 627.970 65.520 628.290 65.580 ;
        RECT 317.010 65.380 628.290 65.520 ;
        RECT 317.010 65.320 317.330 65.380 ;
        RECT 627.970 65.320 628.290 65.380 ;
        RECT 311.950 16.900 312.270 16.960 ;
        RECT 317.010 16.900 317.330 16.960 ;
        RECT 311.950 16.760 317.330 16.900 ;
        RECT 311.950 16.700 312.270 16.760 ;
        RECT 317.010 16.700 317.330 16.760 ;
      LAYER via ;
        RECT 628.000 472.640 628.260 472.900 ;
        RECT 632.140 472.640 632.400 472.900 ;
        RECT 317.040 65.320 317.300 65.580 ;
        RECT 628.000 65.320 628.260 65.580 ;
        RECT 311.980 16.700 312.240 16.960 ;
        RECT 317.040 16.700 317.300 16.960 ;
      LAYER met2 ;
        RECT 633.650 510.410 633.930 514.000 ;
        RECT 632.200 510.270 633.930 510.410 ;
        RECT 632.200 472.930 632.340 510.270 ;
        RECT 633.650 510.000 633.930 510.270 ;
        RECT 628.000 472.610 628.260 472.930 ;
        RECT 632.140 472.610 632.400 472.930 ;
        RECT 628.060 65.610 628.200 472.610 ;
        RECT 317.040 65.290 317.300 65.610 ;
        RECT 628.000 65.290 628.260 65.610 ;
        RECT 317.100 16.990 317.240 65.290 ;
        RECT 311.980 16.670 312.240 16.990 ;
        RECT 317.040 16.670 317.300 16.990 ;
        RECT 312.040 2.400 312.180 16.670 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.590 500.040 603.910 500.100 ;
        RECT 646.370 500.040 646.690 500.100 ;
        RECT 603.590 499.900 646.690 500.040 ;
        RECT 603.590 499.840 603.910 499.900 ;
        RECT 646.370 499.840 646.690 499.900 ;
        RECT 330.810 72.320 331.130 72.380 ;
        RECT 603.590 72.320 603.910 72.380 ;
        RECT 330.810 72.180 603.910 72.320 ;
        RECT 330.810 72.120 331.130 72.180 ;
        RECT 603.590 72.120 603.910 72.180 ;
      LAYER via ;
        RECT 603.620 499.840 603.880 500.100 ;
        RECT 646.400 499.840 646.660 500.100 ;
        RECT 330.840 72.120 331.100 72.380 ;
        RECT 603.620 72.120 603.880 72.380 ;
      LAYER met2 ;
        RECT 646.530 510.340 646.810 514.000 ;
        RECT 646.460 510.000 646.810 510.340 ;
        RECT 646.460 500.130 646.600 510.000 ;
        RECT 603.620 499.810 603.880 500.130 ;
        RECT 646.400 499.810 646.660 500.130 ;
        RECT 603.680 72.410 603.820 499.810 ;
        RECT 330.840 72.090 331.100 72.410 ;
        RECT 603.620 72.090 603.880 72.410 ;
        RECT 330.900 17.410 331.040 72.090 ;
        RECT 329.980 17.270 331.040 17.410 ;
        RECT 329.980 2.400 330.120 17.270 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 134.540 351.830 134.600 ;
        RECT 655.570 134.540 655.890 134.600 ;
        RECT 351.510 134.400 655.890 134.540 ;
        RECT 351.510 134.340 351.830 134.400 ;
        RECT 655.570 134.340 655.890 134.400 ;
        RECT 347.370 17.240 347.690 17.300 ;
        RECT 351.510 17.240 351.830 17.300 ;
        RECT 347.370 17.100 351.830 17.240 ;
        RECT 347.370 17.040 347.690 17.100 ;
        RECT 351.510 17.040 351.830 17.100 ;
      LAYER via ;
        RECT 351.540 134.340 351.800 134.600 ;
        RECT 655.600 134.340 655.860 134.600 ;
        RECT 347.400 17.040 347.660 17.300 ;
        RECT 351.540 17.040 351.800 17.300 ;
      LAYER met2 ;
        RECT 659.410 510.410 659.690 514.000 ;
        RECT 655.660 510.270 659.690 510.410 ;
        RECT 655.660 134.630 655.800 510.270 ;
        RECT 659.410 510.000 659.690 510.270 ;
        RECT 351.540 134.310 351.800 134.630 ;
        RECT 655.600 134.310 655.860 134.630 ;
        RECT 351.600 17.330 351.740 134.310 ;
        RECT 347.400 17.010 347.660 17.330 ;
        RECT 351.540 17.010 351.800 17.330 ;
        RECT 347.460 2.400 347.600 17.010 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 479.640 365.630 479.700 ;
        RECT 671.670 479.640 671.990 479.700 ;
        RECT 365.310 479.500 671.990 479.640 ;
        RECT 365.310 479.440 365.630 479.500 ;
        RECT 671.670 479.440 671.990 479.500 ;
      LAYER via ;
        RECT 365.340 479.440 365.600 479.700 ;
        RECT 671.700 479.440 671.960 479.700 ;
      LAYER met2 ;
        RECT 671.830 510.340 672.110 514.000 ;
        RECT 671.760 510.000 672.110 510.340 ;
        RECT 671.760 479.730 671.900 510.000 ;
        RECT 365.340 479.410 365.600 479.730 ;
        RECT 671.700 479.410 671.960 479.730 ;
        RECT 365.400 2.400 365.540 479.410 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 658.790 500.040 659.110 500.100 ;
        RECT 684.550 500.040 684.870 500.100 ;
        RECT 658.790 499.900 684.870 500.040 ;
        RECT 658.790 499.840 659.110 499.900 ;
        RECT 684.550 499.840 684.870 499.900 ;
        RECT 386.010 79.460 386.330 79.520 ;
        RECT 658.790 79.460 659.110 79.520 ;
        RECT 386.010 79.320 659.110 79.460 ;
        RECT 386.010 79.260 386.330 79.320 ;
        RECT 658.790 79.260 659.110 79.320 ;
        RECT 383.250 17.580 383.570 17.640 ;
        RECT 386.010 17.580 386.330 17.640 ;
        RECT 383.250 17.440 386.330 17.580 ;
        RECT 383.250 17.380 383.570 17.440 ;
        RECT 386.010 17.380 386.330 17.440 ;
      LAYER via ;
        RECT 658.820 499.840 659.080 500.100 ;
        RECT 684.580 499.840 684.840 500.100 ;
        RECT 386.040 79.260 386.300 79.520 ;
        RECT 658.820 79.260 659.080 79.520 ;
        RECT 383.280 17.380 383.540 17.640 ;
        RECT 386.040 17.380 386.300 17.640 ;
      LAYER met2 ;
        RECT 684.710 510.340 684.990 514.000 ;
        RECT 684.640 510.000 684.990 510.340 ;
        RECT 684.640 500.130 684.780 510.000 ;
        RECT 658.820 499.810 659.080 500.130 ;
        RECT 684.580 499.810 684.840 500.130 ;
        RECT 658.880 79.550 659.020 499.810 ;
        RECT 386.040 79.230 386.300 79.550 ;
        RECT 658.820 79.230 659.080 79.550 ;
        RECT 386.100 17.670 386.240 79.230 ;
        RECT 383.280 17.350 383.540 17.670 ;
        RECT 386.040 17.350 386.300 17.670 ;
        RECT 383.340 2.400 383.480 17.350 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.710 203.560 407.030 203.620 ;
        RECT 697.430 203.560 697.750 203.620 ;
        RECT 406.710 203.420 697.750 203.560 ;
        RECT 406.710 203.360 407.030 203.420 ;
        RECT 697.430 203.360 697.750 203.420 ;
        RECT 401.190 15.880 401.510 15.940 ;
        RECT 406.710 15.880 407.030 15.940 ;
        RECT 401.190 15.740 407.030 15.880 ;
        RECT 401.190 15.680 401.510 15.740 ;
        RECT 406.710 15.680 407.030 15.740 ;
      LAYER via ;
        RECT 406.740 203.360 407.000 203.620 ;
        RECT 697.460 203.360 697.720 203.620 ;
        RECT 401.220 15.680 401.480 15.940 ;
        RECT 406.740 15.680 407.000 15.940 ;
      LAYER met2 ;
        RECT 697.590 510.340 697.870 514.000 ;
        RECT 697.520 510.000 697.870 510.340 ;
        RECT 697.520 203.650 697.660 510.000 ;
        RECT 406.740 203.330 407.000 203.650 ;
        RECT 697.460 203.330 697.720 203.650 ;
        RECT 406.800 15.970 406.940 203.330 ;
        RECT 401.220 15.650 401.480 15.970 ;
        RECT 406.740 15.650 407.000 15.970 ;
        RECT 401.280 2.400 401.420 15.650 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.610 472.500 68.930 472.560 ;
        RECT 454.090 472.500 454.410 472.560 ;
        RECT 68.610 472.360 454.410 472.500 ;
        RECT 68.610 472.300 68.930 472.360 ;
        RECT 454.090 472.300 454.410 472.360 ;
        RECT 62.170 20.640 62.490 20.700 ;
        RECT 68.610 20.640 68.930 20.700 ;
        RECT 62.170 20.500 68.930 20.640 ;
        RECT 62.170 20.440 62.490 20.500 ;
        RECT 68.610 20.440 68.930 20.500 ;
      LAYER via ;
        RECT 68.640 472.300 68.900 472.560 ;
        RECT 454.120 472.300 454.380 472.560 ;
        RECT 62.200 20.440 62.460 20.700 ;
        RECT 68.640 20.440 68.900 20.700 ;
      LAYER met2 ;
        RECT 454.250 510.340 454.530 514.000 ;
        RECT 454.180 510.000 454.530 510.340 ;
        RECT 454.180 472.590 454.320 510.000 ;
        RECT 68.640 472.270 68.900 472.590 ;
        RECT 454.120 472.270 454.380 472.590 ;
        RECT 68.700 20.730 68.840 472.270 ;
        RECT 62.200 20.410 62.460 20.730 ;
        RECT 68.640 20.410 68.900 20.730 ;
        RECT 62.260 2.400 62.400 20.410 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.870 472.840 704.190 472.900 ;
        RECT 708.470 472.840 708.790 472.900 ;
        RECT 703.870 472.700 708.790 472.840 ;
        RECT 703.870 472.640 704.190 472.700 ;
        RECT 708.470 472.640 708.790 472.700 ;
        RECT 420.510 148.140 420.830 148.200 ;
        RECT 703.870 148.140 704.190 148.200 ;
        RECT 420.510 148.000 704.190 148.140 ;
        RECT 420.510 147.940 420.830 148.000 ;
        RECT 703.870 147.940 704.190 148.000 ;
        RECT 419.130 14.180 419.450 14.240 ;
        RECT 420.510 14.180 420.830 14.240 ;
        RECT 419.130 14.040 420.830 14.180 ;
        RECT 419.130 13.980 419.450 14.040 ;
        RECT 420.510 13.980 420.830 14.040 ;
      LAYER via ;
        RECT 703.900 472.640 704.160 472.900 ;
        RECT 708.500 472.640 708.760 472.900 ;
        RECT 420.540 147.940 420.800 148.200 ;
        RECT 703.900 147.940 704.160 148.200 ;
        RECT 419.160 13.980 419.420 14.240 ;
        RECT 420.540 13.980 420.800 14.240 ;
      LAYER met2 ;
        RECT 710.470 510.410 710.750 514.000 ;
        RECT 708.560 510.270 710.750 510.410 ;
        RECT 708.560 472.930 708.700 510.270 ;
        RECT 710.470 510.000 710.750 510.270 ;
        RECT 703.900 472.610 704.160 472.930 ;
        RECT 708.500 472.610 708.760 472.930 ;
        RECT 703.960 148.230 704.100 472.610 ;
        RECT 420.540 147.910 420.800 148.230 ;
        RECT 703.900 147.910 704.160 148.230 ;
        RECT 420.600 14.270 420.740 147.910 ;
        RECT 419.160 13.950 419.420 14.270 ;
        RECT 420.540 13.950 420.800 14.270 ;
        RECT 419.220 2.400 419.360 13.950 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 458.900 441.530 458.960 ;
        RECT 720.430 458.900 720.750 458.960 ;
        RECT 441.210 458.760 720.750 458.900 ;
        RECT 441.210 458.700 441.530 458.760 ;
        RECT 720.430 458.700 720.750 458.760 ;
        RECT 436.610 14.520 436.930 14.580 ;
        RECT 441.210 14.520 441.530 14.580 ;
        RECT 436.610 14.380 441.530 14.520 ;
        RECT 436.610 14.320 436.930 14.380 ;
        RECT 441.210 14.320 441.530 14.380 ;
      LAYER via ;
        RECT 441.240 458.700 441.500 458.960 ;
        RECT 720.460 458.700 720.720 458.960 ;
        RECT 436.640 14.320 436.900 14.580 ;
        RECT 441.240 14.320 441.500 14.580 ;
      LAYER met2 ;
        RECT 723.350 510.410 723.630 514.000 ;
        RECT 720.520 510.270 723.630 510.410 ;
        RECT 720.520 458.990 720.660 510.270 ;
        RECT 723.350 510.000 723.630 510.270 ;
        RECT 441.240 458.670 441.500 458.990 ;
        RECT 720.460 458.670 720.720 458.990 ;
        RECT 441.300 14.610 441.440 458.670 ;
        RECT 436.640 14.290 436.900 14.610 ;
        RECT 441.240 14.290 441.500 14.610 ;
        RECT 436.700 2.400 436.840 14.290 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 731.470 472.840 731.790 472.900 ;
        RECT 734.230 472.840 734.550 472.900 ;
        RECT 731.470 472.700 734.550 472.840 ;
        RECT 731.470 472.640 731.790 472.700 ;
        RECT 734.230 472.640 734.550 472.700 ;
        RECT 454.550 217.160 454.870 217.220 ;
        RECT 731.470 217.160 731.790 217.220 ;
        RECT 454.550 217.020 731.790 217.160 ;
        RECT 454.550 216.960 454.870 217.020 ;
        RECT 731.470 216.960 731.790 217.020 ;
      LAYER via ;
        RECT 731.500 472.640 731.760 472.900 ;
        RECT 734.260 472.640 734.520 472.900 ;
        RECT 454.580 216.960 454.840 217.220 ;
        RECT 731.500 216.960 731.760 217.220 ;
      LAYER met2 ;
        RECT 736.230 510.410 736.510 514.000 ;
        RECT 734.320 510.270 736.510 510.410 ;
        RECT 734.320 472.930 734.460 510.270 ;
        RECT 736.230 510.000 736.510 510.270 ;
        RECT 731.500 472.610 731.760 472.930 ;
        RECT 734.260 472.610 734.520 472.930 ;
        RECT 731.560 217.250 731.700 472.610 ;
        RECT 454.580 216.930 454.840 217.250 ;
        RECT 731.500 216.930 731.760 217.250 ;
        RECT 454.640 2.400 454.780 216.930 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 86.260 476.030 86.320 ;
        RECT 745.270 86.260 745.590 86.320 ;
        RECT 475.710 86.120 745.590 86.260 ;
        RECT 475.710 86.060 476.030 86.120 ;
        RECT 745.270 86.060 745.590 86.120 ;
        RECT 472.490 17.580 472.810 17.640 ;
        RECT 475.710 17.580 476.030 17.640 ;
        RECT 472.490 17.440 476.030 17.580 ;
        RECT 472.490 17.380 472.810 17.440 ;
        RECT 475.710 17.380 476.030 17.440 ;
      LAYER via ;
        RECT 475.740 86.060 476.000 86.320 ;
        RECT 745.300 86.060 745.560 86.320 ;
        RECT 472.520 17.380 472.780 17.640 ;
        RECT 475.740 17.380 476.000 17.640 ;
      LAYER met2 ;
        RECT 748.650 510.410 748.930 514.000 ;
        RECT 745.360 510.270 748.930 510.410 ;
        RECT 745.360 86.350 745.500 510.270 ;
        RECT 748.650 510.000 748.930 510.270 ;
        RECT 475.740 86.030 476.000 86.350 ;
        RECT 745.300 86.030 745.560 86.350 ;
        RECT 475.800 17.670 475.940 86.030 ;
        RECT 472.520 17.350 472.780 17.670 ;
        RECT 475.740 17.350 476.000 17.670 ;
        RECT 472.580 2.400 472.720 17.350 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 93.060 496.270 93.120 ;
        RECT 759.070 93.060 759.390 93.120 ;
        RECT 495.950 92.920 759.390 93.060 ;
        RECT 495.950 92.860 496.270 92.920 ;
        RECT 759.070 92.860 759.390 92.920 ;
        RECT 490.430 17.580 490.750 17.640 ;
        RECT 495.950 17.580 496.270 17.640 ;
        RECT 490.430 17.440 496.270 17.580 ;
        RECT 490.430 17.380 490.750 17.440 ;
        RECT 495.950 17.380 496.270 17.440 ;
      LAYER via ;
        RECT 495.980 92.860 496.240 93.120 ;
        RECT 759.100 92.860 759.360 93.120 ;
        RECT 490.460 17.380 490.720 17.640 ;
        RECT 495.980 17.380 496.240 17.640 ;
      LAYER met2 ;
        RECT 761.530 510.410 761.810 514.000 ;
        RECT 759.160 510.270 761.810 510.410 ;
        RECT 759.160 93.150 759.300 510.270 ;
        RECT 761.530 510.000 761.810 510.270 ;
        RECT 495.980 92.830 496.240 93.150 ;
        RECT 759.100 92.830 759.360 93.150 ;
        RECT 496.040 17.670 496.180 92.830 ;
        RECT 490.460 17.350 490.720 17.670 ;
        RECT 495.980 17.350 496.240 17.670 ;
        RECT 490.520 2.400 490.660 17.350 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 99.860 510.530 99.920 ;
        RECT 772.870 99.860 773.190 99.920 ;
        RECT 510.210 99.720 773.190 99.860 ;
        RECT 510.210 99.660 510.530 99.720 ;
        RECT 772.870 99.660 773.190 99.720 ;
        RECT 507.910 17.580 508.230 17.640 ;
        RECT 510.210 17.580 510.530 17.640 ;
        RECT 507.910 17.440 510.530 17.580 ;
        RECT 507.910 17.380 508.230 17.440 ;
        RECT 510.210 17.380 510.530 17.440 ;
      LAYER via ;
        RECT 510.240 99.660 510.500 99.920 ;
        RECT 772.900 99.660 773.160 99.920 ;
        RECT 507.940 17.380 508.200 17.640 ;
        RECT 510.240 17.380 510.500 17.640 ;
      LAYER met2 ;
        RECT 774.410 510.410 774.690 514.000 ;
        RECT 772.960 510.270 774.690 510.410 ;
        RECT 772.960 99.950 773.100 510.270 ;
        RECT 774.410 510.000 774.690 510.270 ;
        RECT 510.240 99.630 510.500 99.950 ;
        RECT 772.900 99.630 773.160 99.950 ;
        RECT 510.300 17.670 510.440 99.630 ;
        RECT 507.940 17.350 508.200 17.670 ;
        RECT 510.240 17.350 510.500 17.670 ;
        RECT 508.000 2.400 508.140 17.350 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 782.990 496.980 783.310 497.040 ;
        RECT 787.130 496.980 787.450 497.040 ;
        RECT 782.990 496.840 787.450 496.980 ;
        RECT 782.990 496.780 783.310 496.840 ;
        RECT 787.130 496.780 787.450 496.840 ;
        RECT 530.910 120.600 531.230 120.660 ;
        RECT 782.990 120.600 783.310 120.660 ;
        RECT 530.910 120.460 783.310 120.600 ;
        RECT 530.910 120.400 531.230 120.460 ;
        RECT 782.990 120.400 783.310 120.460 ;
        RECT 525.850 16.900 526.170 16.960 ;
        RECT 530.910 16.900 531.230 16.960 ;
        RECT 525.850 16.760 531.230 16.900 ;
        RECT 525.850 16.700 526.170 16.760 ;
        RECT 530.910 16.700 531.230 16.760 ;
      LAYER via ;
        RECT 783.020 496.780 783.280 497.040 ;
        RECT 787.160 496.780 787.420 497.040 ;
        RECT 530.940 120.400 531.200 120.660 ;
        RECT 783.020 120.400 783.280 120.660 ;
        RECT 525.880 16.700 526.140 16.960 ;
        RECT 530.940 16.700 531.200 16.960 ;
      LAYER met2 ;
        RECT 787.290 510.340 787.570 514.000 ;
        RECT 787.220 510.000 787.570 510.340 ;
        RECT 787.220 497.070 787.360 510.000 ;
        RECT 783.020 496.750 783.280 497.070 ;
        RECT 787.160 496.750 787.420 497.070 ;
        RECT 783.080 120.690 783.220 496.750 ;
        RECT 530.940 120.370 531.200 120.690 ;
        RECT 783.020 120.370 783.280 120.690 ;
        RECT 531.000 16.990 531.140 120.370 ;
        RECT 525.880 16.670 526.140 16.990 ;
        RECT 530.940 16.670 531.200 16.990 ;
        RECT 525.940 2.400 526.080 16.670 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 794.105 144.925 794.275 193.035 ;
      LAYER mcon ;
        RECT 794.105 192.865 794.275 193.035 ;
      LAYER met1 ;
        RECT 794.490 448.700 794.810 448.760 ;
        RECT 798.170 448.700 798.490 448.760 ;
        RECT 794.490 448.560 798.490 448.700 ;
        RECT 794.490 448.500 794.810 448.560 ;
        RECT 798.170 448.500 798.490 448.560 ;
        RECT 794.030 351.940 794.350 352.200 ;
        RECT 794.120 351.460 794.260 351.940 ;
        RECT 794.490 351.460 794.810 351.520 ;
        RECT 794.120 351.320 794.810 351.460 ;
        RECT 794.490 351.260 794.810 351.320 ;
        RECT 794.030 193.020 794.350 193.080 ;
        RECT 793.835 192.880 794.350 193.020 ;
        RECT 794.030 192.820 794.350 192.880 ;
        RECT 794.045 145.080 794.335 145.125 ;
        RECT 794.950 145.080 795.270 145.140 ;
        RECT 794.045 144.940 795.270 145.080 ;
        RECT 794.045 144.895 794.335 144.940 ;
        RECT 794.950 144.880 795.270 144.940 ;
        RECT 544.710 113.800 545.030 113.860 ;
        RECT 795.410 113.800 795.730 113.860 ;
        RECT 544.710 113.660 795.730 113.800 ;
        RECT 544.710 113.600 545.030 113.660 ;
        RECT 795.410 113.600 795.730 113.660 ;
      LAYER via ;
        RECT 794.520 448.500 794.780 448.760 ;
        RECT 798.200 448.500 798.460 448.760 ;
        RECT 794.060 351.940 794.320 352.200 ;
        RECT 794.520 351.260 794.780 351.520 ;
        RECT 794.060 192.820 794.320 193.080 ;
        RECT 794.980 144.880 795.240 145.140 ;
        RECT 544.740 113.600 545.000 113.860 ;
        RECT 795.440 113.600 795.700 113.860 ;
      LAYER met2 ;
        RECT 800.170 510.410 800.450 514.000 ;
        RECT 798.260 510.270 800.450 510.410 ;
        RECT 798.260 448.790 798.400 510.270 ;
        RECT 800.170 510.000 800.450 510.270 ;
        RECT 794.520 448.470 794.780 448.790 ;
        RECT 798.200 448.470 798.460 448.790 ;
        RECT 794.580 400.930 794.720 448.470 ;
        RECT 794.120 400.790 794.720 400.930 ;
        RECT 794.120 352.230 794.260 400.790 ;
        RECT 794.060 351.910 794.320 352.230 ;
        RECT 794.520 351.230 794.780 351.550 ;
        RECT 794.580 207.130 794.720 351.230 ;
        RECT 794.120 206.990 794.720 207.130 ;
        RECT 794.120 193.110 794.260 206.990 ;
        RECT 794.060 192.790 794.320 193.110 ;
        RECT 794.980 144.850 795.240 145.170 ;
        RECT 795.040 144.570 795.180 144.850 ;
        RECT 795.040 144.430 795.640 144.570 ;
        RECT 795.500 113.890 795.640 144.430 ;
        RECT 544.740 113.570 545.000 113.890 ;
        RECT 795.440 113.570 795.700 113.890 ;
        RECT 544.800 3.130 544.940 113.570 ;
        RECT 543.880 2.990 544.940 3.130 ;
        RECT 543.880 2.400 544.020 2.990 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 808.365 96.645 808.535 144.755 ;
      LAYER mcon ;
        RECT 808.365 144.585 808.535 144.755 ;
      LAYER met1 ;
        RECT 808.750 400.760 809.070 400.820 ;
        RECT 808.380 400.620 809.070 400.760 ;
        RECT 808.380 400.480 808.520 400.620 ;
        RECT 808.750 400.560 809.070 400.620 ;
        RECT 808.290 400.220 808.610 400.480 ;
        RECT 808.290 352.280 808.610 352.540 ;
        RECT 808.380 351.180 808.520 352.280 ;
        RECT 808.290 350.920 808.610 351.180 ;
        RECT 808.290 144.740 808.610 144.800 ;
        RECT 808.095 144.600 808.610 144.740 ;
        RECT 808.290 144.540 808.610 144.600 ;
        RECT 808.305 96.800 808.595 96.845 ;
        RECT 809.210 96.800 809.530 96.860 ;
        RECT 808.305 96.660 809.530 96.800 ;
        RECT 808.305 96.615 808.595 96.660 ;
        RECT 809.210 96.600 809.530 96.660 ;
        RECT 561.730 30.840 562.050 30.900 ;
        RECT 809.210 30.840 809.530 30.900 ;
        RECT 561.730 30.700 809.530 30.840 ;
        RECT 561.730 30.640 562.050 30.700 ;
        RECT 809.210 30.640 809.530 30.700 ;
      LAYER via ;
        RECT 808.780 400.560 809.040 400.820 ;
        RECT 808.320 400.220 808.580 400.480 ;
        RECT 808.320 352.280 808.580 352.540 ;
        RECT 808.320 350.920 808.580 351.180 ;
        RECT 808.320 144.540 808.580 144.800 ;
        RECT 809.240 96.600 809.500 96.860 ;
        RECT 561.760 30.640 562.020 30.900 ;
        RECT 809.240 30.640 809.500 30.900 ;
      LAYER met2 ;
        RECT 813.050 510.410 813.330 514.000 ;
        RECT 810.680 510.270 813.330 510.410 ;
        RECT 810.680 449.210 810.820 510.270 ;
        RECT 813.050 510.000 813.330 510.270 ;
        RECT 808.840 449.070 810.820 449.210 ;
        RECT 808.840 400.850 808.980 449.070 ;
        RECT 808.780 400.530 809.040 400.850 ;
        RECT 808.320 400.190 808.580 400.510 ;
        RECT 808.380 352.570 808.520 400.190 ;
        RECT 808.320 352.250 808.580 352.570 ;
        RECT 808.320 350.890 808.580 351.210 ;
        RECT 808.380 207.130 808.520 350.890 ;
        RECT 807.920 206.990 808.520 207.130 ;
        RECT 807.920 177.890 808.060 206.990 ;
        RECT 807.920 177.750 808.520 177.890 ;
        RECT 808.380 144.830 808.520 177.750 ;
        RECT 808.320 144.510 808.580 144.830 ;
        RECT 809.240 96.570 809.500 96.890 ;
        RECT 809.300 30.930 809.440 96.570 ;
        RECT 561.760 30.610 562.020 30.930 ;
        RECT 809.240 30.610 809.500 30.930 ;
        RECT 561.820 2.400 561.960 30.610 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 822.165 379.525 822.335 427.635 ;
        RECT 821.705 338.045 821.875 362.355 ;
      LAYER mcon ;
        RECT 822.165 427.465 822.335 427.635 ;
        RECT 821.705 362.185 821.875 362.355 ;
      LAYER met1 ;
        RECT 822.090 476.240 822.410 476.300 ;
        RECT 825.770 476.240 826.090 476.300 ;
        RECT 822.090 476.100 826.090 476.240 ;
        RECT 822.090 476.040 822.410 476.100 ;
        RECT 825.770 476.040 826.090 476.100 ;
        RECT 822.090 427.620 822.410 427.680 ;
        RECT 821.895 427.480 822.410 427.620 ;
        RECT 822.090 427.420 822.410 427.480 ;
        RECT 822.090 379.680 822.410 379.740 ;
        RECT 821.895 379.540 822.410 379.680 ;
        RECT 822.090 379.480 822.410 379.540 ;
        RECT 821.645 362.340 821.935 362.385 ;
        RECT 822.090 362.340 822.410 362.400 ;
        RECT 821.645 362.200 822.410 362.340 ;
        RECT 821.645 362.155 821.935 362.200 ;
        RECT 822.090 362.140 822.410 362.200 ;
        RECT 821.630 338.200 821.950 338.260 ;
        RECT 821.435 338.060 821.950 338.200 ;
        RECT 821.630 338.000 821.950 338.060 ;
        RECT 586.110 182.820 586.430 182.880 ;
        RECT 821.630 182.820 821.950 182.880 ;
        RECT 586.110 182.680 821.950 182.820 ;
        RECT 586.110 182.620 586.430 182.680 ;
        RECT 821.630 182.620 821.950 182.680 ;
        RECT 579.670 20.640 579.990 20.700 ;
        RECT 586.110 20.640 586.430 20.700 ;
        RECT 579.670 20.500 586.430 20.640 ;
        RECT 579.670 20.440 579.990 20.500 ;
        RECT 586.110 20.440 586.430 20.500 ;
      LAYER via ;
        RECT 822.120 476.040 822.380 476.300 ;
        RECT 825.800 476.040 826.060 476.300 ;
        RECT 822.120 427.420 822.380 427.680 ;
        RECT 822.120 379.480 822.380 379.740 ;
        RECT 822.120 362.140 822.380 362.400 ;
        RECT 821.660 338.000 821.920 338.260 ;
        RECT 586.140 182.620 586.400 182.880 ;
        RECT 821.660 182.620 821.920 182.880 ;
        RECT 579.700 20.440 579.960 20.700 ;
        RECT 586.140 20.440 586.400 20.700 ;
      LAYER met2 ;
        RECT 825.930 510.340 826.210 514.000 ;
        RECT 825.860 510.000 826.210 510.340 ;
        RECT 825.860 476.330 826.000 510.000 ;
        RECT 822.120 476.010 822.380 476.330 ;
        RECT 825.800 476.010 826.060 476.330 ;
        RECT 822.180 427.710 822.320 476.010 ;
        RECT 822.120 427.390 822.380 427.710 ;
        RECT 822.120 379.450 822.380 379.770 ;
        RECT 822.180 362.430 822.320 379.450 ;
        RECT 822.120 362.110 822.380 362.430 ;
        RECT 821.660 337.970 821.920 338.290 ;
        RECT 821.720 337.805 821.860 337.970 ;
        RECT 821.650 337.435 821.930 337.805 ;
        RECT 822.110 336.755 822.390 337.125 ;
        RECT 822.180 207.130 822.320 336.755 ;
        RECT 821.720 206.990 822.320 207.130 ;
        RECT 821.720 182.910 821.860 206.990 ;
        RECT 586.140 182.590 586.400 182.910 ;
        RECT 821.660 182.590 821.920 182.910 ;
        RECT 586.200 20.730 586.340 182.590 ;
        RECT 579.700 20.410 579.960 20.730 ;
        RECT 586.140 20.410 586.400 20.730 ;
        RECT 579.760 2.400 579.900 20.410 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 821.650 337.480 821.930 337.760 ;
        RECT 822.110 336.800 822.390 337.080 ;
      LAYER met3 ;
        RECT 821.625 337.770 821.955 337.785 ;
        RECT 820.950 337.470 821.955 337.770 ;
        RECT 820.950 337.090 821.250 337.470 ;
        RECT 821.625 337.455 821.955 337.470 ;
        RECT 822.085 337.090 822.415 337.105 ;
        RECT 820.950 336.790 822.415 337.090 ;
        RECT 822.085 336.775 822.415 336.790 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 458.690 496.980 459.010 497.040 ;
        RECT 471.110 496.980 471.430 497.040 ;
        RECT 458.690 496.840 471.430 496.980 ;
        RECT 458.690 496.780 459.010 496.840 ;
        RECT 471.110 496.780 471.430 496.840 ;
        RECT 89.310 396.680 89.630 396.740 ;
        RECT 458.690 396.680 459.010 396.740 ;
        RECT 89.310 396.540 459.010 396.680 ;
        RECT 89.310 396.480 89.630 396.540 ;
        RECT 458.690 396.480 459.010 396.540 ;
        RECT 86.090 20.640 86.410 20.700 ;
        RECT 89.310 20.640 89.630 20.700 ;
        RECT 86.090 20.500 89.630 20.640 ;
        RECT 86.090 20.440 86.410 20.500 ;
        RECT 89.310 20.440 89.630 20.500 ;
      LAYER via ;
        RECT 458.720 496.780 458.980 497.040 ;
        RECT 471.140 496.780 471.400 497.040 ;
        RECT 89.340 396.480 89.600 396.740 ;
        RECT 458.720 396.480 458.980 396.740 ;
        RECT 86.120 20.440 86.380 20.700 ;
        RECT 89.340 20.440 89.600 20.700 ;
      LAYER met2 ;
        RECT 471.270 510.340 471.550 514.000 ;
        RECT 471.200 510.000 471.550 510.340 ;
        RECT 471.200 497.070 471.340 510.000 ;
        RECT 458.720 496.750 458.980 497.070 ;
        RECT 471.140 496.750 471.400 497.070 ;
        RECT 458.780 396.770 458.920 496.750 ;
        RECT 89.340 396.450 89.600 396.770 ;
        RECT 458.720 396.450 458.980 396.770 ;
        RECT 89.400 20.730 89.540 396.450 ;
        RECT 86.120 20.410 86.380 20.730 ;
        RECT 89.340 20.410 89.600 20.730 ;
        RECT 86.180 2.400 86.320 20.410 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 189.620 600.230 189.680 ;
        RECT 834.970 189.620 835.290 189.680 ;
        RECT 599.910 189.480 835.290 189.620 ;
        RECT 599.910 189.420 600.230 189.480 ;
        RECT 834.970 189.420 835.290 189.480 ;
        RECT 597.150 16.900 597.470 16.960 ;
        RECT 599.910 16.900 600.230 16.960 ;
        RECT 597.150 16.760 600.230 16.900 ;
        RECT 597.150 16.700 597.470 16.760 ;
        RECT 599.910 16.700 600.230 16.760 ;
      LAYER via ;
        RECT 599.940 189.420 600.200 189.680 ;
        RECT 835.000 189.420 835.260 189.680 ;
        RECT 597.180 16.700 597.440 16.960 ;
        RECT 599.940 16.700 600.200 16.960 ;
      LAYER met2 ;
        RECT 838.350 510.410 838.630 514.000 ;
        RECT 835.060 510.270 838.630 510.410 ;
        RECT 835.060 189.710 835.200 510.270 ;
        RECT 838.350 510.000 838.630 510.270 ;
        RECT 599.940 189.390 600.200 189.710 ;
        RECT 835.000 189.390 835.260 189.710 ;
        RECT 600.000 16.990 600.140 189.390 ;
        RECT 597.180 16.670 597.440 16.990 ;
        RECT 599.940 16.670 600.200 16.990 ;
        RECT 597.240 2.400 597.380 16.670 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 245.040 620.930 245.100 ;
        RECT 848.770 245.040 849.090 245.100 ;
        RECT 620.610 244.900 849.090 245.040 ;
        RECT 620.610 244.840 620.930 244.900 ;
        RECT 848.770 244.840 849.090 244.900 ;
        RECT 615.090 16.900 615.410 16.960 ;
        RECT 620.610 16.900 620.930 16.960 ;
        RECT 615.090 16.760 620.930 16.900 ;
        RECT 615.090 16.700 615.410 16.760 ;
        RECT 620.610 16.700 620.930 16.760 ;
      LAYER via ;
        RECT 620.640 244.840 620.900 245.100 ;
        RECT 848.800 244.840 849.060 245.100 ;
        RECT 615.120 16.700 615.380 16.960 ;
        RECT 620.640 16.700 620.900 16.960 ;
      LAYER met2 ;
        RECT 851.230 510.410 851.510 514.000 ;
        RECT 848.860 510.270 851.510 510.410 ;
        RECT 848.860 245.130 849.000 510.270 ;
        RECT 851.230 510.000 851.510 510.270 ;
        RECT 620.640 244.810 620.900 245.130 ;
        RECT 848.800 244.810 849.060 245.130 ;
        RECT 620.700 16.990 620.840 244.810 ;
        RECT 615.120 16.670 615.380 16.990 ;
        RECT 620.640 16.670 620.900 16.990 ;
        RECT 615.180 2.400 615.320 16.670 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 465.700 110.330 465.760 ;
        RECT 485.830 465.700 486.150 465.760 ;
        RECT 110.010 465.560 486.150 465.700 ;
        RECT 110.010 465.500 110.330 465.560 ;
        RECT 485.830 465.500 486.150 465.560 ;
      LAYER via ;
        RECT 110.040 465.500 110.300 465.760 ;
        RECT 485.860 465.500 486.120 465.760 ;
      LAYER met2 ;
        RECT 488.750 510.410 489.030 514.000 ;
        RECT 485.920 510.270 489.030 510.410 ;
        RECT 485.920 465.790 486.060 510.270 ;
        RECT 488.750 510.000 489.030 510.270 ;
        RECT 110.040 465.470 110.300 465.790 ;
        RECT 485.860 465.470 486.120 465.790 ;
        RECT 110.100 14.010 110.240 465.470 ;
        RECT 109.640 13.870 110.240 14.010 ;
        RECT 109.640 2.400 109.780 13.870 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 451.760 137.930 451.820 ;
        RECT 504.230 451.760 504.550 451.820 ;
        RECT 137.610 451.620 504.550 451.760 ;
        RECT 137.610 451.560 137.930 451.620 ;
        RECT 504.230 451.560 504.550 451.620 ;
        RECT 133.470 15.540 133.790 15.600 ;
        RECT 137.610 15.540 137.930 15.600 ;
        RECT 133.470 15.400 137.930 15.540 ;
        RECT 133.470 15.340 133.790 15.400 ;
        RECT 137.610 15.340 137.930 15.400 ;
      LAYER via ;
        RECT 137.640 451.560 137.900 451.820 ;
        RECT 504.260 451.560 504.520 451.820 ;
        RECT 133.500 15.340 133.760 15.600 ;
        RECT 137.640 15.340 137.900 15.600 ;
      LAYER met2 ;
        RECT 505.770 510.410 506.050 514.000 ;
        RECT 504.320 510.270 506.050 510.410 ;
        RECT 504.320 451.850 504.460 510.270 ;
        RECT 505.770 510.000 506.050 510.270 ;
        RECT 137.640 451.530 137.900 451.850 ;
        RECT 504.260 451.530 504.520 451.850 ;
        RECT 137.700 15.630 137.840 451.530 ;
        RECT 133.500 15.310 133.760 15.630 ;
        RECT 137.640 15.310 137.900 15.630 ;
        RECT 133.560 2.400 133.700 15.310 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 150.950 113.800 151.270 113.860 ;
        RECT 517.570 113.800 517.890 113.860 ;
        RECT 150.950 113.660 517.890 113.800 ;
        RECT 150.950 113.600 151.270 113.660 ;
        RECT 517.570 113.600 517.890 113.660 ;
      LAYER via ;
        RECT 150.980 113.600 151.240 113.860 ;
        RECT 517.600 113.600 517.860 113.860 ;
      LAYER met2 ;
        RECT 518.190 510.410 518.470 514.000 ;
        RECT 517.660 510.270 518.470 510.410 ;
        RECT 517.660 113.890 517.800 510.270 ;
        RECT 518.190 510.000 518.470 510.270 ;
        RECT 150.980 113.570 151.240 113.890 ;
        RECT 517.600 113.570 517.860 113.890 ;
        RECT 151.040 18.090 151.180 113.570 ;
        RECT 151.040 17.950 151.640 18.090 ;
        RECT 151.500 2.400 151.640 17.950 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 444.960 172.430 445.020 ;
        RECT 527.690 444.960 528.010 445.020 ;
        RECT 172.110 444.820 528.010 444.960 ;
        RECT 172.110 444.760 172.430 444.820 ;
        RECT 527.690 444.760 528.010 444.820 ;
        RECT 169.350 20.640 169.670 20.700 ;
        RECT 172.110 20.640 172.430 20.700 ;
        RECT 169.350 20.500 172.430 20.640 ;
        RECT 169.350 20.440 169.670 20.500 ;
        RECT 172.110 20.440 172.430 20.500 ;
      LAYER via ;
        RECT 172.140 444.760 172.400 445.020 ;
        RECT 527.720 444.760 527.980 445.020 ;
        RECT 169.380 20.440 169.640 20.700 ;
        RECT 172.140 20.440 172.400 20.700 ;
      LAYER met2 ;
        RECT 531.070 510.340 531.350 514.000 ;
        RECT 531.000 510.000 531.350 510.340 ;
        RECT 531.000 483.325 531.140 510.000 ;
        RECT 527.710 482.955 527.990 483.325 ;
        RECT 530.930 482.955 531.210 483.325 ;
        RECT 527.780 445.050 527.920 482.955 ;
        RECT 172.140 444.730 172.400 445.050 ;
        RECT 527.720 444.730 527.980 445.050 ;
        RECT 172.200 20.730 172.340 444.730 ;
        RECT 169.380 20.410 169.640 20.730 ;
        RECT 172.140 20.410 172.400 20.730 ;
        RECT 169.440 2.400 169.580 20.410 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 527.710 483.000 527.990 483.280 ;
        RECT 530.930 483.000 531.210 483.280 ;
      LAYER met3 ;
        RECT 527.685 483.290 528.015 483.305 ;
        RECT 530.905 483.290 531.235 483.305 ;
        RECT 527.685 482.990 531.235 483.290 ;
        RECT 527.685 482.975 528.015 482.990 ;
        RECT 530.905 482.975 531.235 482.990 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 438.160 193.130 438.220 ;
        RECT 541.490 438.160 541.810 438.220 ;
        RECT 192.810 438.020 541.810 438.160 ;
        RECT 192.810 437.960 193.130 438.020 ;
        RECT 541.490 437.960 541.810 438.020 ;
        RECT 186.830 20.640 187.150 20.700 ;
        RECT 192.810 20.640 193.130 20.700 ;
        RECT 186.830 20.500 193.130 20.640 ;
        RECT 186.830 20.440 187.150 20.500 ;
        RECT 192.810 20.440 193.130 20.500 ;
      LAYER via ;
        RECT 192.840 437.960 193.100 438.220 ;
        RECT 541.520 437.960 541.780 438.220 ;
        RECT 186.860 20.440 187.120 20.700 ;
        RECT 192.840 20.440 193.100 20.700 ;
      LAYER met2 ;
        RECT 543.950 510.340 544.230 514.000 ;
        RECT 543.880 510.000 544.230 510.340 ;
        RECT 543.880 483.325 544.020 510.000 ;
        RECT 541.510 482.955 541.790 483.325 ;
        RECT 543.810 482.955 544.090 483.325 ;
        RECT 541.580 438.250 541.720 482.955 ;
        RECT 192.840 437.930 193.100 438.250 ;
        RECT 541.520 437.930 541.780 438.250 ;
        RECT 192.900 20.730 193.040 437.930 ;
        RECT 186.860 20.410 187.120 20.730 ;
        RECT 192.840 20.410 193.100 20.730 ;
        RECT 186.920 2.400 187.060 20.410 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 541.510 483.000 541.790 483.280 ;
        RECT 543.810 483.000 544.090 483.280 ;
      LAYER met3 ;
        RECT 541.485 483.290 541.815 483.305 ;
        RECT 543.785 483.290 544.115 483.305 ;
        RECT 541.485 482.990 544.115 483.290 ;
        RECT 541.485 482.975 541.815 482.990 ;
        RECT 543.785 482.975 544.115 482.990 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 552.605 386.325 552.775 434.775 ;
        RECT 553.525 241.485 553.695 289.595 ;
      LAYER mcon ;
        RECT 552.605 434.605 552.775 434.775 ;
        RECT 553.525 289.425 553.695 289.595 ;
      LAYER met1 ;
        RECT 552.545 434.760 552.835 434.805 ;
        RECT 552.990 434.760 553.310 434.820 ;
        RECT 552.545 434.620 553.310 434.760 ;
        RECT 552.545 434.575 552.835 434.620 ;
        RECT 552.990 434.560 553.310 434.620 ;
        RECT 552.530 386.480 552.850 386.540 ;
        RECT 552.335 386.340 552.850 386.480 ;
        RECT 552.530 386.280 552.850 386.340 ;
        RECT 552.530 338.200 552.850 338.260 ;
        RECT 552.990 338.200 553.310 338.260 ;
        RECT 552.530 338.060 553.310 338.200 ;
        RECT 552.530 338.000 552.850 338.060 ;
        RECT 552.990 338.000 553.310 338.060 ;
        RECT 553.450 289.580 553.770 289.640 ;
        RECT 553.255 289.440 553.770 289.580 ;
        RECT 553.450 289.380 553.770 289.440 ;
        RECT 553.465 241.640 553.755 241.685 ;
        RECT 553.910 241.640 554.230 241.700 ;
        RECT 553.465 241.500 554.230 241.640 ;
        RECT 553.465 241.455 553.755 241.500 ;
        RECT 553.910 241.440 554.230 241.500 ;
        RECT 553.450 193.360 553.770 193.420 ;
        RECT 553.910 193.360 554.230 193.420 ;
        RECT 553.450 193.220 554.230 193.360 ;
        RECT 553.450 193.160 553.770 193.220 ;
        RECT 553.910 193.160 554.230 193.220 ;
        RECT 206.610 127.740 206.930 127.800 ;
        RECT 553.450 127.740 553.770 127.800 ;
        RECT 206.610 127.600 553.770 127.740 ;
        RECT 206.610 127.540 206.930 127.600 ;
        RECT 553.450 127.540 553.770 127.600 ;
        RECT 204.770 14.180 205.090 14.240 ;
        RECT 206.610 14.180 206.930 14.240 ;
        RECT 204.770 14.040 206.930 14.180 ;
        RECT 204.770 13.980 205.090 14.040 ;
        RECT 206.610 13.980 206.930 14.040 ;
      LAYER via ;
        RECT 553.020 434.560 553.280 434.820 ;
        RECT 552.560 386.280 552.820 386.540 ;
        RECT 552.560 338.000 552.820 338.260 ;
        RECT 553.020 338.000 553.280 338.260 ;
        RECT 553.480 289.380 553.740 289.640 ;
        RECT 553.940 241.440 554.200 241.700 ;
        RECT 553.480 193.160 553.740 193.420 ;
        RECT 553.940 193.160 554.200 193.420 ;
        RECT 206.640 127.540 206.900 127.800 ;
        RECT 553.480 127.540 553.740 127.800 ;
        RECT 204.800 13.980 205.060 14.240 ;
        RECT 206.640 13.980 206.900 14.240 ;
      LAYER met2 ;
        RECT 556.830 510.410 557.110 514.000 ;
        RECT 554.920 510.270 557.110 510.410 ;
        RECT 554.920 449.210 555.060 510.270 ;
        RECT 556.830 510.000 557.110 510.270 ;
        RECT 554.000 449.070 555.060 449.210 ;
        RECT 554.000 448.530 554.140 449.070 ;
        RECT 553.080 448.390 554.140 448.530 ;
        RECT 553.080 434.850 553.220 448.390 ;
        RECT 553.020 434.530 553.280 434.850 ;
        RECT 552.560 386.250 552.820 386.570 ;
        RECT 552.620 338.290 552.760 386.250 ;
        RECT 552.560 337.970 552.820 338.290 ;
        RECT 553.020 337.970 553.280 338.290 ;
        RECT 553.080 303.010 553.220 337.970 ;
        RECT 553.080 302.870 553.680 303.010 ;
        RECT 553.540 289.670 553.680 302.870 ;
        RECT 553.480 289.350 553.740 289.670 ;
        RECT 553.940 241.410 554.200 241.730 ;
        RECT 554.000 193.450 554.140 241.410 ;
        RECT 553.480 193.130 553.740 193.450 ;
        RECT 553.940 193.130 554.200 193.450 ;
        RECT 553.540 127.830 553.680 193.130 ;
        RECT 206.640 127.510 206.900 127.830 ;
        RECT 553.480 127.510 553.740 127.830 ;
        RECT 206.700 14.270 206.840 127.510 ;
        RECT 204.800 13.950 205.060 14.270 ;
        RECT 206.640 13.950 206.900 14.270 ;
        RECT 204.860 2.400 205.000 13.950 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.870 255.240 566.190 255.300 ;
        RECT 566.790 255.240 567.110 255.300 ;
        RECT 565.870 255.100 567.110 255.240 ;
        RECT 565.870 255.040 566.190 255.100 ;
        RECT 566.790 255.040 567.110 255.100 ;
        RECT 566.790 207.100 567.110 207.360 ;
        RECT 566.880 206.680 567.020 207.100 ;
        RECT 566.790 206.420 567.110 206.680 ;
        RECT 227.310 141.340 227.630 141.400 ;
        RECT 566.790 141.340 567.110 141.400 ;
        RECT 227.310 141.200 567.110 141.340 ;
        RECT 227.310 141.140 227.630 141.200 ;
        RECT 566.790 141.140 567.110 141.200 ;
        RECT 222.710 20.640 223.030 20.700 ;
        RECT 227.310 20.640 227.630 20.700 ;
        RECT 222.710 20.500 227.630 20.640 ;
        RECT 222.710 20.440 223.030 20.500 ;
        RECT 227.310 20.440 227.630 20.500 ;
      LAYER via ;
        RECT 565.900 255.040 566.160 255.300 ;
        RECT 566.820 255.040 567.080 255.300 ;
        RECT 566.820 207.100 567.080 207.360 ;
        RECT 566.820 206.420 567.080 206.680 ;
        RECT 227.340 141.140 227.600 141.400 ;
        RECT 566.820 141.140 567.080 141.400 ;
        RECT 222.740 20.440 223.000 20.700 ;
        RECT 227.340 20.440 227.600 20.700 ;
      LAYER met2 ;
        RECT 569.710 510.410 569.990 514.000 ;
        RECT 567.340 510.270 569.990 510.410 ;
        RECT 567.340 449.210 567.480 510.270 ;
        RECT 569.710 510.000 569.990 510.270 ;
        RECT 566.880 449.070 567.480 449.210 ;
        RECT 566.880 351.970 567.020 449.070 ;
        RECT 565.960 351.830 567.020 351.970 ;
        RECT 565.960 351.290 566.100 351.830 ;
        RECT 565.960 351.150 566.560 351.290 ;
        RECT 566.420 255.410 566.560 351.150 ;
        RECT 565.960 255.330 566.560 255.410 ;
        RECT 565.900 255.270 566.560 255.330 ;
        RECT 565.900 255.010 566.160 255.270 ;
        RECT 566.820 255.010 567.080 255.330 ;
        RECT 565.960 254.855 566.100 255.010 ;
        RECT 566.880 207.390 567.020 255.010 ;
        RECT 566.820 207.070 567.080 207.390 ;
        RECT 566.820 206.390 567.080 206.710 ;
        RECT 566.880 141.430 567.020 206.390 ;
        RECT 227.340 141.110 227.600 141.430 ;
        RECT 566.820 141.110 567.080 141.430 ;
        RECT 227.400 20.730 227.540 141.110 ;
        RECT 222.740 20.410 223.000 20.730 ;
        RECT 227.340 20.410 227.600 20.730 ;
        RECT 222.800 2.400 222.940 20.410 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 86.260 45.470 86.320 ;
        RECT 420.970 86.260 421.290 86.320 ;
        RECT 45.150 86.120 421.290 86.260 ;
        RECT 45.150 86.060 45.470 86.120 ;
        RECT 420.970 86.060 421.290 86.120 ;
        RECT 20.310 20.300 20.630 20.360 ;
        RECT 45.150 20.300 45.470 20.360 ;
        RECT 20.310 20.160 45.470 20.300 ;
        RECT 20.310 20.100 20.630 20.160 ;
        RECT 45.150 20.100 45.470 20.160 ;
      LAYER via ;
        RECT 45.180 86.060 45.440 86.320 ;
        RECT 421.000 86.060 421.260 86.320 ;
        RECT 20.340 20.100 20.600 20.360 ;
        RECT 45.180 20.100 45.440 20.360 ;
      LAYER met2 ;
        RECT 424.350 510.410 424.630 514.000 ;
        RECT 421.060 510.270 424.630 510.410 ;
        RECT 421.060 86.350 421.200 510.270 ;
        RECT 424.350 510.000 424.630 510.270 ;
        RECT 45.180 86.030 45.440 86.350 ;
        RECT 421.000 86.030 421.260 86.350 ;
        RECT 45.240 20.390 45.380 86.030 ;
        RECT 20.340 20.070 20.600 20.390 ;
        RECT 45.180 20.070 45.440 20.390 ;
        RECT 20.400 2.400 20.540 20.070 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 435.765 282.965 435.935 331.075 ;
      LAYER mcon ;
        RECT 435.765 330.905 435.935 331.075 ;
      LAYER met1 ;
        RECT 436.150 386.480 436.470 386.540 ;
        RECT 437.990 386.480 438.310 386.540 ;
        RECT 436.150 386.340 438.310 386.480 ;
        RECT 436.150 386.280 436.470 386.340 ;
        RECT 437.990 386.280 438.310 386.340 ;
        RECT 435.690 331.060 436.010 331.120 ;
        RECT 435.495 330.920 436.010 331.060 ;
        RECT 435.690 330.860 436.010 330.920 ;
        RECT 435.690 283.120 436.010 283.180 ;
        RECT 435.495 282.980 436.010 283.120 ;
        RECT 435.690 282.920 436.010 282.980 ;
        RECT 52.050 245.040 52.370 245.100 ;
        RECT 435.690 245.040 436.010 245.100 ;
        RECT 52.050 244.900 436.010 245.040 ;
        RECT 52.050 244.840 52.370 244.900 ;
        RECT 435.690 244.840 436.010 244.900 ;
        RECT 44.230 20.640 44.550 20.700 ;
        RECT 52.050 20.640 52.370 20.700 ;
        RECT 44.230 20.500 52.370 20.640 ;
        RECT 44.230 20.440 44.550 20.500 ;
        RECT 52.050 20.440 52.370 20.500 ;
      LAYER via ;
        RECT 436.180 386.280 436.440 386.540 ;
        RECT 438.020 386.280 438.280 386.540 ;
        RECT 435.720 330.860 435.980 331.120 ;
        RECT 435.720 282.920 435.980 283.180 ;
        RECT 52.080 244.840 52.340 245.100 ;
        RECT 435.720 244.840 435.980 245.100 ;
        RECT 44.260 20.440 44.520 20.700 ;
        RECT 52.080 20.440 52.340 20.700 ;
      LAYER met2 ;
        RECT 441.370 510.410 441.650 514.000 ;
        RECT 439.000 510.270 441.650 510.410 ;
        RECT 439.000 449.210 439.140 510.270 ;
        RECT 441.370 510.000 441.650 510.270 ;
        RECT 438.080 449.070 439.140 449.210 ;
        RECT 438.080 386.570 438.220 449.070 ;
        RECT 436.180 386.250 436.440 386.570 ;
        RECT 438.020 386.250 438.280 386.570 ;
        RECT 436.240 331.570 436.380 386.250 ;
        RECT 435.780 331.430 436.380 331.570 ;
        RECT 435.780 331.150 435.920 331.430 ;
        RECT 435.720 330.830 435.980 331.150 ;
        RECT 435.720 282.890 435.980 283.210 ;
        RECT 435.780 245.130 435.920 282.890 ;
        RECT 52.080 244.810 52.340 245.130 ;
        RECT 435.720 244.810 435.980 245.130 ;
        RECT 52.140 20.730 52.280 244.810 ;
        RECT 44.260 20.410 44.520 20.730 ;
        RECT 52.080 20.410 52.340 20.730 ;
        RECT 44.320 2.400 44.460 20.410 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 431.360 248.330 431.420 ;
        RECT 587.030 431.360 587.350 431.420 ;
        RECT 248.010 431.220 587.350 431.360 ;
        RECT 248.010 431.160 248.330 431.220 ;
        RECT 587.030 431.160 587.350 431.220 ;
      LAYER via ;
        RECT 248.040 431.160 248.300 431.420 ;
        RECT 587.060 431.160 587.320 431.420 ;
      LAYER met2 ;
        RECT 586.730 510.340 587.010 514.000 ;
        RECT 586.660 510.000 587.010 510.340 ;
        RECT 586.660 473.690 586.800 510.000 ;
        RECT 586.660 473.550 587.260 473.690 ;
        RECT 587.120 431.450 587.260 473.550 ;
        RECT 248.040 431.130 248.300 431.450 ;
        RECT 587.060 431.130 587.320 431.450 ;
        RECT 248.100 16.730 248.240 431.130 ;
        RECT 246.720 16.590 248.240 16.730 ;
        RECT 246.720 2.400 246.860 16.590 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.930 448.700 594.250 448.760 ;
        RECT 597.610 448.700 597.930 448.760 ;
        RECT 593.930 448.560 597.930 448.700 ;
        RECT 593.930 448.500 594.250 448.560 ;
        RECT 597.610 448.500 597.930 448.560 ;
        RECT 268.710 424.220 269.030 424.280 ;
        RECT 593.930 424.220 594.250 424.280 ;
        RECT 268.710 424.080 594.250 424.220 ;
        RECT 268.710 424.020 269.030 424.080 ;
        RECT 593.930 424.020 594.250 424.080 ;
        RECT 264.110 17.240 264.430 17.300 ;
        RECT 268.710 17.240 269.030 17.300 ;
        RECT 264.110 17.100 269.030 17.240 ;
        RECT 264.110 17.040 264.430 17.100 ;
        RECT 268.710 17.040 269.030 17.100 ;
      LAYER via ;
        RECT 593.960 448.500 594.220 448.760 ;
        RECT 597.640 448.500 597.900 448.760 ;
        RECT 268.740 424.020 269.000 424.280 ;
        RECT 593.960 424.020 594.220 424.280 ;
        RECT 264.140 17.040 264.400 17.300 ;
        RECT 268.740 17.040 269.000 17.300 ;
      LAYER met2 ;
        RECT 599.610 510.410 599.890 514.000 ;
        RECT 598.160 510.270 599.890 510.410 ;
        RECT 598.160 449.210 598.300 510.270 ;
        RECT 599.610 510.000 599.890 510.270 ;
        RECT 597.700 449.070 598.300 449.210 ;
        RECT 597.700 448.790 597.840 449.070 ;
        RECT 593.960 448.470 594.220 448.790 ;
        RECT 597.640 448.470 597.900 448.790 ;
        RECT 594.020 424.310 594.160 448.470 ;
        RECT 268.740 423.990 269.000 424.310 ;
        RECT 593.960 423.990 594.220 424.310 ;
        RECT 268.800 17.330 268.940 423.990 ;
        RECT 264.140 17.010 264.400 17.330 ;
        RECT 268.740 17.010 269.000 17.330 ;
        RECT 264.200 2.400 264.340 17.010 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 608.265 193.205 608.435 241.315 ;
      LAYER mcon ;
        RECT 608.265 241.145 608.435 241.315 ;
      LAYER met1 ;
        RECT 607.270 255.240 607.590 255.300 ;
        RECT 608.190 255.240 608.510 255.300 ;
        RECT 607.270 255.100 608.510 255.240 ;
        RECT 607.270 255.040 607.590 255.100 ;
        RECT 608.190 255.040 608.510 255.100 ;
        RECT 608.190 241.300 608.510 241.360 ;
        RECT 607.995 241.160 608.510 241.300 ;
        RECT 608.190 241.100 608.510 241.160 ;
        RECT 608.205 193.360 608.495 193.405 ;
        RECT 608.650 193.360 608.970 193.420 ;
        RECT 608.205 193.220 608.970 193.360 ;
        RECT 608.205 193.175 608.495 193.220 ;
        RECT 608.650 193.160 608.970 193.220 ;
        RECT 282.050 155.280 282.370 155.340 ;
        RECT 608.650 155.280 608.970 155.340 ;
        RECT 282.050 155.140 608.970 155.280 ;
        RECT 282.050 155.080 282.370 155.140 ;
        RECT 608.650 155.080 608.970 155.140 ;
      LAYER via ;
        RECT 607.300 255.040 607.560 255.300 ;
        RECT 608.220 255.040 608.480 255.300 ;
        RECT 608.220 241.100 608.480 241.360 ;
        RECT 608.680 193.160 608.940 193.420 ;
        RECT 282.080 155.080 282.340 155.340 ;
        RECT 608.680 155.080 608.940 155.340 ;
      LAYER met2 ;
        RECT 612.490 510.410 612.770 514.000 ;
        RECT 608.740 510.270 612.770 510.410 ;
        RECT 608.740 449.210 608.880 510.270 ;
        RECT 612.490 510.000 612.770 510.270 ;
        RECT 608.280 449.070 608.880 449.210 ;
        RECT 608.280 351.970 608.420 449.070 ;
        RECT 607.360 351.830 608.420 351.970 ;
        RECT 607.360 351.290 607.500 351.830 ;
        RECT 607.360 351.150 607.960 351.290 ;
        RECT 607.820 255.410 607.960 351.150 ;
        RECT 607.360 255.330 607.960 255.410 ;
        RECT 607.300 255.270 607.960 255.330 ;
        RECT 607.300 255.010 607.560 255.270 ;
        RECT 608.220 255.010 608.480 255.330 ;
        RECT 607.360 254.855 607.500 255.010 ;
        RECT 608.280 241.390 608.420 255.010 ;
        RECT 608.220 241.070 608.480 241.390 ;
        RECT 608.680 193.130 608.940 193.450 ;
        RECT 608.740 155.370 608.880 193.130 ;
        RECT 282.080 155.050 282.340 155.370 ;
        RECT 608.680 155.050 608.940 155.370 ;
        RECT 282.140 2.400 282.280 155.050 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 621.145 386.325 621.315 434.775 ;
        RECT 622.065 289.765 622.235 304.215 ;
        RECT 621.605 241.485 621.775 255.595 ;
      LAYER mcon ;
        RECT 621.145 434.605 621.315 434.775 ;
        RECT 622.065 304.045 622.235 304.215 ;
        RECT 621.605 255.425 621.775 255.595 ;
      LAYER met1 ;
        RECT 621.085 434.760 621.375 434.805 ;
        RECT 621.530 434.760 621.850 434.820 ;
        RECT 621.085 434.620 621.850 434.760 ;
        RECT 621.085 434.575 621.375 434.620 ;
        RECT 621.530 434.560 621.850 434.620 ;
        RECT 621.070 386.480 621.390 386.540 ;
        RECT 620.875 386.340 621.390 386.480 ;
        RECT 621.070 386.280 621.390 386.340 ;
        RECT 621.070 351.800 621.390 351.860 ;
        RECT 621.990 351.800 622.310 351.860 ;
        RECT 621.070 351.660 622.310 351.800 ;
        RECT 621.070 351.600 621.390 351.660 ;
        RECT 621.990 351.600 622.310 351.660 ;
        RECT 621.990 304.200 622.310 304.260 ;
        RECT 621.795 304.060 622.310 304.200 ;
        RECT 621.990 304.000 622.310 304.060 ;
        RECT 621.530 289.920 621.850 289.980 ;
        RECT 622.005 289.920 622.295 289.965 ;
        RECT 621.530 289.780 622.295 289.920 ;
        RECT 621.530 289.720 621.850 289.780 ;
        RECT 622.005 289.735 622.295 289.780 ;
        RECT 621.530 255.580 621.850 255.640 ;
        RECT 621.335 255.440 621.850 255.580 ;
        RECT 621.530 255.380 621.850 255.440 ;
        RECT 621.530 241.640 621.850 241.700 ;
        RECT 621.335 241.500 621.850 241.640 ;
        RECT 621.530 241.440 621.850 241.500 ;
        RECT 303.210 162.080 303.530 162.140 ;
        RECT 621.070 162.080 621.390 162.140 ;
        RECT 303.210 161.940 621.390 162.080 ;
        RECT 303.210 161.880 303.530 161.940 ;
        RECT 621.070 161.880 621.390 161.940 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 621.560 434.560 621.820 434.820 ;
        RECT 621.100 386.280 621.360 386.540 ;
        RECT 621.100 351.600 621.360 351.860 ;
        RECT 622.020 351.600 622.280 351.860 ;
        RECT 622.020 304.000 622.280 304.260 ;
        RECT 621.560 289.720 621.820 289.980 ;
        RECT 621.560 255.380 621.820 255.640 ;
        RECT 621.560 241.440 621.820 241.700 ;
        RECT 303.240 161.880 303.500 162.140 ;
        RECT 621.100 161.880 621.360 162.140 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 624.910 510.340 625.190 514.000 ;
        RECT 624.840 510.000 625.190 510.340 ;
        RECT 624.840 483.325 624.980 510.000 ;
        RECT 622.010 482.955 622.290 483.325 ;
        RECT 624.770 482.955 625.050 483.325 ;
        RECT 622.080 448.530 622.220 482.955 ;
        RECT 621.620 448.390 622.220 448.530 ;
        RECT 621.620 434.850 621.760 448.390 ;
        RECT 621.560 434.530 621.820 434.850 ;
        RECT 621.100 386.250 621.360 386.570 ;
        RECT 621.160 351.890 621.300 386.250 ;
        RECT 621.100 351.570 621.360 351.890 ;
        RECT 622.020 351.570 622.280 351.890 ;
        RECT 622.080 304.290 622.220 351.570 ;
        RECT 622.020 303.970 622.280 304.290 ;
        RECT 621.560 289.690 621.820 290.010 ;
        RECT 621.620 255.670 621.760 289.690 ;
        RECT 621.560 255.350 621.820 255.670 ;
        RECT 621.560 241.410 621.820 241.730 ;
        RECT 621.620 241.130 621.760 241.410 ;
        RECT 621.160 240.990 621.760 241.130 ;
        RECT 621.160 162.170 621.300 240.990 ;
        RECT 303.240 161.850 303.500 162.170 ;
        RECT 621.100 161.850 621.360 162.170 ;
        RECT 303.300 16.990 303.440 161.850 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 622.010 483.000 622.290 483.280 ;
        RECT 624.770 483.000 625.050 483.280 ;
      LAYER met3 ;
        RECT 621.985 483.290 622.315 483.305 ;
        RECT 624.745 483.290 625.075 483.305 ;
        RECT 621.985 482.990 625.075 483.290 ;
        RECT 621.985 482.975 622.315 482.990 ;
        RECT 624.745 482.975 625.075 482.990 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 417.420 324.230 417.480 ;
        RECT 634.870 417.420 635.190 417.480 ;
        RECT 323.910 417.280 635.190 417.420 ;
        RECT 323.910 417.220 324.230 417.280 ;
        RECT 634.870 417.220 635.190 417.280 ;
        RECT 317.930 16.560 318.250 16.620 ;
        RECT 323.910 16.560 324.230 16.620 ;
        RECT 317.930 16.420 324.230 16.560 ;
        RECT 317.930 16.360 318.250 16.420 ;
        RECT 323.910 16.360 324.230 16.420 ;
      LAYER via ;
        RECT 323.940 417.220 324.200 417.480 ;
        RECT 634.900 417.220 635.160 417.480 ;
        RECT 317.960 16.360 318.220 16.620 ;
        RECT 323.940 16.360 324.200 16.620 ;
      LAYER met2 ;
        RECT 637.790 510.410 638.070 514.000 ;
        RECT 634.960 510.270 638.070 510.410 ;
        RECT 634.960 417.510 635.100 510.270 ;
        RECT 637.790 510.000 638.070 510.270 ;
        RECT 323.940 417.190 324.200 417.510 ;
        RECT 634.900 417.190 635.160 417.510 ;
        RECT 324.000 16.650 324.140 417.190 ;
        RECT 317.960 16.330 318.220 16.650 ;
        RECT 323.940 16.330 324.200 16.650 ;
        RECT 318.020 2.400 318.160 16.330 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 496.980 645.310 497.040 ;
        RECT 650.510 496.980 650.830 497.040 ;
        RECT 644.990 496.840 650.830 496.980 ;
        RECT 644.990 496.780 645.310 496.840 ;
        RECT 650.510 496.780 650.830 496.840 ;
        RECT 337.710 410.620 338.030 410.680 ;
        RECT 644.990 410.620 645.310 410.680 ;
        RECT 337.710 410.480 645.310 410.620 ;
        RECT 337.710 410.420 338.030 410.480 ;
        RECT 644.990 410.420 645.310 410.480 ;
      LAYER via ;
        RECT 645.020 496.780 645.280 497.040 ;
        RECT 650.540 496.780 650.800 497.040 ;
        RECT 337.740 410.420 338.000 410.680 ;
        RECT 645.020 410.420 645.280 410.680 ;
      LAYER met2 ;
        RECT 650.670 510.340 650.950 514.000 ;
        RECT 650.600 510.000 650.950 510.340 ;
        RECT 650.600 497.070 650.740 510.000 ;
        RECT 645.020 496.750 645.280 497.070 ;
        RECT 650.540 496.750 650.800 497.070 ;
        RECT 645.080 410.710 645.220 496.750 ;
        RECT 337.740 410.390 338.000 410.710 ;
        RECT 645.020 410.390 645.280 410.710 ;
        RECT 337.800 17.410 337.940 410.390 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 403.480 358.730 403.540 ;
        RECT 662.930 403.480 663.250 403.540 ;
        RECT 358.410 403.340 663.250 403.480 ;
        RECT 358.410 403.280 358.730 403.340 ;
        RECT 662.930 403.280 663.250 403.340 ;
        RECT 353.350 17.240 353.670 17.300 ;
        RECT 358.410 17.240 358.730 17.300 ;
        RECT 353.350 17.100 358.730 17.240 ;
        RECT 353.350 17.040 353.670 17.100 ;
        RECT 358.410 17.040 358.730 17.100 ;
      LAYER via ;
        RECT 358.440 403.280 358.700 403.540 ;
        RECT 662.960 403.280 663.220 403.540 ;
        RECT 353.380 17.040 353.640 17.300 ;
        RECT 358.440 17.040 358.700 17.300 ;
      LAYER met2 ;
        RECT 663.550 510.410 663.830 514.000 ;
        RECT 663.020 510.270 663.830 510.410 ;
        RECT 663.020 403.570 663.160 510.270 ;
        RECT 663.550 510.000 663.830 510.270 ;
        RECT 358.440 403.250 358.700 403.570 ;
        RECT 662.960 403.250 663.220 403.570 ;
        RECT 358.500 17.330 358.640 403.250 ;
        RECT 353.380 17.010 353.640 17.330 ;
        RECT 358.440 17.010 358.700 17.330 ;
        RECT 353.440 2.400 353.580 17.010 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 389.880 372.530 389.940 ;
        RECT 676.730 389.880 677.050 389.940 ;
        RECT 372.210 389.740 677.050 389.880 ;
        RECT 372.210 389.680 372.530 389.740 ;
        RECT 676.730 389.680 677.050 389.740 ;
      LAYER via ;
        RECT 372.240 389.680 372.500 389.940 ;
        RECT 676.760 389.680 677.020 389.940 ;
      LAYER met2 ;
        RECT 676.430 510.340 676.710 514.000 ;
        RECT 676.360 510.000 676.710 510.340 ;
        RECT 676.360 473.690 676.500 510.000 ;
        RECT 676.360 473.550 676.960 473.690 ;
        RECT 676.820 389.970 676.960 473.550 ;
        RECT 372.240 389.650 372.500 389.970 ;
        RECT 676.760 389.650 677.020 389.970 ;
        RECT 372.300 17.410 372.440 389.650 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 683.705 338.045 683.875 386.155 ;
        RECT 684.165 241.485 684.335 289.595 ;
      LAYER mcon ;
        RECT 683.705 385.985 683.875 386.155 ;
        RECT 684.165 289.425 684.335 289.595 ;
      LAYER met1 ;
        RECT 683.630 386.140 683.950 386.200 ;
        RECT 683.435 386.000 683.950 386.140 ;
        RECT 683.630 385.940 683.950 386.000 ;
        RECT 683.645 338.200 683.935 338.245 ;
        RECT 684.090 338.200 684.410 338.260 ;
        RECT 683.645 338.060 684.410 338.200 ;
        RECT 683.645 338.015 683.935 338.060 ;
        RECT 684.090 338.000 684.410 338.060 ;
        RECT 684.105 289.580 684.395 289.625 ;
        RECT 684.550 289.580 684.870 289.640 ;
        RECT 684.105 289.440 684.870 289.580 ;
        RECT 684.105 289.395 684.395 289.440 ;
        RECT 684.550 289.380 684.870 289.440 ;
        RECT 684.090 241.640 684.410 241.700 ;
        RECT 683.895 241.500 684.410 241.640 ;
        RECT 684.090 241.440 684.410 241.500 ;
        RECT 392.910 168.880 393.230 168.940 ;
        RECT 684.550 168.880 684.870 168.940 ;
        RECT 392.910 168.740 684.870 168.880 ;
        RECT 392.910 168.680 393.230 168.740 ;
        RECT 684.550 168.680 684.870 168.740 ;
        RECT 389.230 17.580 389.550 17.640 ;
        RECT 392.910 17.580 393.230 17.640 ;
        RECT 389.230 17.440 393.230 17.580 ;
        RECT 389.230 17.380 389.550 17.440 ;
        RECT 392.910 17.380 393.230 17.440 ;
      LAYER via ;
        RECT 683.660 385.940 683.920 386.200 ;
        RECT 684.120 338.000 684.380 338.260 ;
        RECT 684.580 289.380 684.840 289.640 ;
        RECT 684.120 241.440 684.380 241.700 ;
        RECT 392.940 168.680 393.200 168.940 ;
        RECT 684.580 168.680 684.840 168.940 ;
        RECT 389.260 17.380 389.520 17.640 ;
        RECT 392.940 17.380 393.200 17.640 ;
      LAYER met2 ;
        RECT 689.310 510.410 689.590 514.000 ;
        RECT 686.480 510.270 689.590 510.410 ;
        RECT 686.480 449.210 686.620 510.270 ;
        RECT 689.310 510.000 689.590 510.270 ;
        RECT 685.560 449.070 686.620 449.210 ;
        RECT 685.560 448.530 685.700 449.070 ;
        RECT 684.180 448.390 685.700 448.530 ;
        RECT 684.180 400.930 684.320 448.390 ;
        RECT 684.180 400.790 684.780 400.930 ;
        RECT 684.640 387.330 684.780 400.790 ;
        RECT 684.180 387.190 684.780 387.330 ;
        RECT 684.180 386.650 684.320 387.190 ;
        RECT 683.720 386.510 684.320 386.650 ;
        RECT 683.720 386.230 683.860 386.510 ;
        RECT 683.660 385.910 683.920 386.230 ;
        RECT 684.120 337.970 684.380 338.290 ;
        RECT 684.180 303.690 684.320 337.970 ;
        RECT 684.180 303.550 684.780 303.690 ;
        RECT 684.640 289.670 684.780 303.550 ;
        RECT 684.580 289.350 684.840 289.670 ;
        RECT 684.120 241.410 684.380 241.730 ;
        RECT 684.180 207.130 684.320 241.410 ;
        RECT 684.180 206.990 684.780 207.130 ;
        RECT 684.640 168.970 684.780 206.990 ;
        RECT 392.940 168.650 393.200 168.970 ;
        RECT 684.580 168.650 684.840 168.970 ;
        RECT 393.000 17.670 393.140 168.650 ;
        RECT 389.260 17.350 389.520 17.670 ;
        RECT 392.940 17.350 393.200 17.670 ;
        RECT 389.320 2.400 389.460 17.350 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 472.840 697.290 472.900 ;
        RECT 700.190 472.840 700.510 472.900 ;
        RECT 696.970 472.700 700.510 472.840 ;
        RECT 696.970 472.640 697.290 472.700 ;
        RECT 700.190 472.640 700.510 472.700 ;
        RECT 413.150 176.020 413.470 176.080 ;
        RECT 696.970 176.020 697.290 176.080 ;
        RECT 413.150 175.880 697.290 176.020 ;
        RECT 413.150 175.820 413.470 175.880 ;
        RECT 696.970 175.820 697.290 175.880 ;
        RECT 407.170 17.580 407.490 17.640 ;
        RECT 413.150 17.580 413.470 17.640 ;
        RECT 407.170 17.440 413.470 17.580 ;
        RECT 407.170 17.380 407.490 17.440 ;
        RECT 413.150 17.380 413.470 17.440 ;
      LAYER via ;
        RECT 697.000 472.640 697.260 472.900 ;
        RECT 700.220 472.640 700.480 472.900 ;
        RECT 413.180 175.820 413.440 176.080 ;
        RECT 697.000 175.820 697.260 176.080 ;
        RECT 407.200 17.380 407.460 17.640 ;
        RECT 413.180 17.380 413.440 17.640 ;
      LAYER met2 ;
        RECT 701.730 510.410 702.010 514.000 ;
        RECT 700.280 510.270 702.010 510.410 ;
        RECT 700.280 472.930 700.420 510.270 ;
        RECT 701.730 510.000 702.010 510.270 ;
        RECT 697.000 472.610 697.260 472.930 ;
        RECT 700.220 472.610 700.480 472.930 ;
        RECT 697.060 176.110 697.200 472.610 ;
        RECT 413.180 175.790 413.440 176.110 ;
        RECT 697.000 175.790 697.260 176.110 ;
        RECT 413.240 17.670 413.380 175.790 ;
        RECT 407.200 17.350 407.460 17.670 ;
        RECT 413.180 17.350 413.440 17.670 ;
        RECT 407.260 2.400 407.400 17.350 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 93.060 68.470 93.120 ;
        RECT 455.470 93.060 455.790 93.120 ;
        RECT 68.150 92.920 455.790 93.060 ;
        RECT 68.150 92.860 68.470 92.920 ;
        RECT 455.470 92.860 455.790 92.920 ;
      LAYER via ;
        RECT 68.180 92.860 68.440 93.120 ;
        RECT 455.500 92.860 455.760 93.120 ;
      LAYER met2 ;
        RECT 458.850 510.410 459.130 514.000 ;
        RECT 455.560 510.270 459.130 510.410 ;
        RECT 455.560 93.150 455.700 510.270 ;
        RECT 458.850 510.000 459.130 510.270 ;
        RECT 68.180 92.830 68.440 93.150 ;
        RECT 455.500 92.830 455.760 93.150 ;
        RECT 68.240 2.400 68.380 92.830 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 710.845 386.325 711.015 434.775 ;
        RECT 710.845 351.645 711.015 385.815 ;
      LAYER mcon ;
        RECT 710.845 434.605 711.015 434.775 ;
        RECT 710.845 385.645 711.015 385.815 ;
      LAYER met1 ;
        RECT 710.785 434.760 711.075 434.805 ;
        RECT 711.230 434.760 711.550 434.820 ;
        RECT 710.785 434.620 711.550 434.760 ;
        RECT 710.785 434.575 711.075 434.620 ;
        RECT 711.230 434.560 711.550 434.620 ;
        RECT 710.770 386.480 711.090 386.540 ;
        RECT 710.575 386.340 711.090 386.480 ;
        RECT 710.770 386.280 711.090 386.340 ;
        RECT 710.770 385.800 711.090 385.860 ;
        RECT 710.575 385.660 711.090 385.800 ;
        RECT 710.770 385.600 711.090 385.660 ;
        RECT 710.785 351.800 711.075 351.845 ;
        RECT 711.230 351.800 711.550 351.860 ;
        RECT 710.785 351.660 711.550 351.800 ;
        RECT 710.785 351.615 711.075 351.660 ;
        RECT 711.230 351.600 711.550 351.660 ;
        RECT 427.410 210.360 427.730 210.420 ;
        RECT 711.690 210.360 712.010 210.420 ;
        RECT 427.410 210.220 712.010 210.360 ;
        RECT 427.410 210.160 427.730 210.220 ;
        RECT 711.690 210.160 712.010 210.220 ;
        RECT 424.650 17.580 424.970 17.640 ;
        RECT 427.410 17.580 427.730 17.640 ;
        RECT 424.650 17.440 427.730 17.580 ;
        RECT 424.650 17.380 424.970 17.440 ;
        RECT 427.410 17.380 427.730 17.440 ;
      LAYER via ;
        RECT 711.260 434.560 711.520 434.820 ;
        RECT 710.800 386.280 711.060 386.540 ;
        RECT 710.800 385.600 711.060 385.860 ;
        RECT 711.260 351.600 711.520 351.860 ;
        RECT 427.440 210.160 427.700 210.420 ;
        RECT 711.720 210.160 711.980 210.420 ;
        RECT 424.680 17.380 424.940 17.640 ;
        RECT 427.440 17.380 427.700 17.640 ;
      LAYER met2 ;
        RECT 714.610 510.340 714.890 514.000 ;
        RECT 714.540 510.000 714.890 510.340 ;
        RECT 714.540 483.325 714.680 510.000 ;
        RECT 711.710 482.955 711.990 483.325 ;
        RECT 714.470 482.955 714.750 483.325 ;
        RECT 711.780 448.530 711.920 482.955 ;
        RECT 711.320 448.390 711.920 448.530 ;
        RECT 711.320 434.850 711.460 448.390 ;
        RECT 711.260 434.530 711.520 434.850 ;
        RECT 710.800 386.250 711.060 386.570 ;
        RECT 710.860 385.890 711.000 386.250 ;
        RECT 710.800 385.570 711.060 385.890 ;
        RECT 711.260 351.570 711.520 351.890 ;
        RECT 711.320 255.410 711.460 351.570 ;
        RECT 711.320 255.270 711.920 255.410 ;
        RECT 711.780 210.450 711.920 255.270 ;
        RECT 427.440 210.130 427.700 210.450 ;
        RECT 711.720 210.130 711.980 210.450 ;
        RECT 427.500 17.670 427.640 210.130 ;
        RECT 424.680 17.350 424.940 17.670 ;
        RECT 427.440 17.350 427.700 17.670 ;
        RECT 424.740 2.400 424.880 17.350 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 711.710 483.000 711.990 483.280 ;
        RECT 714.470 483.000 714.750 483.280 ;
      LAYER met3 ;
        RECT 711.685 483.290 712.015 483.305 ;
        RECT 714.445 483.290 714.775 483.305 ;
        RECT 711.685 482.990 714.775 483.290 ;
        RECT 711.685 482.975 712.015 482.990 ;
        RECT 714.445 482.975 714.775 482.990 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 224.300 448.430 224.360 ;
        RECT 724.570 224.300 724.890 224.360 ;
        RECT 448.110 224.160 724.890 224.300 ;
        RECT 448.110 224.100 448.430 224.160 ;
        RECT 724.570 224.100 724.890 224.160 ;
        RECT 442.590 17.580 442.910 17.640 ;
        RECT 448.110 17.580 448.430 17.640 ;
        RECT 442.590 17.440 448.430 17.580 ;
        RECT 442.590 17.380 442.910 17.440 ;
        RECT 448.110 17.380 448.430 17.440 ;
      LAYER via ;
        RECT 448.140 224.100 448.400 224.360 ;
        RECT 724.600 224.100 724.860 224.360 ;
        RECT 442.620 17.380 442.880 17.640 ;
        RECT 448.140 17.380 448.400 17.640 ;
      LAYER met2 ;
        RECT 727.490 510.410 727.770 514.000 ;
        RECT 724.660 510.270 727.770 510.410 ;
        RECT 724.660 224.390 724.800 510.270 ;
        RECT 727.490 510.000 727.770 510.270 ;
        RECT 448.140 224.070 448.400 224.390 ;
        RECT 724.600 224.070 724.860 224.390 ;
        RECT 448.200 17.670 448.340 224.070 ;
        RECT 442.620 17.350 442.880 17.670 ;
        RECT 448.140 17.350 448.400 17.670 ;
        RECT 442.680 2.400 442.820 17.350 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 396.680 462.230 396.740 ;
        RECT 738.830 396.680 739.150 396.740 ;
        RECT 461.910 396.540 739.150 396.680 ;
        RECT 461.910 396.480 462.230 396.540 ;
        RECT 738.830 396.480 739.150 396.540 ;
      LAYER via ;
        RECT 461.940 396.480 462.200 396.740 ;
        RECT 738.860 396.480 739.120 396.740 ;
      LAYER met2 ;
        RECT 740.370 510.410 740.650 514.000 ;
        RECT 738.920 510.270 740.650 510.410 ;
        RECT 738.920 396.770 739.060 510.270 ;
        RECT 740.370 510.000 740.650 510.270 ;
        RECT 461.940 396.450 462.200 396.770 ;
        RECT 738.860 396.450 739.120 396.770 ;
        RECT 462.000 16.730 462.140 396.450 ;
        RECT 460.620 16.590 462.140 16.730 ;
        RECT 460.620 2.400 460.760 16.590 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 231.100 482.930 231.160 ;
        RECT 752.630 231.100 752.950 231.160 ;
        RECT 482.610 230.960 752.950 231.100 ;
        RECT 482.610 230.900 482.930 230.960 ;
        RECT 752.630 230.900 752.950 230.960 ;
        RECT 478.470 17.580 478.790 17.640 ;
        RECT 482.610 17.580 482.930 17.640 ;
        RECT 478.470 17.440 482.930 17.580 ;
        RECT 478.470 17.380 478.790 17.440 ;
        RECT 482.610 17.380 482.930 17.440 ;
      LAYER via ;
        RECT 482.640 230.900 482.900 231.160 ;
        RECT 752.660 230.900 752.920 231.160 ;
        RECT 478.500 17.380 478.760 17.640 ;
        RECT 482.640 17.380 482.900 17.640 ;
      LAYER met2 ;
        RECT 753.250 510.410 753.530 514.000 ;
        RECT 752.720 510.270 753.530 510.410 ;
        RECT 752.720 231.190 752.860 510.270 ;
        RECT 753.250 510.000 753.530 510.270 ;
        RECT 482.640 230.870 482.900 231.190 ;
        RECT 752.660 230.870 752.920 231.190 ;
        RECT 482.700 17.670 482.840 230.870 ;
        RECT 478.500 17.350 478.760 17.670 ;
        RECT 482.640 17.350 482.900 17.670 ;
        RECT 478.560 2.400 478.700 17.350 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 500.380 624.610 500.440 ;
        RECT 765.970 500.380 766.290 500.440 ;
        RECT 624.290 500.240 766.290 500.380 ;
        RECT 624.290 500.180 624.610 500.240 ;
        RECT 765.970 500.180 766.290 500.240 ;
        RECT 496.410 24.040 496.730 24.100 ;
        RECT 624.290 24.040 624.610 24.100 ;
        RECT 496.410 23.900 624.610 24.040 ;
        RECT 496.410 23.840 496.730 23.900 ;
        RECT 624.290 23.840 624.610 23.900 ;
      LAYER via ;
        RECT 624.320 500.180 624.580 500.440 ;
        RECT 766.000 500.180 766.260 500.440 ;
        RECT 496.440 23.840 496.700 24.100 ;
        RECT 624.320 23.840 624.580 24.100 ;
      LAYER met2 ;
        RECT 766.130 510.340 766.410 514.000 ;
        RECT 766.060 510.000 766.410 510.340 ;
        RECT 766.060 500.470 766.200 510.000 ;
        RECT 624.320 500.150 624.580 500.470 ;
        RECT 766.000 500.150 766.260 500.470 ;
        RECT 624.380 24.130 624.520 500.150 ;
        RECT 496.440 23.810 496.700 24.130 ;
        RECT 624.320 23.810 624.580 24.130 ;
        RECT 496.500 2.400 496.640 23.810 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 773.865 338.045 774.035 403.835 ;
      LAYER mcon ;
        RECT 773.865 403.665 774.035 403.835 ;
      LAYER met1 ;
        RECT 773.805 403.820 774.095 403.865 ;
        RECT 774.710 403.820 775.030 403.880 ;
        RECT 773.805 403.680 775.030 403.820 ;
        RECT 773.805 403.635 774.095 403.680 ;
        RECT 774.710 403.620 775.030 403.680 ;
        RECT 773.790 338.200 774.110 338.260 ;
        RECT 773.595 338.060 774.110 338.200 ;
        RECT 773.790 338.000 774.110 338.060 ;
        RECT 517.110 237.900 517.430 237.960 ;
        RECT 773.790 237.900 774.110 237.960 ;
        RECT 517.110 237.760 774.110 237.900 ;
        RECT 517.110 237.700 517.430 237.760 ;
        RECT 773.790 237.700 774.110 237.760 ;
        RECT 513.890 16.560 514.210 16.620 ;
        RECT 517.110 16.560 517.430 16.620 ;
        RECT 513.890 16.420 517.430 16.560 ;
        RECT 513.890 16.360 514.210 16.420 ;
        RECT 517.110 16.360 517.430 16.420 ;
      LAYER via ;
        RECT 774.740 403.620 775.000 403.880 ;
        RECT 773.820 338.000 774.080 338.260 ;
        RECT 517.140 237.700 517.400 237.960 ;
        RECT 773.820 237.700 774.080 237.960 ;
        RECT 513.920 16.360 514.180 16.620 ;
        RECT 517.140 16.360 517.400 16.620 ;
      LAYER met2 ;
        RECT 778.550 510.410 778.830 514.000 ;
        RECT 775.720 510.270 778.830 510.410 ;
        RECT 775.720 449.210 775.860 510.270 ;
        RECT 778.550 510.000 778.830 510.270 ;
        RECT 774.800 449.070 775.860 449.210 ;
        RECT 774.800 403.910 774.940 449.070 ;
        RECT 774.740 403.590 775.000 403.910 ;
        RECT 773.820 337.970 774.080 338.290 ;
        RECT 773.880 237.990 774.020 337.970 ;
        RECT 517.140 237.670 517.400 237.990 ;
        RECT 773.820 237.670 774.080 237.990 ;
        RECT 517.200 16.650 517.340 237.670 ;
        RECT 513.920 16.330 514.180 16.650 ;
        RECT 517.140 16.330 517.400 16.650 ;
        RECT 513.980 2.400 514.120 16.330 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 787.590 303.860 787.910 303.920 ;
        RECT 786.760 303.720 787.910 303.860 ;
        RECT 786.760 303.580 786.900 303.720 ;
        RECT 787.590 303.660 787.910 303.720 ;
        RECT 786.670 303.320 786.990 303.580 ;
        RECT 537.810 251.840 538.130 251.900 ;
        RECT 786.670 251.840 786.990 251.900 ;
        RECT 537.810 251.700 786.990 251.840 ;
        RECT 537.810 251.640 538.130 251.700 ;
        RECT 786.670 251.640 786.990 251.700 ;
        RECT 531.830 16.900 532.150 16.960 ;
        RECT 537.810 16.900 538.130 16.960 ;
        RECT 531.830 16.760 538.130 16.900 ;
        RECT 531.830 16.700 532.150 16.760 ;
        RECT 537.810 16.700 538.130 16.760 ;
      LAYER via ;
        RECT 787.620 303.660 787.880 303.920 ;
        RECT 786.700 303.320 786.960 303.580 ;
        RECT 537.840 251.640 538.100 251.900 ;
        RECT 786.700 251.640 786.960 251.900 ;
        RECT 531.860 16.700 532.120 16.960 ;
        RECT 537.840 16.700 538.100 16.960 ;
      LAYER met2 ;
        RECT 791.430 510.410 791.710 514.000 ;
        RECT 788.140 510.270 791.710 510.410 ;
        RECT 788.140 449.210 788.280 510.270 ;
        RECT 791.430 510.000 791.710 510.270 ;
        RECT 787.680 449.070 788.280 449.210 ;
        RECT 787.680 303.950 787.820 449.070 ;
        RECT 787.620 303.630 787.880 303.950 ;
        RECT 786.700 303.290 786.960 303.610 ;
        RECT 786.760 251.930 786.900 303.290 ;
        RECT 537.840 251.610 538.100 251.930 ;
        RECT 786.700 251.610 786.960 251.930 ;
        RECT 537.900 16.990 538.040 251.610 ;
        RECT 531.860 16.670 532.120 16.990 ;
        RECT 537.840 16.670 538.100 16.990 ;
        RECT 531.920 2.400 532.060 16.670 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 801.005 379.525 801.175 427.635 ;
        RECT 801.005 289.765 801.175 337.875 ;
      LAYER mcon ;
        RECT 801.005 427.465 801.175 427.635 ;
        RECT 801.005 337.705 801.175 337.875 ;
      LAYER met1 ;
        RECT 800.470 496.980 800.790 497.040 ;
        RECT 804.150 496.980 804.470 497.040 ;
        RECT 800.470 496.840 804.470 496.980 ;
        RECT 800.470 496.780 800.790 496.840 ;
        RECT 804.150 496.780 804.470 496.840 ;
        RECT 800.470 448.500 800.790 448.760 ;
        RECT 800.560 448.020 800.700 448.500 ;
        RECT 800.930 448.020 801.250 448.080 ;
        RECT 800.560 447.880 801.250 448.020 ;
        RECT 800.930 447.820 801.250 447.880 ;
        RECT 800.930 427.620 801.250 427.680 ;
        RECT 800.735 427.480 801.250 427.620 ;
        RECT 800.930 427.420 801.250 427.480 ;
        RECT 800.930 379.680 801.250 379.740 ;
        RECT 800.735 379.540 801.250 379.680 ;
        RECT 800.930 379.480 801.250 379.540 ;
        RECT 800.930 337.860 801.250 337.920 ;
        RECT 800.735 337.720 801.250 337.860 ;
        RECT 800.930 337.660 801.250 337.720 ;
        RECT 800.930 289.920 801.250 289.980 ;
        RECT 800.735 289.780 801.250 289.920 ;
        RECT 800.930 289.720 801.250 289.780 ;
        RECT 551.610 258.640 551.930 258.700 ;
        RECT 800.930 258.640 801.250 258.700 ;
        RECT 551.610 258.500 801.250 258.640 ;
        RECT 551.610 258.440 551.930 258.500 ;
        RECT 800.930 258.440 801.250 258.500 ;
        RECT 549.770 2.960 550.090 3.020 ;
        RECT 551.610 2.960 551.930 3.020 ;
        RECT 549.770 2.820 551.930 2.960 ;
        RECT 549.770 2.760 550.090 2.820 ;
        RECT 551.610 2.760 551.930 2.820 ;
      LAYER via ;
        RECT 800.500 496.780 800.760 497.040 ;
        RECT 804.180 496.780 804.440 497.040 ;
        RECT 800.500 448.500 800.760 448.760 ;
        RECT 800.960 447.820 801.220 448.080 ;
        RECT 800.960 427.420 801.220 427.680 ;
        RECT 800.960 379.480 801.220 379.740 ;
        RECT 800.960 337.660 801.220 337.920 ;
        RECT 800.960 289.720 801.220 289.980 ;
        RECT 551.640 258.440 551.900 258.700 ;
        RECT 800.960 258.440 801.220 258.700 ;
        RECT 549.800 2.760 550.060 3.020 ;
        RECT 551.640 2.760 551.900 3.020 ;
      LAYER met2 ;
        RECT 804.310 510.340 804.590 514.000 ;
        RECT 804.240 510.000 804.590 510.340 ;
        RECT 804.240 497.070 804.380 510.000 ;
        RECT 800.500 496.750 800.760 497.070 ;
        RECT 804.180 496.750 804.440 497.070 ;
        RECT 800.560 448.790 800.700 496.750 ;
        RECT 800.500 448.470 800.760 448.790 ;
        RECT 800.960 447.790 801.220 448.110 ;
        RECT 801.020 427.710 801.160 447.790 ;
        RECT 800.960 427.390 801.220 427.710 ;
        RECT 800.960 379.450 801.220 379.770 ;
        RECT 801.020 337.950 801.160 379.450 ;
        RECT 800.960 337.630 801.220 337.950 ;
        RECT 800.960 289.690 801.220 290.010 ;
        RECT 801.020 258.730 801.160 289.690 ;
        RECT 551.640 258.410 551.900 258.730 ;
        RECT 800.960 258.410 801.220 258.730 ;
        RECT 551.700 3.050 551.840 258.410 ;
        RECT 549.800 2.730 550.060 3.050 ;
        RECT 551.640 2.730 551.900 3.050 ;
        RECT 549.860 2.400 550.000 2.730 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 265.440 572.630 265.500 ;
        RECT 814.270 265.440 814.590 265.500 ;
        RECT 572.310 265.300 814.590 265.440 ;
        RECT 572.310 265.240 572.630 265.300 ;
        RECT 814.270 265.240 814.590 265.300 ;
        RECT 567.710 20.640 568.030 20.700 ;
        RECT 572.310 20.640 572.630 20.700 ;
        RECT 567.710 20.500 572.630 20.640 ;
        RECT 567.710 20.440 568.030 20.500 ;
        RECT 572.310 20.440 572.630 20.500 ;
      LAYER via ;
        RECT 572.340 265.240 572.600 265.500 ;
        RECT 814.300 265.240 814.560 265.500 ;
        RECT 567.740 20.440 568.000 20.700 ;
        RECT 572.340 20.440 572.600 20.700 ;
      LAYER met2 ;
        RECT 817.190 510.410 817.470 514.000 ;
        RECT 814.360 510.270 817.470 510.410 ;
        RECT 814.360 265.530 814.500 510.270 ;
        RECT 817.190 510.000 817.470 510.270 ;
        RECT 572.340 265.210 572.600 265.530 ;
        RECT 814.300 265.210 814.560 265.530 ;
        RECT 572.400 20.730 572.540 265.210 ;
        RECT 567.740 20.410 568.000 20.730 ;
        RECT 572.340 20.410 572.600 20.730 ;
        RECT 567.800 2.400 567.940 20.410 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 789.890 503.440 790.210 503.500 ;
        RECT 829.910 503.440 830.230 503.500 ;
        RECT 789.890 503.300 830.230 503.440 ;
        RECT 789.890 503.240 790.210 503.300 ;
        RECT 829.910 503.240 830.230 503.300 ;
        RECT 585.650 72.660 585.970 72.720 ;
        RECT 789.890 72.660 790.210 72.720 ;
        RECT 585.650 72.520 790.210 72.660 ;
        RECT 585.650 72.460 585.970 72.520 ;
        RECT 789.890 72.460 790.210 72.520 ;
      LAYER via ;
        RECT 789.920 503.240 790.180 503.500 ;
        RECT 829.940 503.240 830.200 503.500 ;
        RECT 585.680 72.460 585.940 72.720 ;
        RECT 789.920 72.460 790.180 72.720 ;
      LAYER met2 ;
        RECT 830.070 510.340 830.350 514.000 ;
        RECT 830.000 510.000 830.350 510.340 ;
        RECT 830.000 503.530 830.140 510.000 ;
        RECT 789.920 503.210 790.180 503.530 ;
        RECT 829.940 503.210 830.200 503.530 ;
        RECT 789.980 72.750 790.120 503.210 ;
        RECT 585.680 72.430 585.940 72.750 ;
        RECT 789.920 72.430 790.180 72.750 ;
        RECT 585.740 2.400 585.880 72.430 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 469.730 241.640 470.050 241.700 ;
        RECT 470.190 241.640 470.510 241.700 ;
        RECT 469.730 241.500 470.510 241.640 ;
        RECT 469.730 241.440 470.050 241.500 ;
        RECT 470.190 241.440 470.510 241.500 ;
        RECT 96.210 99.860 96.530 99.920 ;
        RECT 470.650 99.860 470.970 99.920 ;
        RECT 96.210 99.720 470.970 99.860 ;
        RECT 96.210 99.660 96.530 99.720 ;
        RECT 470.650 99.660 470.970 99.720 ;
        RECT 91.610 20.640 91.930 20.700 ;
        RECT 96.210 20.640 96.530 20.700 ;
        RECT 91.610 20.500 96.530 20.640 ;
        RECT 91.610 20.440 91.930 20.500 ;
        RECT 96.210 20.440 96.530 20.500 ;
      LAYER via ;
        RECT 469.760 241.440 470.020 241.700 ;
        RECT 470.220 241.440 470.480 241.700 ;
        RECT 96.240 99.660 96.500 99.920 ;
        RECT 470.680 99.660 470.940 99.920 ;
        RECT 91.640 20.440 91.900 20.700 ;
        RECT 96.240 20.440 96.500 20.700 ;
      LAYER met2 ;
        RECT 475.870 510.410 476.150 514.000 ;
        RECT 472.580 510.270 476.150 510.410 ;
        RECT 472.580 472.330 472.720 510.270 ;
        RECT 475.870 510.000 476.150 510.270 ;
        RECT 469.820 472.190 472.720 472.330 ;
        RECT 469.820 400.930 469.960 472.190 ;
        RECT 469.360 400.790 469.960 400.930 ;
        RECT 469.360 400.250 469.500 400.790 ;
        RECT 469.360 400.110 469.960 400.250 ;
        RECT 469.820 399.570 469.960 400.110 ;
        RECT 469.820 399.430 470.420 399.570 ;
        RECT 470.280 241.730 470.420 399.430 ;
        RECT 469.760 241.410 470.020 241.730 ;
        RECT 470.220 241.410 470.480 241.730 ;
        RECT 469.820 207.130 469.960 241.410 ;
        RECT 469.820 206.990 470.420 207.130 ;
        RECT 470.280 158.850 470.420 206.990 ;
        RECT 470.280 158.710 470.880 158.850 ;
        RECT 470.740 99.950 470.880 158.710 ;
        RECT 96.240 99.630 96.500 99.950 ;
        RECT 470.680 99.630 470.940 99.950 ;
        RECT 96.300 20.730 96.440 99.630 ;
        RECT 91.640 20.410 91.900 20.730 ;
        RECT 96.240 20.410 96.500 20.730 ;
        RECT 91.700 2.400 91.840 20.410 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 272.580 607.130 272.640 ;
        RECT 842.330 272.580 842.650 272.640 ;
        RECT 606.810 272.440 842.650 272.580 ;
        RECT 606.810 272.380 607.130 272.440 ;
        RECT 842.330 272.380 842.650 272.440 ;
        RECT 603.130 16.900 603.450 16.960 ;
        RECT 606.810 16.900 607.130 16.960 ;
        RECT 603.130 16.760 607.130 16.900 ;
        RECT 603.130 16.700 603.450 16.760 ;
        RECT 606.810 16.700 607.130 16.760 ;
      LAYER via ;
        RECT 606.840 272.380 607.100 272.640 ;
        RECT 842.360 272.380 842.620 272.640 ;
        RECT 603.160 16.700 603.420 16.960 ;
        RECT 606.840 16.700 607.100 16.960 ;
      LAYER met2 ;
        RECT 842.950 510.410 843.230 514.000 ;
        RECT 842.420 510.270 843.230 510.410 ;
        RECT 842.420 272.670 842.560 510.270 ;
        RECT 842.950 510.000 843.230 510.270 ;
        RECT 606.840 272.350 607.100 272.670 ;
        RECT 842.360 272.350 842.620 272.670 ;
        RECT 606.900 16.990 607.040 272.350 ;
        RECT 603.160 16.670 603.420 16.990 ;
        RECT 606.840 16.670 607.100 16.990 ;
        RECT 603.220 2.400 603.360 16.670 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 849.765 379.525 849.935 427.635 ;
      LAYER mcon ;
        RECT 849.765 427.465 849.935 427.635 ;
      LAYER met1 ;
        RECT 849.690 448.700 850.010 448.760 ;
        RECT 851.990 448.700 852.310 448.760 ;
        RECT 849.690 448.560 852.310 448.700 ;
        RECT 849.690 448.500 850.010 448.560 ;
        RECT 851.990 448.500 852.310 448.560 ;
        RECT 849.690 427.620 850.010 427.680 ;
        RECT 849.495 427.480 850.010 427.620 ;
        RECT 849.690 427.420 850.010 427.480 ;
        RECT 849.690 379.680 850.010 379.740 ;
        RECT 849.495 379.540 850.010 379.680 ;
        RECT 849.690 379.480 850.010 379.540 ;
        RECT 849.690 351.940 850.010 352.200 ;
        RECT 849.780 351.460 849.920 351.940 ;
        RECT 850.150 351.460 850.470 351.520 ;
        RECT 849.780 351.320 850.470 351.460 ;
        RECT 850.150 351.260 850.470 351.320 ;
        RECT 849.230 337.860 849.550 337.920 ;
        RECT 850.150 337.860 850.470 337.920 ;
        RECT 849.230 337.720 850.470 337.860 ;
        RECT 849.230 337.660 849.550 337.720 ;
        RECT 850.150 337.660 850.470 337.720 ;
        RECT 627.510 279.380 627.830 279.440 ;
        RECT 849.230 279.380 849.550 279.440 ;
        RECT 627.510 279.240 849.550 279.380 ;
        RECT 627.510 279.180 627.830 279.240 ;
        RECT 849.230 279.180 849.550 279.240 ;
        RECT 621.070 16.900 621.390 16.960 ;
        RECT 627.510 16.900 627.830 16.960 ;
        RECT 621.070 16.760 627.830 16.900 ;
        RECT 621.070 16.700 621.390 16.760 ;
        RECT 627.510 16.700 627.830 16.760 ;
      LAYER via ;
        RECT 849.720 448.500 849.980 448.760 ;
        RECT 852.020 448.500 852.280 448.760 ;
        RECT 849.720 427.420 849.980 427.680 ;
        RECT 849.720 379.480 849.980 379.740 ;
        RECT 849.720 351.940 849.980 352.200 ;
        RECT 850.180 351.260 850.440 351.520 ;
        RECT 849.260 337.660 849.520 337.920 ;
        RECT 850.180 337.660 850.440 337.920 ;
        RECT 627.540 279.180 627.800 279.440 ;
        RECT 849.260 279.180 849.520 279.440 ;
        RECT 621.100 16.700 621.360 16.960 ;
        RECT 627.540 16.700 627.800 16.960 ;
      LAYER met2 ;
        RECT 855.370 510.410 855.650 514.000 ;
        RECT 852.540 510.270 855.650 510.410 ;
        RECT 852.540 449.210 852.680 510.270 ;
        RECT 855.370 510.000 855.650 510.270 ;
        RECT 852.080 449.070 852.680 449.210 ;
        RECT 852.080 448.790 852.220 449.070 ;
        RECT 849.720 448.470 849.980 448.790 ;
        RECT 852.020 448.470 852.280 448.790 ;
        RECT 849.780 427.710 849.920 448.470 ;
        RECT 849.720 427.390 849.980 427.710 ;
        RECT 849.720 379.450 849.980 379.770 ;
        RECT 849.780 352.230 849.920 379.450 ;
        RECT 849.720 351.910 849.980 352.230 ;
        RECT 850.180 351.230 850.440 351.550 ;
        RECT 850.240 337.950 850.380 351.230 ;
        RECT 849.260 337.630 849.520 337.950 ;
        RECT 850.180 337.630 850.440 337.950 ;
        RECT 849.320 279.470 849.460 337.630 ;
        RECT 627.540 279.150 627.800 279.470 ;
        RECT 849.260 279.150 849.520 279.470 ;
        RECT 627.600 16.990 627.740 279.150 ;
        RECT 621.100 16.670 621.360 16.990 ;
        RECT 627.540 16.670 627.800 16.990 ;
        RECT 621.160 2.400 621.300 16.670 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 120.600 117.230 120.660 ;
        RECT 489.970 120.600 490.290 120.660 ;
        RECT 116.910 120.460 490.290 120.600 ;
        RECT 116.910 120.400 117.230 120.460 ;
        RECT 489.970 120.400 490.290 120.460 ;
        RECT 115.530 14.180 115.850 14.240 ;
        RECT 116.910 14.180 117.230 14.240 ;
        RECT 115.530 14.040 117.230 14.180 ;
        RECT 115.530 13.980 115.850 14.040 ;
        RECT 116.910 13.980 117.230 14.040 ;
      LAYER via ;
        RECT 116.940 120.400 117.200 120.660 ;
        RECT 490.000 120.400 490.260 120.660 ;
        RECT 115.560 13.980 115.820 14.240 ;
        RECT 116.940 13.980 117.200 14.240 ;
      LAYER met2 ;
        RECT 492.890 510.410 493.170 514.000 ;
        RECT 490.060 510.270 493.170 510.410 ;
        RECT 490.060 120.690 490.200 510.270 ;
        RECT 492.890 510.000 493.170 510.270 ;
        RECT 116.940 120.370 117.200 120.690 ;
        RECT 490.000 120.370 490.260 120.690 ;
        RECT 117.000 14.270 117.140 120.370 ;
        RECT 115.560 13.950 115.820 14.270 ;
        RECT 116.940 13.950 117.200 14.270 ;
        RECT 115.620 2.400 115.760 13.950 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.770 400.420 504.090 400.480 ;
        RECT 507.450 400.420 507.770 400.480 ;
        RECT 503.770 400.280 507.770 400.420 ;
        RECT 503.770 400.220 504.090 400.280 ;
        RECT 507.450 400.220 507.770 400.280 ;
        RECT 144.510 382.740 144.830 382.800 ;
        RECT 503.770 382.740 504.090 382.800 ;
        RECT 144.510 382.600 504.090 382.740 ;
        RECT 144.510 382.540 144.830 382.600 ;
        RECT 503.770 382.540 504.090 382.600 ;
        RECT 139.450 20.640 139.770 20.700 ;
        RECT 144.510 20.640 144.830 20.700 ;
        RECT 139.450 20.500 144.830 20.640 ;
        RECT 139.450 20.440 139.770 20.500 ;
        RECT 144.510 20.440 144.830 20.500 ;
      LAYER via ;
        RECT 503.800 400.220 504.060 400.480 ;
        RECT 507.480 400.220 507.740 400.480 ;
        RECT 144.540 382.540 144.800 382.800 ;
        RECT 503.800 382.540 504.060 382.800 ;
        RECT 139.480 20.440 139.740 20.700 ;
        RECT 144.540 20.440 144.800 20.700 ;
      LAYER met2 ;
        RECT 509.910 510.340 510.190 514.000 ;
        RECT 509.840 510.000 510.190 510.340 ;
        RECT 509.840 483.325 509.980 510.000 ;
        RECT 507.930 482.955 508.210 483.325 ;
        RECT 509.770 482.955 510.050 483.325 ;
        RECT 508.000 400.930 508.140 482.955 ;
        RECT 507.540 400.790 508.140 400.930 ;
        RECT 507.540 400.510 507.680 400.790 ;
        RECT 503.800 400.190 504.060 400.510 ;
        RECT 507.480 400.190 507.740 400.510 ;
        RECT 503.860 382.830 504.000 400.190 ;
        RECT 144.540 382.510 144.800 382.830 ;
        RECT 503.800 382.510 504.060 382.830 ;
        RECT 144.600 20.730 144.740 382.510 ;
        RECT 139.480 20.410 139.740 20.730 ;
        RECT 144.540 20.410 144.800 20.730 ;
        RECT 139.540 2.400 139.680 20.410 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 507.930 483.000 508.210 483.280 ;
        RECT 509.770 483.000 510.050 483.280 ;
      LAYER met3 ;
        RECT 507.905 483.290 508.235 483.305 ;
        RECT 509.745 483.290 510.075 483.305 ;
        RECT 507.905 482.990 510.075 483.290 ;
        RECT 507.905 482.975 508.235 482.990 ;
        RECT 509.745 482.975 510.075 482.990 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 158.385 338.045 158.555 375.955 ;
        RECT 158.385 241.485 158.555 289.595 ;
        RECT 158.385 144.925 158.555 193.035 ;
        RECT 157.465 2.805 157.635 48.195 ;
      LAYER mcon ;
        RECT 158.385 375.785 158.555 375.955 ;
        RECT 158.385 289.425 158.555 289.595 ;
        RECT 158.385 192.865 158.555 193.035 ;
        RECT 157.465 48.025 157.635 48.195 ;
      LAYER met1 ;
        RECT 518.030 386.480 518.350 386.540 ;
        RECT 520.330 386.480 520.650 386.540 ;
        RECT 518.030 386.340 520.650 386.480 ;
        RECT 518.030 386.280 518.350 386.340 ;
        RECT 520.330 386.280 520.650 386.340 ;
        RECT 158.325 375.940 158.615 375.985 ;
        RECT 518.030 375.940 518.350 376.000 ;
        RECT 158.325 375.800 518.350 375.940 ;
        RECT 158.325 375.755 158.615 375.800 ;
        RECT 518.030 375.740 518.350 375.800 ;
        RECT 158.310 338.200 158.630 338.260 ;
        RECT 158.115 338.060 158.630 338.200 ;
        RECT 158.310 338.000 158.630 338.060 ;
        RECT 158.310 289.580 158.630 289.640 ;
        RECT 158.115 289.440 158.630 289.580 ;
        RECT 158.310 289.380 158.630 289.440 ;
        RECT 158.310 241.640 158.630 241.700 ;
        RECT 158.115 241.500 158.630 241.640 ;
        RECT 158.310 241.440 158.630 241.500 ;
        RECT 158.310 193.020 158.630 193.080 ;
        RECT 158.115 192.880 158.630 193.020 ;
        RECT 158.310 192.820 158.630 192.880 ;
        RECT 158.310 145.080 158.630 145.140 ;
        RECT 158.115 144.940 158.630 145.080 ;
        RECT 158.310 144.880 158.630 144.940 ;
        RECT 157.390 96.460 157.710 96.520 ;
        RECT 158.310 96.460 158.630 96.520 ;
        RECT 157.390 96.320 158.630 96.460 ;
        RECT 157.390 96.260 157.710 96.320 ;
        RECT 158.310 96.260 158.630 96.320 ;
        RECT 157.405 48.180 157.695 48.225 ;
        RECT 158.310 48.180 158.630 48.240 ;
        RECT 157.405 48.040 158.630 48.180 ;
        RECT 157.405 47.995 157.695 48.040 ;
        RECT 158.310 47.980 158.630 48.040 ;
        RECT 157.390 2.960 157.710 3.020 ;
        RECT 157.195 2.820 157.710 2.960 ;
        RECT 157.390 2.760 157.710 2.820 ;
      LAYER via ;
        RECT 518.060 386.280 518.320 386.540 ;
        RECT 520.360 386.280 520.620 386.540 ;
        RECT 518.060 375.740 518.320 376.000 ;
        RECT 158.340 338.000 158.600 338.260 ;
        RECT 158.340 289.380 158.600 289.640 ;
        RECT 158.340 241.440 158.600 241.700 ;
        RECT 158.340 192.820 158.600 193.080 ;
        RECT 158.340 144.880 158.600 145.140 ;
        RECT 157.420 96.260 157.680 96.520 ;
        RECT 158.340 96.260 158.600 96.520 ;
        RECT 158.340 47.980 158.600 48.240 ;
        RECT 157.420 2.760 157.680 3.020 ;
      LAYER met2 ;
        RECT 522.790 510.340 523.070 514.000 ;
        RECT 522.720 510.000 523.070 510.340 ;
        RECT 522.720 483.325 522.860 510.000 ;
        RECT 520.350 482.955 520.630 483.325 ;
        RECT 522.650 482.955 522.930 483.325 ;
        RECT 520.420 386.570 520.560 482.955 ;
        RECT 518.060 386.250 518.320 386.570 ;
        RECT 520.360 386.250 520.620 386.570 ;
        RECT 518.120 376.030 518.260 386.250 ;
        RECT 518.060 375.710 518.320 376.030 ;
        RECT 158.340 337.970 158.600 338.290 ;
        RECT 158.400 289.670 158.540 337.970 ;
        RECT 158.340 289.350 158.600 289.670 ;
        RECT 158.340 241.410 158.600 241.730 ;
        RECT 158.400 193.110 158.540 241.410 ;
        RECT 158.340 192.790 158.600 193.110 ;
        RECT 158.340 144.850 158.600 145.170 ;
        RECT 158.400 96.550 158.540 144.850 ;
        RECT 157.420 96.230 157.680 96.550 ;
        RECT 158.340 96.230 158.600 96.550 ;
        RECT 157.480 48.805 157.620 96.230 ;
        RECT 157.410 48.435 157.690 48.805 ;
        RECT 158.330 48.435 158.610 48.805 ;
        RECT 158.400 48.270 158.540 48.435 ;
        RECT 158.340 47.950 158.600 48.270 ;
        RECT 157.420 2.730 157.680 3.050 ;
        RECT 157.480 2.400 157.620 2.730 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 520.350 483.000 520.630 483.280 ;
        RECT 522.650 483.000 522.930 483.280 ;
        RECT 157.410 48.480 157.690 48.760 ;
        RECT 158.330 48.480 158.610 48.760 ;
      LAYER met3 ;
        RECT 520.325 483.290 520.655 483.305 ;
        RECT 522.625 483.290 522.955 483.305 ;
        RECT 520.325 482.990 522.955 483.290 ;
        RECT 520.325 482.975 520.655 482.990 ;
        RECT 522.625 482.975 522.955 482.990 ;
        RECT 157.385 48.770 157.715 48.785 ;
        RECT 158.305 48.770 158.635 48.785 ;
        RECT 157.385 48.470 158.635 48.770 ;
        RECT 157.385 48.455 157.715 48.470 ;
        RECT 158.305 48.455 158.635 48.470 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.370 386.480 531.690 386.540 ;
        RECT 533.210 386.480 533.530 386.540 ;
        RECT 531.370 386.340 533.530 386.480 ;
        RECT 531.370 386.280 531.690 386.340 ;
        RECT 533.210 386.280 533.530 386.340 ;
        RECT 179.010 258.640 179.330 258.700 ;
        RECT 532.290 258.640 532.610 258.700 ;
        RECT 179.010 258.500 532.610 258.640 ;
        RECT 179.010 258.440 179.330 258.500 ;
        RECT 532.290 258.440 532.610 258.500 ;
        RECT 174.870 15.200 175.190 15.260 ;
        RECT 179.010 15.200 179.330 15.260 ;
        RECT 174.870 15.060 179.330 15.200 ;
        RECT 174.870 15.000 175.190 15.060 ;
        RECT 179.010 15.000 179.330 15.060 ;
      LAYER via ;
        RECT 531.400 386.280 531.660 386.540 ;
        RECT 533.240 386.280 533.500 386.540 ;
        RECT 179.040 258.440 179.300 258.700 ;
        RECT 532.320 258.440 532.580 258.700 ;
        RECT 174.900 15.000 175.160 15.260 ;
        RECT 179.040 15.000 179.300 15.260 ;
      LAYER met2 ;
        RECT 535.670 510.340 535.950 514.000 ;
        RECT 535.600 510.000 535.950 510.340 ;
        RECT 535.600 483.325 535.740 510.000 ;
        RECT 533.230 482.955 533.510 483.325 ;
        RECT 535.530 482.955 535.810 483.325 ;
        RECT 533.300 386.570 533.440 482.955 ;
        RECT 531.400 386.250 531.660 386.570 ;
        RECT 533.240 386.250 533.500 386.570 ;
        RECT 531.460 351.970 531.600 386.250 ;
        RECT 531.460 351.830 532.520 351.970 ;
        RECT 532.380 258.730 532.520 351.830 ;
        RECT 179.040 258.410 179.300 258.730 ;
        RECT 532.320 258.410 532.580 258.730 ;
        RECT 179.100 15.290 179.240 258.410 ;
        RECT 174.900 14.970 175.160 15.290 ;
        RECT 179.040 14.970 179.300 15.290 ;
        RECT 174.960 2.400 175.100 14.970 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 533.230 483.000 533.510 483.280 ;
        RECT 535.530 483.000 535.810 483.280 ;
      LAYER met3 ;
        RECT 533.205 483.290 533.535 483.305 ;
        RECT 535.505 483.290 535.835 483.305 ;
        RECT 533.205 482.990 535.835 483.290 ;
        RECT 533.205 482.975 533.535 482.990 ;
        RECT 535.505 482.975 535.835 482.990 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 265.440 192.670 265.500 ;
        RECT 545.170 265.440 545.490 265.500 ;
        RECT 192.350 265.300 545.490 265.440 ;
        RECT 192.350 265.240 192.670 265.300 ;
        RECT 545.170 265.240 545.490 265.300 ;
      LAYER via ;
        RECT 192.380 265.240 192.640 265.500 ;
        RECT 545.200 265.240 545.460 265.500 ;
      LAYER met2 ;
        RECT 548.090 510.410 548.370 514.000 ;
        RECT 545.260 510.270 548.370 510.410 ;
        RECT 545.260 265.530 545.400 510.270 ;
        RECT 548.090 510.000 548.370 510.270 ;
        RECT 192.380 265.210 192.640 265.530 ;
        RECT 545.200 265.210 545.460 265.530 ;
        RECT 192.440 20.130 192.580 265.210 ;
        RECT 192.440 19.990 193.040 20.130 ;
        RECT 192.900 2.400 193.040 19.990 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 534.590 496.980 534.910 497.040 ;
        RECT 560.810 496.980 561.130 497.040 ;
        RECT 534.590 496.840 561.130 496.980 ;
        RECT 534.590 496.780 534.910 496.840 ;
        RECT 560.810 496.780 561.130 496.840 ;
        RECT 213.510 369.140 213.830 369.200 ;
        RECT 534.590 369.140 534.910 369.200 ;
        RECT 213.510 369.000 534.910 369.140 ;
        RECT 213.510 368.940 213.830 369.000 ;
        RECT 534.590 368.940 534.910 369.000 ;
        RECT 210.750 20.640 211.070 20.700 ;
        RECT 213.510 20.640 213.830 20.700 ;
        RECT 210.750 20.500 213.830 20.640 ;
        RECT 210.750 20.440 211.070 20.500 ;
        RECT 213.510 20.440 213.830 20.500 ;
      LAYER via ;
        RECT 534.620 496.780 534.880 497.040 ;
        RECT 560.840 496.780 561.100 497.040 ;
        RECT 213.540 368.940 213.800 369.200 ;
        RECT 534.620 368.940 534.880 369.200 ;
        RECT 210.780 20.440 211.040 20.700 ;
        RECT 213.540 20.440 213.800 20.700 ;
      LAYER met2 ;
        RECT 560.970 510.340 561.250 514.000 ;
        RECT 560.900 510.000 561.250 510.340 ;
        RECT 560.900 497.070 561.040 510.000 ;
        RECT 534.620 496.750 534.880 497.070 ;
        RECT 560.840 496.750 561.100 497.070 ;
        RECT 534.680 369.230 534.820 496.750 ;
        RECT 213.540 368.910 213.800 369.230 ;
        RECT 534.620 368.910 534.880 369.230 ;
        RECT 213.600 20.730 213.740 368.910 ;
        RECT 210.780 20.410 211.040 20.730 ;
        RECT 213.540 20.410 213.800 20.730 ;
        RECT 210.840 2.400 210.980 20.410 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 362.340 234.530 362.400 ;
        RECT 573.230 362.340 573.550 362.400 ;
        RECT 234.210 362.200 573.550 362.340 ;
        RECT 234.210 362.140 234.530 362.200 ;
        RECT 573.230 362.140 573.550 362.200 ;
        RECT 228.690 17.240 229.010 17.300 ;
        RECT 234.210 17.240 234.530 17.300 ;
        RECT 228.690 17.100 234.530 17.240 ;
        RECT 228.690 17.040 229.010 17.100 ;
        RECT 234.210 17.040 234.530 17.100 ;
      LAYER via ;
        RECT 234.240 362.140 234.500 362.400 ;
        RECT 573.260 362.140 573.520 362.400 ;
        RECT 228.720 17.040 228.980 17.300 ;
        RECT 234.240 17.040 234.500 17.300 ;
      LAYER met2 ;
        RECT 573.850 510.410 574.130 514.000 ;
        RECT 573.320 510.270 574.130 510.410 ;
        RECT 573.320 362.430 573.460 510.270 ;
        RECT 573.850 510.000 574.130 510.270 ;
        RECT 234.240 362.110 234.500 362.430 ;
        RECT 573.260 362.110 573.520 362.430 ;
        RECT 234.300 17.330 234.440 362.110 ;
        RECT 228.720 17.010 228.980 17.330 ;
        RECT 234.240 17.010 234.500 17.330 ;
        RECT 228.780 2.400 228.920 17.010 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 442.665 386.325 442.835 434.775 ;
        RECT 441.745 282.965 441.915 331.075 ;
      LAYER mcon ;
        RECT 442.665 434.605 442.835 434.775 ;
        RECT 441.745 330.905 441.915 331.075 ;
      LAYER met1 ;
        RECT 442.590 434.760 442.910 434.820 ;
        RECT 442.395 434.620 442.910 434.760 ;
        RECT 442.590 434.560 442.910 434.620 ;
        RECT 442.590 386.480 442.910 386.540 ;
        RECT 442.395 386.340 442.910 386.480 ;
        RECT 442.590 386.280 442.910 386.340 ;
        RECT 441.685 331.060 441.975 331.105 ;
        RECT 442.130 331.060 442.450 331.120 ;
        RECT 441.685 330.920 442.450 331.060 ;
        RECT 441.685 330.875 441.975 330.920 ;
        RECT 442.130 330.860 442.450 330.920 ;
        RECT 441.670 283.120 441.990 283.180 ;
        RECT 441.475 282.980 441.990 283.120 ;
        RECT 441.670 282.920 441.990 282.980 ;
        RECT 441.670 241.640 441.990 241.700 ;
        RECT 442.130 241.640 442.450 241.700 ;
        RECT 441.670 241.500 442.450 241.640 ;
        RECT 441.670 241.440 441.990 241.500 ;
        RECT 442.130 241.440 442.450 241.500 ;
        RECT 442.130 207.300 442.450 207.360 ;
        RECT 441.760 207.160 442.450 207.300 ;
        RECT 441.760 207.020 441.900 207.160 ;
        RECT 442.130 207.100 442.450 207.160 ;
        RECT 441.670 206.760 441.990 207.020 ;
        RECT 54.810 182.820 55.130 182.880 ;
        RECT 441.670 182.820 441.990 182.880 ;
        RECT 54.810 182.680 441.990 182.820 ;
        RECT 54.810 182.620 55.130 182.680 ;
        RECT 441.670 182.620 441.990 182.680 ;
        RECT 50.210 17.920 50.530 17.980 ;
        RECT 54.810 17.920 55.130 17.980 ;
        RECT 50.210 17.780 55.130 17.920 ;
        RECT 50.210 17.720 50.530 17.780 ;
        RECT 54.810 17.720 55.130 17.780 ;
      LAYER via ;
        RECT 442.620 434.560 442.880 434.820 ;
        RECT 442.620 386.280 442.880 386.540 ;
        RECT 442.160 330.860 442.420 331.120 ;
        RECT 441.700 282.920 441.960 283.180 ;
        RECT 441.700 241.440 441.960 241.700 ;
        RECT 442.160 241.440 442.420 241.700 ;
        RECT 442.160 207.100 442.420 207.360 ;
        RECT 441.700 206.760 441.960 207.020 ;
        RECT 54.840 182.620 55.100 182.880 ;
        RECT 441.700 182.620 441.960 182.880 ;
        RECT 50.240 17.720 50.500 17.980 ;
        RECT 54.840 17.720 55.100 17.980 ;
      LAYER met2 ;
        RECT 445.970 510.340 446.250 514.000 ;
        RECT 445.900 510.000 446.250 510.340 ;
        RECT 445.900 483.325 446.040 510.000 ;
        RECT 442.610 482.955 442.890 483.325 ;
        RECT 445.830 482.955 446.110 483.325 ;
        RECT 442.680 434.850 442.820 482.955 ;
        RECT 442.620 434.530 442.880 434.850 ;
        RECT 442.620 386.250 442.880 386.570 ;
        RECT 442.680 331.570 442.820 386.250 ;
        RECT 442.220 331.430 442.820 331.570 ;
        RECT 442.220 331.150 442.360 331.430 ;
        RECT 442.160 330.830 442.420 331.150 ;
        RECT 441.700 282.890 441.960 283.210 ;
        RECT 441.760 241.730 441.900 282.890 ;
        RECT 441.700 241.410 441.960 241.730 ;
        RECT 442.160 241.410 442.420 241.730 ;
        RECT 442.220 207.390 442.360 241.410 ;
        RECT 442.160 207.070 442.420 207.390 ;
        RECT 441.700 206.730 441.960 207.050 ;
        RECT 441.760 182.910 441.900 206.730 ;
        RECT 54.840 182.590 55.100 182.910 ;
        RECT 441.700 182.590 441.960 182.910 ;
        RECT 54.900 18.010 55.040 182.590 ;
        RECT 50.240 17.690 50.500 18.010 ;
        RECT 54.840 17.690 55.100 18.010 ;
        RECT 50.300 2.400 50.440 17.690 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 442.610 483.000 442.890 483.280 ;
        RECT 445.830 483.000 446.110 483.280 ;
      LAYER met3 ;
        RECT 442.585 483.290 442.915 483.305 ;
        RECT 445.805 483.290 446.135 483.305 ;
        RECT 442.585 482.990 446.135 483.290 ;
        RECT 442.585 482.975 442.915 482.990 ;
        RECT 445.805 482.975 446.135 482.990 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 586.570 472.840 586.890 472.900 ;
        RECT 588.870 472.840 589.190 472.900 ;
        RECT 586.570 472.700 589.190 472.840 ;
        RECT 586.570 472.640 586.890 472.700 ;
        RECT 588.870 472.640 589.190 472.700 ;
        RECT 254.910 189.620 255.230 189.680 ;
        RECT 586.570 189.620 586.890 189.680 ;
        RECT 254.910 189.480 586.890 189.620 ;
        RECT 254.910 189.420 255.230 189.480 ;
        RECT 586.570 189.420 586.890 189.480 ;
        RECT 252.610 17.240 252.930 17.300 ;
        RECT 254.910 17.240 255.230 17.300 ;
        RECT 252.610 17.100 255.230 17.240 ;
        RECT 252.610 17.040 252.930 17.100 ;
        RECT 254.910 17.040 255.230 17.100 ;
      LAYER via ;
        RECT 586.600 472.640 586.860 472.900 ;
        RECT 588.900 472.640 589.160 472.900 ;
        RECT 254.940 189.420 255.200 189.680 ;
        RECT 586.600 189.420 586.860 189.680 ;
        RECT 252.640 17.040 252.900 17.300 ;
        RECT 254.940 17.040 255.200 17.300 ;
      LAYER met2 ;
        RECT 590.870 510.410 591.150 514.000 ;
        RECT 588.960 510.270 591.150 510.410 ;
        RECT 588.960 472.930 589.100 510.270 ;
        RECT 590.870 510.000 591.150 510.270 ;
        RECT 586.600 472.610 586.860 472.930 ;
        RECT 588.900 472.610 589.160 472.930 ;
        RECT 586.660 189.710 586.800 472.610 ;
        RECT 254.940 189.390 255.200 189.710 ;
        RECT 586.600 189.390 586.860 189.710 ;
        RECT 255.000 17.330 255.140 189.390 ;
        RECT 252.640 17.010 252.900 17.330 ;
        RECT 254.940 17.010 255.200 17.330 ;
        RECT 252.700 2.400 252.840 17.010 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 272.580 275.930 272.640 ;
        RECT 600.370 272.580 600.690 272.640 ;
        RECT 275.610 272.440 600.690 272.580 ;
        RECT 275.610 272.380 275.930 272.440 ;
        RECT 600.370 272.380 600.690 272.440 ;
        RECT 270.090 17.240 270.410 17.300 ;
        RECT 275.610 17.240 275.930 17.300 ;
        RECT 270.090 17.100 275.930 17.240 ;
        RECT 270.090 17.040 270.410 17.100 ;
        RECT 275.610 17.040 275.930 17.100 ;
      LAYER via ;
        RECT 275.640 272.380 275.900 272.640 ;
        RECT 600.400 272.380 600.660 272.640 ;
        RECT 270.120 17.040 270.380 17.300 ;
        RECT 275.640 17.040 275.900 17.300 ;
      LAYER met2 ;
        RECT 603.750 510.410 604.030 514.000 ;
        RECT 600.460 510.270 604.030 510.410 ;
        RECT 600.460 272.670 600.600 510.270 ;
        RECT 603.750 510.000 604.030 510.270 ;
        RECT 275.640 272.350 275.900 272.670 ;
        RECT 600.400 272.350 600.660 272.670 ;
        RECT 275.700 17.330 275.840 272.350 ;
        RECT 270.120 17.010 270.380 17.330 ;
        RECT 275.640 17.010 275.900 17.330 ;
        RECT 270.180 2.400 270.320 17.010 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 355.200 289.730 355.260 ;
        RECT 614.630 355.200 614.950 355.260 ;
        RECT 289.410 355.060 614.950 355.200 ;
        RECT 289.410 355.000 289.730 355.060 ;
        RECT 614.630 355.000 614.950 355.060 ;
      LAYER via ;
        RECT 289.440 355.000 289.700 355.260 ;
        RECT 614.660 355.000 614.920 355.260 ;
      LAYER met2 ;
        RECT 616.630 510.410 616.910 514.000 ;
        RECT 614.720 510.270 616.910 510.410 ;
        RECT 614.720 355.290 614.860 510.270 ;
        RECT 616.630 510.000 616.910 510.270 ;
        RECT 289.440 354.970 289.700 355.290 ;
        RECT 614.660 354.970 614.920 355.290 ;
        RECT 289.500 17.410 289.640 354.970 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 348.400 310.430 348.460 ;
        RECT 628.430 348.400 628.750 348.460 ;
        RECT 310.110 348.260 628.750 348.400 ;
        RECT 310.110 348.200 310.430 348.260 ;
        RECT 628.430 348.200 628.750 348.260 ;
        RECT 305.970 16.900 306.290 16.960 ;
        RECT 310.110 16.900 310.430 16.960 ;
        RECT 305.970 16.760 310.430 16.900 ;
        RECT 305.970 16.700 306.290 16.760 ;
        RECT 310.110 16.700 310.430 16.760 ;
      LAYER via ;
        RECT 310.140 348.200 310.400 348.460 ;
        RECT 628.460 348.200 628.720 348.460 ;
        RECT 306.000 16.700 306.260 16.960 ;
        RECT 310.140 16.700 310.400 16.960 ;
      LAYER met2 ;
        RECT 629.510 510.410 629.790 514.000 ;
        RECT 628.520 510.270 629.790 510.410 ;
        RECT 628.520 348.490 628.660 510.270 ;
        RECT 629.510 510.000 629.790 510.270 ;
        RECT 310.140 348.170 310.400 348.490 ;
        RECT 628.460 348.170 628.720 348.490 ;
        RECT 310.200 16.990 310.340 348.170 ;
        RECT 306.000 16.670 306.260 16.990 ;
        RECT 310.140 16.670 310.400 16.990 ;
        RECT 306.060 2.400 306.200 16.670 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.450 196.760 323.770 196.820 ;
        RECT 642.230 196.760 642.550 196.820 ;
        RECT 323.450 196.620 642.550 196.760 ;
        RECT 323.450 196.560 323.770 196.620 ;
        RECT 642.230 196.560 642.550 196.620 ;
      LAYER via ;
        RECT 323.480 196.560 323.740 196.820 ;
        RECT 642.260 196.560 642.520 196.820 ;
      LAYER met2 ;
        RECT 642.390 510.340 642.670 514.000 ;
        RECT 642.320 510.000 642.670 510.340 ;
        RECT 642.320 196.850 642.460 510.000 ;
        RECT 323.480 196.530 323.740 196.850 ;
        RECT 642.260 196.530 642.520 196.850 ;
        RECT 323.540 7.890 323.680 196.530 ;
        RECT 323.540 7.750 324.140 7.890 ;
        RECT 324.000 2.400 324.140 7.750 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 649.205 386.325 649.375 434.775 ;
      LAYER mcon ;
        RECT 649.205 434.605 649.375 434.775 ;
      LAYER met1 ;
        RECT 648.670 448.700 648.990 448.760 ;
        RECT 651.890 448.700 652.210 448.760 ;
        RECT 648.670 448.560 652.210 448.700 ;
        RECT 648.670 448.500 648.990 448.560 ;
        RECT 651.890 448.500 652.210 448.560 ;
        RECT 649.145 434.760 649.435 434.805 ;
        RECT 649.590 434.760 649.910 434.820 ;
        RECT 649.145 434.620 649.910 434.760 ;
        RECT 649.145 434.575 649.435 434.620 ;
        RECT 649.590 434.560 649.910 434.620 ;
        RECT 649.130 386.480 649.450 386.540 ;
        RECT 648.935 386.340 649.450 386.480 ;
        RECT 649.130 386.280 649.450 386.340 ;
        RECT 344.610 341.600 344.930 341.660 ;
        RECT 650.050 341.600 650.370 341.660 ;
        RECT 344.610 341.460 650.370 341.600 ;
        RECT 344.610 341.400 344.930 341.460 ;
        RECT 650.050 341.400 650.370 341.460 ;
        RECT 341.390 17.240 341.710 17.300 ;
        RECT 344.610 17.240 344.930 17.300 ;
        RECT 341.390 17.100 344.930 17.240 ;
        RECT 341.390 17.040 341.710 17.100 ;
        RECT 344.610 17.040 344.930 17.100 ;
      LAYER via ;
        RECT 648.700 448.500 648.960 448.760 ;
        RECT 651.920 448.500 652.180 448.760 ;
        RECT 649.620 434.560 649.880 434.820 ;
        RECT 649.160 386.280 649.420 386.540 ;
        RECT 344.640 341.400 344.900 341.660 ;
        RECT 650.080 341.400 650.340 341.660 ;
        RECT 341.420 17.040 341.680 17.300 ;
        RECT 344.640 17.040 344.900 17.300 ;
      LAYER met2 ;
        RECT 654.810 510.410 655.090 514.000 ;
        RECT 652.440 510.270 655.090 510.410 ;
        RECT 652.440 449.210 652.580 510.270 ;
        RECT 654.810 510.000 655.090 510.270 ;
        RECT 651.980 449.070 652.580 449.210 ;
        RECT 651.980 448.790 652.120 449.070 ;
        RECT 648.700 448.530 648.960 448.790 ;
        RECT 648.700 448.470 649.820 448.530 ;
        RECT 651.920 448.470 652.180 448.790 ;
        RECT 648.760 448.390 649.820 448.470 ;
        RECT 649.680 434.850 649.820 448.390 ;
        RECT 649.620 434.530 649.880 434.850 ;
        RECT 649.160 386.250 649.420 386.570 ;
        RECT 649.220 351.970 649.360 386.250 ;
        RECT 649.220 351.830 650.280 351.970 ;
        RECT 650.140 341.690 650.280 351.830 ;
        RECT 344.640 341.370 344.900 341.690 ;
        RECT 650.080 341.370 650.340 341.690 ;
        RECT 344.700 17.330 344.840 341.370 ;
        RECT 341.420 17.010 341.680 17.330 ;
        RECT 344.640 17.010 344.900 17.330 ;
        RECT 341.480 2.400 341.620 17.010 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.470 472.840 662.790 472.900 ;
        RECT 666.150 472.840 666.470 472.900 ;
        RECT 662.470 472.700 666.470 472.840 ;
        RECT 662.470 472.640 662.790 472.700 ;
        RECT 666.150 472.640 666.470 472.700 ;
        RECT 359.330 37.980 359.650 38.040 ;
        RECT 662.470 37.980 662.790 38.040 ;
        RECT 359.330 37.840 662.790 37.980 ;
        RECT 359.330 37.780 359.650 37.840 ;
        RECT 662.470 37.780 662.790 37.840 ;
      LAYER via ;
        RECT 662.500 472.640 662.760 472.900 ;
        RECT 666.180 472.640 666.440 472.900 ;
        RECT 359.360 37.780 359.620 38.040 ;
        RECT 662.500 37.780 662.760 38.040 ;
      LAYER met2 ;
        RECT 667.690 510.410 667.970 514.000 ;
        RECT 666.240 510.270 667.970 510.410 ;
        RECT 666.240 472.930 666.380 510.270 ;
        RECT 667.690 510.000 667.970 510.270 ;
        RECT 662.500 472.610 662.760 472.930 ;
        RECT 666.180 472.610 666.440 472.930 ;
        RECT 662.560 38.070 662.700 472.610 ;
        RECT 359.360 37.750 359.620 38.070 ;
        RECT 662.500 37.750 662.760 38.070 ;
        RECT 359.420 2.400 359.560 37.750 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 676.270 472.840 676.590 472.900 ;
        RECT 679.030 472.840 679.350 472.900 ;
        RECT 676.270 472.700 679.350 472.840 ;
        RECT 676.270 472.640 676.590 472.700 ;
        RECT 679.030 472.640 679.350 472.700 ;
        RECT 379.110 286.180 379.430 286.240 ;
        RECT 676.270 286.180 676.590 286.240 ;
        RECT 379.110 286.040 676.590 286.180 ;
        RECT 379.110 285.980 379.430 286.040 ;
        RECT 676.270 285.980 676.590 286.040 ;
      LAYER via ;
        RECT 676.300 472.640 676.560 472.900 ;
        RECT 679.060 472.640 679.320 472.900 ;
        RECT 379.140 285.980 379.400 286.240 ;
        RECT 676.300 285.980 676.560 286.240 ;
      LAYER met2 ;
        RECT 680.570 510.410 680.850 514.000 ;
        RECT 679.120 510.270 680.850 510.410 ;
        RECT 679.120 472.930 679.260 510.270 ;
        RECT 680.570 510.000 680.850 510.270 ;
        RECT 676.300 472.610 676.560 472.930 ;
        RECT 679.060 472.610 679.320 472.930 ;
        RECT 676.360 286.270 676.500 472.610 ;
        RECT 379.140 285.950 379.400 286.270 ;
        RECT 676.300 285.950 676.560 286.270 ;
        RECT 379.200 16.730 379.340 285.950 ;
        RECT 377.360 16.590 379.340 16.730 ;
        RECT 377.360 2.400 377.500 16.590 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 44.780 395.530 44.840 ;
        RECT 690.070 44.780 690.390 44.840 ;
        RECT 395.210 44.640 690.390 44.780 ;
        RECT 395.210 44.580 395.530 44.640 ;
        RECT 690.070 44.580 690.390 44.640 ;
      LAYER via ;
        RECT 395.240 44.580 395.500 44.840 ;
        RECT 690.100 44.580 690.360 44.840 ;
      LAYER met2 ;
        RECT 693.450 510.410 693.730 514.000 ;
        RECT 690.160 510.270 693.730 510.410 ;
        RECT 690.160 44.870 690.300 510.270 ;
        RECT 693.450 510.000 693.730 510.270 ;
        RECT 395.240 44.550 395.500 44.870 ;
        RECT 690.100 44.550 690.360 44.870 ;
        RECT 395.300 2.400 395.440 44.550 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.610 293.320 413.930 293.380 ;
        RECT 704.330 293.320 704.650 293.380 ;
        RECT 413.610 293.180 704.650 293.320 ;
        RECT 413.610 293.120 413.930 293.180 ;
        RECT 704.330 293.120 704.650 293.180 ;
      LAYER via ;
        RECT 413.640 293.120 413.900 293.380 ;
        RECT 704.360 293.120 704.620 293.380 ;
      LAYER met2 ;
        RECT 706.330 510.410 706.610 514.000 ;
        RECT 704.420 510.270 706.610 510.410 ;
        RECT 704.420 293.410 704.560 510.270 ;
        RECT 706.330 510.000 706.610 510.270 ;
        RECT 413.640 293.090 413.900 293.410 ;
        RECT 704.360 293.090 704.620 293.410 ;
        RECT 413.700 16.050 413.840 293.090 ;
        RECT 413.240 15.910 413.840 16.050 ;
        RECT 413.240 2.400 413.380 15.910 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 334.460 75.830 334.520 ;
        RECT 462.830 334.460 463.150 334.520 ;
        RECT 75.510 334.320 463.150 334.460 ;
        RECT 75.510 334.260 75.830 334.320 ;
        RECT 462.830 334.260 463.150 334.320 ;
        RECT 74.130 14.180 74.450 14.240 ;
        RECT 75.510 14.180 75.830 14.240 ;
        RECT 74.130 14.040 75.830 14.180 ;
        RECT 74.130 13.980 74.450 14.040 ;
        RECT 75.510 13.980 75.830 14.040 ;
      LAYER via ;
        RECT 75.540 334.260 75.800 334.520 ;
        RECT 462.860 334.260 463.120 334.520 ;
        RECT 74.160 13.980 74.420 14.240 ;
        RECT 75.540 13.980 75.800 14.240 ;
      LAYER met2 ;
        RECT 462.990 510.340 463.270 514.000 ;
        RECT 462.920 510.000 463.270 510.340 ;
        RECT 462.920 334.550 463.060 510.000 ;
        RECT 75.540 334.230 75.800 334.550 ;
        RECT 462.860 334.230 463.120 334.550 ;
        RECT 75.600 14.270 75.740 334.230 ;
        RECT 74.160 13.950 74.420 14.270 ;
        RECT 75.540 13.950 75.800 14.270 ;
        RECT 74.220 2.400 74.360 13.950 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 107.000 434.630 107.060 ;
        RECT 717.670 107.000 717.990 107.060 ;
        RECT 434.310 106.860 717.990 107.000 ;
        RECT 434.310 106.800 434.630 106.860 ;
        RECT 717.670 106.800 717.990 106.860 ;
        RECT 430.630 17.580 430.950 17.640 ;
        RECT 434.310 17.580 434.630 17.640 ;
        RECT 430.630 17.440 434.630 17.580 ;
        RECT 430.630 17.380 430.950 17.440 ;
        RECT 434.310 17.380 434.630 17.440 ;
      LAYER via ;
        RECT 434.340 106.800 434.600 107.060 ;
        RECT 717.700 106.800 717.960 107.060 ;
        RECT 430.660 17.380 430.920 17.640 ;
        RECT 434.340 17.380 434.600 17.640 ;
      LAYER met2 ;
        RECT 719.210 510.410 719.490 514.000 ;
        RECT 717.760 510.270 719.490 510.410 ;
        RECT 717.760 107.090 717.900 510.270 ;
        RECT 719.210 510.000 719.490 510.270 ;
        RECT 434.340 106.770 434.600 107.090 ;
        RECT 717.700 106.770 717.960 107.090 ;
        RECT 434.400 17.670 434.540 106.770 ;
        RECT 430.660 17.350 430.920 17.670 ;
        RECT 434.340 17.350 434.600 17.670 ;
        RECT 430.720 2.400 430.860 17.350 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.010 300.120 455.330 300.180 ;
        RECT 731.930 300.120 732.250 300.180 ;
        RECT 455.010 299.980 732.250 300.120 ;
        RECT 455.010 299.920 455.330 299.980 ;
        RECT 731.930 299.920 732.250 299.980 ;
        RECT 448.570 15.200 448.890 15.260 ;
        RECT 455.010 15.200 455.330 15.260 ;
        RECT 448.570 15.060 455.330 15.200 ;
        RECT 448.570 15.000 448.890 15.060 ;
        RECT 455.010 15.000 455.330 15.060 ;
      LAYER via ;
        RECT 455.040 299.920 455.300 300.180 ;
        RECT 731.960 299.920 732.220 300.180 ;
        RECT 448.600 15.000 448.860 15.260 ;
        RECT 455.040 15.000 455.300 15.260 ;
      LAYER met2 ;
        RECT 731.630 510.340 731.910 514.000 ;
        RECT 731.560 510.000 731.910 510.340 ;
        RECT 731.560 473.690 731.700 510.000 ;
        RECT 731.560 473.550 732.160 473.690 ;
        RECT 732.020 300.210 732.160 473.550 ;
        RECT 455.040 299.890 455.300 300.210 ;
        RECT 731.960 299.890 732.220 300.210 ;
        RECT 455.100 15.290 455.240 299.890 ;
        RECT 448.600 14.970 448.860 15.290 ;
        RECT 455.040 14.970 455.300 15.290 ;
        RECT 448.660 2.400 448.800 14.970 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 739.825 193.205 739.995 207.315 ;
      LAYER mcon ;
        RECT 739.825 207.145 739.995 207.315 ;
      LAYER met1 ;
        RECT 738.370 400.420 738.690 400.480 ;
        RECT 739.290 400.420 739.610 400.480 ;
        RECT 738.370 400.280 739.610 400.420 ;
        RECT 738.370 400.220 738.690 400.280 ;
        RECT 739.290 400.220 739.610 400.280 ;
        RECT 739.290 303.320 739.610 303.580 ;
        RECT 739.380 303.180 739.520 303.320 ;
        RECT 739.750 303.180 740.070 303.240 ;
        RECT 739.380 303.040 740.070 303.180 ;
        RECT 739.750 302.980 740.070 303.040 ;
        RECT 739.750 207.300 740.070 207.360 ;
        RECT 739.555 207.160 740.070 207.300 ;
        RECT 739.750 207.100 740.070 207.160 ;
        RECT 739.750 193.360 740.070 193.420 ;
        RECT 739.555 193.220 740.070 193.360 ;
        RECT 739.750 193.160 740.070 193.220 ;
        RECT 466.510 17.240 466.830 17.300 ;
        RECT 466.510 17.100 725.260 17.240 ;
        RECT 466.510 17.040 466.830 17.100 ;
        RECT 725.120 16.900 725.260 17.100 ;
        RECT 740.210 16.900 740.530 16.960 ;
        RECT 725.120 16.760 740.530 16.900 ;
        RECT 740.210 16.700 740.530 16.760 ;
      LAYER via ;
        RECT 738.400 400.220 738.660 400.480 ;
        RECT 739.320 400.220 739.580 400.480 ;
        RECT 739.320 303.320 739.580 303.580 ;
        RECT 739.780 302.980 740.040 303.240 ;
        RECT 739.780 207.100 740.040 207.360 ;
        RECT 739.780 193.160 740.040 193.420 ;
        RECT 466.540 17.040 466.800 17.300 ;
        RECT 740.240 16.700 740.500 16.960 ;
      LAYER met2 ;
        RECT 744.510 510.410 744.790 514.000 ;
        RECT 741.680 510.270 744.790 510.410 ;
        RECT 741.680 449.210 741.820 510.270 ;
        RECT 744.510 510.000 744.790 510.270 ;
        RECT 739.840 449.070 741.820 449.210 ;
        RECT 739.840 400.930 739.980 449.070 ;
        RECT 739.380 400.790 739.980 400.930 ;
        RECT 739.380 400.510 739.520 400.790 ;
        RECT 738.400 400.190 738.660 400.510 ;
        RECT 739.320 400.190 739.580 400.510 ;
        RECT 738.460 376.450 738.600 400.190 ;
        RECT 738.460 376.310 739.060 376.450 ;
        RECT 738.920 351.290 739.060 376.310 ;
        RECT 738.920 351.150 739.520 351.290 ;
        RECT 739.380 303.610 739.520 351.150 ;
        RECT 739.320 303.290 739.580 303.610 ;
        RECT 739.780 302.950 740.040 303.270 ;
        RECT 739.840 207.390 739.980 302.950 ;
        RECT 739.780 207.070 740.040 207.390 ;
        RECT 739.780 193.130 740.040 193.450 ;
        RECT 739.840 109.890 739.980 193.130 ;
        RECT 739.840 109.750 740.440 109.890 ;
        RECT 466.540 17.010 466.800 17.330 ;
        RECT 466.600 2.400 466.740 17.010 ;
        RECT 740.300 16.990 740.440 109.750 ;
        RECT 740.240 16.670 740.500 16.990 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 511.205 16.745 511.375 17.935 ;
      LAYER mcon ;
        RECT 511.205 17.765 511.375 17.935 ;
      LAYER met1 ;
        RECT 752.170 472.840 752.490 472.900 ;
        RECT 755.390 472.840 755.710 472.900 ;
        RECT 752.170 472.700 755.710 472.840 ;
        RECT 752.170 472.640 752.490 472.700 ;
        RECT 755.390 472.640 755.710 472.700 ;
        RECT 511.145 17.920 511.435 17.965 ;
        RECT 751.710 17.920 752.030 17.980 ;
        RECT 511.145 17.780 752.030 17.920 ;
        RECT 511.145 17.735 511.435 17.780 ;
        RECT 751.710 17.720 752.030 17.780 ;
        RECT 484.450 16.900 484.770 16.960 ;
        RECT 511.145 16.900 511.435 16.945 ;
        RECT 484.450 16.760 511.435 16.900 ;
        RECT 484.450 16.700 484.770 16.760 ;
        RECT 511.145 16.715 511.435 16.760 ;
      LAYER via ;
        RECT 752.200 472.640 752.460 472.900 ;
        RECT 755.420 472.640 755.680 472.900 ;
        RECT 751.740 17.720 752.000 17.980 ;
        RECT 484.480 16.700 484.740 16.960 ;
      LAYER met2 ;
        RECT 757.390 510.410 757.670 514.000 ;
        RECT 755.480 510.270 757.670 510.410 ;
        RECT 755.480 472.930 755.620 510.270 ;
        RECT 757.390 510.000 757.670 510.270 ;
        RECT 752.200 472.610 752.460 472.930 ;
        RECT 755.420 472.610 755.680 472.930 ;
        RECT 752.260 18.090 752.400 472.610 ;
        RECT 751.800 18.010 752.400 18.090 ;
        RECT 751.740 17.950 752.400 18.010 ;
        RECT 751.740 17.690 752.000 17.950 ;
        RECT 484.480 16.670 484.740 16.990 ;
        RECT 484.540 2.400 484.680 16.670 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 767.425 145.265 767.595 159.035 ;
        RECT 766.505 89.845 766.675 137.955 ;
      LAYER mcon ;
        RECT 767.425 158.865 767.595 159.035 ;
        RECT 766.505 137.785 766.675 137.955 ;
      LAYER met1 ;
        RECT 766.890 193.700 767.210 193.760 ;
        RECT 767.350 193.700 767.670 193.760 ;
        RECT 766.890 193.560 767.670 193.700 ;
        RECT 766.890 193.500 767.210 193.560 ;
        RECT 767.350 193.500 767.670 193.560 ;
        RECT 767.350 159.020 767.670 159.080 ;
        RECT 767.155 158.880 767.670 159.020 ;
        RECT 767.350 158.820 767.670 158.880 ;
        RECT 766.890 145.420 767.210 145.480 ;
        RECT 767.365 145.420 767.655 145.465 ;
        RECT 766.890 145.280 767.655 145.420 ;
        RECT 766.890 145.220 767.210 145.280 ;
        RECT 767.365 145.235 767.655 145.280 ;
        RECT 766.430 137.940 766.750 138.000 ;
        RECT 766.235 137.800 766.750 137.940 ;
        RECT 766.430 137.740 766.750 137.800 ;
        RECT 766.445 90.000 766.735 90.045 ;
        RECT 766.890 90.000 767.210 90.060 ;
        RECT 766.445 89.860 767.210 90.000 ;
        RECT 766.445 89.815 766.735 89.860 ;
        RECT 766.890 89.800 767.210 89.860 ;
        RECT 502.390 17.920 502.710 17.980 ;
        RECT 502.390 17.780 510.900 17.920 ;
        RECT 502.390 17.720 502.710 17.780 ;
        RECT 510.760 17.580 510.900 17.780 ;
        RECT 510.760 17.440 728.020 17.580 ;
        RECT 727.880 17.240 728.020 17.440 ;
        RECT 767.350 17.240 767.670 17.300 ;
        RECT 727.880 17.100 767.670 17.240 ;
        RECT 767.350 17.040 767.670 17.100 ;
      LAYER via ;
        RECT 766.920 193.500 767.180 193.760 ;
        RECT 767.380 193.500 767.640 193.760 ;
        RECT 767.380 158.820 767.640 159.080 ;
        RECT 766.920 145.220 767.180 145.480 ;
        RECT 766.460 137.740 766.720 138.000 ;
        RECT 766.920 89.800 767.180 90.060 ;
        RECT 502.420 17.720 502.680 17.980 ;
        RECT 767.380 17.040 767.640 17.300 ;
      LAYER met2 ;
        RECT 770.270 510.340 770.550 514.000 ;
        RECT 770.200 510.000 770.550 510.340 ;
        RECT 770.200 483.325 770.340 510.000 ;
        RECT 766.910 482.955 767.190 483.325 ;
        RECT 770.130 482.955 770.410 483.325 ;
        RECT 766.980 193.790 767.120 482.955 ;
        RECT 766.920 193.470 767.180 193.790 ;
        RECT 767.380 193.470 767.640 193.790 ;
        RECT 767.440 159.110 767.580 193.470 ;
        RECT 767.380 158.790 767.640 159.110 ;
        RECT 766.920 145.250 767.180 145.510 ;
        RECT 766.520 145.190 767.180 145.250 ;
        RECT 766.520 145.110 767.120 145.190 ;
        RECT 766.520 138.030 766.660 145.110 ;
        RECT 766.460 137.710 766.720 138.030 ;
        RECT 766.920 89.770 767.180 90.090 ;
        RECT 766.980 48.010 767.120 89.770 ;
        RECT 766.980 47.870 767.580 48.010 ;
        RECT 502.420 17.690 502.680 18.010 ;
        RECT 502.480 2.400 502.620 17.690 ;
        RECT 767.440 17.330 767.580 47.870 ;
        RECT 767.380 17.010 767.640 17.330 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 766.910 483.000 767.190 483.280 ;
        RECT 770.130 483.000 770.410 483.280 ;
      LAYER met3 ;
        RECT 766.885 483.290 767.215 483.305 ;
        RECT 770.105 483.290 770.435 483.305 ;
        RECT 766.885 482.990 770.435 483.290 ;
        RECT 766.885 482.975 767.215 482.990 ;
        RECT 770.105 482.975 770.435 482.990 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 18.260 520.190 18.320 ;
        RECT 779.770 18.260 780.090 18.320 ;
        RECT 519.870 18.120 780.090 18.260 ;
        RECT 519.870 18.060 520.190 18.120 ;
        RECT 779.770 18.060 780.090 18.120 ;
      LAYER via ;
        RECT 519.900 18.060 520.160 18.320 ;
        RECT 779.800 18.060 780.060 18.320 ;
      LAYER met2 ;
        RECT 783.150 510.410 783.430 514.000 ;
        RECT 779.860 510.270 783.430 510.410 ;
        RECT 779.860 18.350 780.000 510.270 ;
        RECT 783.150 510.000 783.430 510.270 ;
        RECT 519.900 18.030 520.160 18.350 ;
        RECT 779.800 18.030 780.060 18.350 ;
        RECT 519.960 2.400 520.100 18.030 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.350 18.600 537.670 18.660 ;
        RECT 794.030 18.600 794.350 18.660 ;
        RECT 537.350 18.460 794.350 18.600 ;
        RECT 537.350 18.400 537.670 18.460 ;
        RECT 794.030 18.400 794.350 18.460 ;
      LAYER via ;
        RECT 537.380 18.400 537.640 18.660 ;
        RECT 794.060 18.400 794.320 18.660 ;
      LAYER met2 ;
        RECT 796.030 510.410 796.310 514.000 ;
        RECT 793.660 510.270 796.310 510.410 ;
        RECT 793.660 21.490 793.800 510.270 ;
        RECT 796.030 510.000 796.310 510.270 ;
        RECT 793.660 21.350 794.260 21.490 ;
        RECT 794.120 18.690 794.260 21.350 ;
        RECT 537.380 18.370 537.640 18.690 ;
        RECT 794.060 18.370 794.320 18.690 ;
        RECT 537.440 9.250 537.580 18.370 ;
        RECT 537.440 9.110 538.040 9.250 ;
        RECT 537.900 2.400 538.040 9.110 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 18.940 556.070 19.000 ;
        RECT 807.370 18.940 807.690 19.000 ;
        RECT 555.750 18.800 807.690 18.940 ;
        RECT 555.750 18.740 556.070 18.800 ;
        RECT 807.370 18.740 807.690 18.800 ;
      LAYER via ;
        RECT 555.780 18.740 556.040 19.000 ;
        RECT 807.400 18.740 807.660 19.000 ;
      LAYER met2 ;
        RECT 808.450 510.410 808.730 514.000 ;
        RECT 807.460 510.270 808.730 510.410 ;
        RECT 807.460 19.030 807.600 510.270 ;
        RECT 808.450 510.000 808.730 510.270 ;
        RECT 555.780 18.710 556.040 19.030 ;
        RECT 807.400 18.710 807.660 19.030 ;
        RECT 555.840 2.400 555.980 18.710 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 821.170 19.620 821.490 19.680 ;
        RECT 787.220 19.480 821.490 19.620 ;
        RECT 573.690 19.280 574.010 19.340 ;
        RECT 787.220 19.280 787.360 19.480 ;
        RECT 821.170 19.420 821.490 19.480 ;
        RECT 573.690 19.140 787.360 19.280 ;
        RECT 573.690 19.080 574.010 19.140 ;
      LAYER via ;
        RECT 573.720 19.080 573.980 19.340 ;
        RECT 821.200 19.420 821.460 19.680 ;
      LAYER met2 ;
        RECT 821.330 510.340 821.610 514.000 ;
        RECT 821.260 510.000 821.610 510.340 ;
        RECT 821.260 19.710 821.400 510.000 ;
        RECT 821.200 19.390 821.460 19.710 ;
        RECT 573.720 19.050 573.980 19.370 ;
        RECT 573.780 2.400 573.920 19.050 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 786.745 18.105 786.915 19.635 ;
      LAYER mcon ;
        RECT 786.745 19.465 786.915 19.635 ;
      LAYER met1 ;
        RECT 828.530 448.700 828.850 448.760 ;
        RECT 831.750 448.700 832.070 448.760 ;
        RECT 828.530 448.560 832.070 448.700 ;
        RECT 828.530 448.500 828.850 448.560 ;
        RECT 831.750 448.500 832.070 448.560 ;
        RECT 828.990 110.740 829.310 110.800 ;
        RECT 828.620 110.600 829.310 110.740 ;
        RECT 828.620 110.460 828.760 110.600 ;
        RECT 828.990 110.540 829.310 110.600 ;
        RECT 828.530 110.200 828.850 110.460 ;
        RECT 591.170 19.620 591.490 19.680 ;
        RECT 786.685 19.620 786.975 19.665 ;
        RECT 591.170 19.480 786.975 19.620 ;
        RECT 591.170 19.420 591.490 19.480 ;
        RECT 786.685 19.435 786.975 19.480 ;
        RECT 786.685 18.260 786.975 18.305 ;
        RECT 828.990 18.260 829.310 18.320 ;
        RECT 786.685 18.120 829.310 18.260 ;
        RECT 786.685 18.075 786.975 18.120 ;
        RECT 828.990 18.060 829.310 18.120 ;
      LAYER via ;
        RECT 828.560 448.500 828.820 448.760 ;
        RECT 831.780 448.500 832.040 448.760 ;
        RECT 829.020 110.540 829.280 110.800 ;
        RECT 828.560 110.200 828.820 110.460 ;
        RECT 591.200 19.420 591.460 19.680 ;
        RECT 829.020 18.060 829.280 18.320 ;
      LAYER met2 ;
        RECT 834.210 510.410 834.490 514.000 ;
        RECT 831.840 510.270 834.490 510.410 ;
        RECT 831.840 448.790 831.980 510.270 ;
        RECT 834.210 510.000 834.490 510.270 ;
        RECT 828.560 448.470 828.820 448.790 ;
        RECT 831.780 448.470 832.040 448.790 ;
        RECT 828.620 206.450 828.760 448.470 ;
        RECT 828.620 206.310 829.220 206.450 ;
        RECT 829.080 110.830 829.220 206.310 ;
        RECT 829.020 110.510 829.280 110.830 ;
        RECT 828.560 110.170 828.820 110.490 ;
        RECT 828.620 62.290 828.760 110.170 ;
        RECT 828.620 62.150 829.220 62.290 ;
        RECT 591.200 19.390 591.460 19.710 ;
        RECT 591.260 2.400 591.400 19.390 ;
        RECT 829.080 18.350 829.220 62.150 ;
        RECT 829.020 18.030 829.280 18.350 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 477.625 324.445 477.795 372.555 ;
      LAYER mcon ;
        RECT 477.625 372.385 477.795 372.555 ;
      LAYER met1 ;
        RECT 478.010 434.900 478.330 435.160 ;
        RECT 478.100 434.420 478.240 434.900 ;
        RECT 478.470 434.420 478.790 434.480 ;
        RECT 478.100 434.280 478.790 434.420 ;
        RECT 478.470 434.220 478.790 434.280 ;
        RECT 477.565 372.540 477.855 372.585 ;
        RECT 478.930 372.540 479.250 372.600 ;
        RECT 477.565 372.400 479.250 372.540 ;
        RECT 477.565 372.355 477.855 372.400 ;
        RECT 478.930 372.340 479.250 372.400 ;
        RECT 477.550 324.600 477.870 324.660 ;
        RECT 477.355 324.460 477.870 324.600 ;
        RECT 477.550 324.400 477.870 324.460 ;
        RECT 476.630 276.320 476.950 276.380 ;
        RECT 477.090 276.320 477.410 276.380 ;
        RECT 476.630 276.180 477.410 276.320 ;
        RECT 476.630 276.120 476.950 276.180 ;
        RECT 477.090 276.120 477.410 276.180 ;
        RECT 103.110 231.100 103.430 231.160 ;
        RECT 477.090 231.100 477.410 231.160 ;
        RECT 103.110 230.960 477.410 231.100 ;
        RECT 103.110 230.900 103.430 230.960 ;
        RECT 477.090 230.900 477.410 230.960 ;
        RECT 97.590 20.640 97.910 20.700 ;
        RECT 103.110 20.640 103.430 20.700 ;
        RECT 97.590 20.500 103.430 20.640 ;
        RECT 97.590 20.440 97.910 20.500 ;
        RECT 103.110 20.440 103.430 20.500 ;
      LAYER via ;
        RECT 478.040 434.900 478.300 435.160 ;
        RECT 478.500 434.220 478.760 434.480 ;
        RECT 478.960 372.340 479.220 372.600 ;
        RECT 477.580 324.400 477.840 324.660 ;
        RECT 476.660 276.120 476.920 276.380 ;
        RECT 477.120 276.120 477.380 276.380 ;
        RECT 103.140 230.900 103.400 231.160 ;
        RECT 477.120 230.900 477.380 231.160 ;
        RECT 97.620 20.440 97.880 20.700 ;
        RECT 103.140 20.440 103.400 20.700 ;
      LAYER met2 ;
        RECT 480.010 510.410 480.290 514.000 ;
        RECT 478.100 510.270 480.290 510.410 ;
        RECT 478.100 435.190 478.240 510.270 ;
        RECT 480.010 510.000 480.290 510.270 ;
        RECT 478.040 434.870 478.300 435.190 ;
        RECT 478.500 434.190 478.760 434.510 ;
        RECT 478.560 387.330 478.700 434.190 ;
        RECT 478.560 387.190 479.160 387.330 ;
        RECT 479.020 372.630 479.160 387.190 ;
        RECT 478.960 372.310 479.220 372.630 ;
        RECT 477.580 324.370 477.840 324.690 ;
        RECT 477.640 304.370 477.780 324.370 ;
        RECT 477.180 304.230 477.780 304.370 ;
        RECT 477.180 276.410 477.320 304.230 ;
        RECT 476.660 276.090 476.920 276.410 ;
        RECT 477.120 276.090 477.380 276.410 ;
        RECT 476.720 255.410 476.860 276.090 ;
        RECT 476.720 255.270 477.320 255.410 ;
        RECT 477.180 231.190 477.320 255.270 ;
        RECT 103.140 230.870 103.400 231.190 ;
        RECT 477.120 230.870 477.380 231.190 ;
        RECT 103.200 20.730 103.340 230.870 ;
        RECT 97.620 20.410 97.880 20.730 ;
        RECT 103.140 20.410 103.400 20.730 ;
        RECT 97.680 2.400 97.820 20.410 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 841.870 472.840 842.190 472.900 ;
        RECT 845.550 472.840 845.870 472.900 ;
        RECT 841.870 472.700 845.870 472.840 ;
        RECT 841.870 472.640 842.190 472.700 ;
        RECT 845.550 472.640 845.870 472.700 ;
        RECT 841.870 20.300 842.190 20.360 ;
        RECT 821.720 20.160 842.190 20.300 ;
        RECT 609.110 19.960 609.430 20.020 ;
        RECT 821.720 19.960 821.860 20.160 ;
        RECT 841.870 20.100 842.190 20.160 ;
        RECT 609.110 19.820 821.860 19.960 ;
        RECT 609.110 19.760 609.430 19.820 ;
      LAYER via ;
        RECT 841.900 472.640 842.160 472.900 ;
        RECT 845.580 472.640 845.840 472.900 ;
        RECT 609.140 19.760 609.400 20.020 ;
        RECT 841.900 20.100 842.160 20.360 ;
      LAYER met2 ;
        RECT 847.090 510.410 847.370 514.000 ;
        RECT 845.640 510.270 847.370 510.410 ;
        RECT 845.640 472.930 845.780 510.270 ;
        RECT 847.090 510.000 847.370 510.270 ;
        RECT 841.900 472.610 842.160 472.930 ;
        RECT 845.580 472.610 845.840 472.930 ;
        RECT 841.960 20.390 842.100 472.610 ;
        RECT 841.900 20.070 842.160 20.390 ;
        RECT 609.140 19.730 609.400 20.050 ;
        RECT 609.200 2.400 609.340 19.730 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 855.745 96.645 855.915 144.755 ;
        RECT 835.045 19.465 835.215 20.655 ;
      LAYER mcon ;
        RECT 855.745 144.585 855.915 144.755 ;
        RECT 835.045 20.485 835.215 20.655 ;
      LAYER met1 ;
        RECT 855.670 144.740 855.990 144.800 ;
        RECT 855.475 144.600 855.990 144.740 ;
        RECT 855.670 144.540 855.990 144.600 ;
        RECT 855.685 96.800 855.975 96.845 ;
        RECT 856.590 96.800 856.910 96.860 ;
        RECT 855.685 96.660 856.910 96.800 ;
        RECT 855.685 96.615 855.975 96.660 ;
        RECT 856.590 96.600 856.910 96.660 ;
        RECT 834.985 20.640 835.275 20.685 ;
        RECT 821.260 20.500 835.275 20.640 ;
        RECT 627.050 20.300 627.370 20.360 ;
        RECT 821.260 20.300 821.400 20.500 ;
        RECT 834.985 20.455 835.275 20.500 ;
        RECT 627.050 20.160 821.400 20.300 ;
        RECT 627.050 20.100 627.370 20.160 ;
        RECT 834.985 19.620 835.275 19.665 ;
        RECT 856.590 19.620 856.910 19.680 ;
        RECT 834.985 19.480 856.910 19.620 ;
        RECT 834.985 19.435 835.275 19.480 ;
        RECT 856.590 19.420 856.910 19.480 ;
      LAYER via ;
        RECT 855.700 144.540 855.960 144.800 ;
        RECT 856.620 96.600 856.880 96.860 ;
        RECT 627.080 20.100 627.340 20.360 ;
        RECT 856.620 19.420 856.880 19.680 ;
      LAYER met2 ;
        RECT 859.970 510.410 860.250 514.000 ;
        RECT 856.220 510.270 860.250 510.410 ;
        RECT 856.220 449.210 856.360 510.270 ;
        RECT 859.970 510.000 860.250 510.270 ;
        RECT 855.760 449.070 856.360 449.210 ;
        RECT 855.760 144.830 855.900 449.070 ;
        RECT 855.700 144.510 855.960 144.830 ;
        RECT 856.620 96.570 856.880 96.890 ;
        RECT 627.080 20.070 627.340 20.390 ;
        RECT 627.140 2.400 627.280 20.070 ;
        RECT 856.680 19.710 856.820 96.570 ;
        RECT 856.620 19.390 856.880 19.710 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 327.660 124.130 327.720 ;
        RECT 497.330 327.660 497.650 327.720 ;
        RECT 123.810 327.520 497.650 327.660 ;
        RECT 123.810 327.460 124.130 327.520 ;
        RECT 497.330 327.460 497.650 327.520 ;
        RECT 121.510 20.640 121.830 20.700 ;
        RECT 123.810 20.640 124.130 20.700 ;
        RECT 121.510 20.500 124.130 20.640 ;
        RECT 121.510 20.440 121.830 20.500 ;
        RECT 123.810 20.440 124.130 20.500 ;
      LAYER via ;
        RECT 123.840 327.460 124.100 327.720 ;
        RECT 497.360 327.460 497.620 327.720 ;
        RECT 121.540 20.440 121.800 20.700 ;
        RECT 123.840 20.440 124.100 20.700 ;
      LAYER met2 ;
        RECT 497.030 510.340 497.310 514.000 ;
        RECT 496.960 510.000 497.310 510.340 ;
        RECT 496.960 473.690 497.100 510.000 ;
        RECT 496.960 473.550 497.560 473.690 ;
        RECT 497.420 327.750 497.560 473.550 ;
        RECT 123.840 327.430 124.100 327.750 ;
        RECT 497.360 327.430 497.620 327.750 ;
        RECT 123.900 20.730 124.040 327.430 ;
        RECT 121.540 20.410 121.800 20.730 ;
        RECT 123.840 20.410 124.100 20.730 ;
        RECT 121.600 2.400 121.740 20.410 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 151.410 237.900 151.730 237.960 ;
        RECT 510.670 237.900 510.990 237.960 ;
        RECT 151.410 237.760 510.990 237.900 ;
        RECT 151.410 237.700 151.730 237.760 ;
        RECT 510.670 237.700 510.990 237.760 ;
        RECT 145.430 19.280 145.750 19.340 ;
        RECT 151.410 19.280 151.730 19.340 ;
        RECT 145.430 19.140 151.730 19.280 ;
        RECT 145.430 19.080 145.750 19.140 ;
        RECT 151.410 19.080 151.730 19.140 ;
      LAYER via ;
        RECT 151.440 237.700 151.700 237.960 ;
        RECT 510.700 237.700 510.960 237.960 ;
        RECT 145.460 19.080 145.720 19.340 ;
        RECT 151.440 19.080 151.700 19.340 ;
      LAYER met2 ;
        RECT 514.050 510.410 514.330 514.000 ;
        RECT 510.760 510.270 514.330 510.410 ;
        RECT 510.760 237.990 510.900 510.270 ;
        RECT 514.050 510.000 514.330 510.270 ;
        RECT 151.440 237.670 151.700 237.990 ;
        RECT 510.700 237.670 510.960 237.990 ;
        RECT 151.500 19.370 151.640 237.670 ;
        RECT 145.460 19.050 145.720 19.370 ;
        RECT 151.440 19.050 151.700 19.370 ;
        RECT 145.520 2.400 145.660 19.050 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 19.280 163.690 19.340 ;
        RECT 163.370 19.140 497.560 19.280 ;
        RECT 163.370 19.080 163.690 19.140 ;
        RECT 497.420 18.940 497.560 19.140 ;
        RECT 524.470 18.940 524.790 19.000 ;
        RECT 497.420 18.800 524.790 18.940 ;
        RECT 524.470 18.740 524.790 18.800 ;
      LAYER via ;
        RECT 163.400 19.080 163.660 19.340 ;
        RECT 524.500 18.740 524.760 19.000 ;
      LAYER met2 ;
        RECT 526.930 510.410 527.210 514.000 ;
        RECT 524.560 510.270 527.210 510.410 ;
        RECT 163.400 19.050 163.660 19.370 ;
        RECT 163.460 2.400 163.600 19.050 ;
        RECT 524.560 19.030 524.700 510.270 ;
        RECT 526.930 510.000 527.210 510.270 ;
        RECT 524.500 18.710 524.760 19.030 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 19.960 181.170 20.020 ;
        RECT 538.270 19.960 538.590 20.020 ;
        RECT 180.850 19.820 538.590 19.960 ;
        RECT 180.850 19.760 181.170 19.820 ;
        RECT 538.270 19.760 538.590 19.820 ;
      LAYER via ;
        RECT 180.880 19.760 181.140 20.020 ;
        RECT 538.300 19.760 538.560 20.020 ;
      LAYER met2 ;
        RECT 539.810 510.410 540.090 514.000 ;
        RECT 538.360 510.270 540.090 510.410 ;
        RECT 538.360 20.050 538.500 510.270 ;
        RECT 539.810 510.000 540.090 510.270 ;
        RECT 180.880 19.730 181.140 20.050 ;
        RECT 538.300 19.730 538.560 20.050 ;
        RECT 180.940 2.400 181.080 19.730 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 19.620 199.110 19.680 ;
        RECT 552.070 19.620 552.390 19.680 ;
        RECT 198.790 19.480 552.390 19.620 ;
        RECT 198.790 19.420 199.110 19.480 ;
        RECT 552.070 19.420 552.390 19.480 ;
      LAYER via ;
        RECT 198.820 19.420 199.080 19.680 ;
        RECT 552.100 19.420 552.360 19.680 ;
      LAYER met2 ;
        RECT 552.690 510.410 552.970 514.000 ;
        RECT 552.160 510.270 552.970 510.410 ;
        RECT 552.160 19.710 552.300 510.270 ;
        RECT 552.690 510.000 552.970 510.270 ;
        RECT 198.820 19.390 199.080 19.710 ;
        RECT 552.100 19.390 552.360 19.710 ;
        RECT 198.880 2.400 199.020 19.390 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 559.505 282.965 559.675 331.075 ;
        RECT 560.425 59.245 560.595 96.475 ;
      LAYER mcon ;
        RECT 559.505 330.905 559.675 331.075 ;
        RECT 560.425 96.305 560.595 96.475 ;
      LAYER met1 ;
        RECT 558.970 386.480 559.290 386.540 ;
        RECT 560.350 386.480 560.670 386.540 ;
        RECT 558.970 386.340 560.670 386.480 ;
        RECT 558.970 386.280 559.290 386.340 ;
        RECT 560.350 386.280 560.670 386.340 ;
        RECT 558.970 331.060 559.290 331.120 ;
        RECT 559.445 331.060 559.735 331.105 ;
        RECT 558.970 330.920 559.735 331.060 ;
        RECT 558.970 330.860 559.290 330.920 ;
        RECT 559.445 330.875 559.735 330.920 ;
        RECT 559.430 283.120 559.750 283.180 ;
        RECT 559.235 282.980 559.750 283.120 ;
        RECT 559.430 282.920 559.750 282.980 ;
        RECT 558.970 145.080 559.290 145.140 ;
        RECT 560.350 145.080 560.670 145.140 ;
        RECT 558.970 144.940 560.670 145.080 ;
        RECT 558.970 144.880 559.290 144.940 ;
        RECT 560.350 144.880 560.670 144.940 ;
        RECT 559.430 110.400 559.750 110.460 ;
        RECT 560.350 110.400 560.670 110.460 ;
        RECT 559.430 110.260 560.670 110.400 ;
        RECT 559.430 110.200 559.750 110.260 ;
        RECT 560.350 110.200 560.670 110.260 ;
        RECT 560.350 96.460 560.670 96.520 ;
        RECT 560.155 96.320 560.670 96.460 ;
        RECT 560.350 96.260 560.670 96.320 ;
        RECT 560.350 59.400 560.670 59.460 ;
        RECT 560.155 59.260 560.670 59.400 ;
        RECT 560.350 59.200 560.670 59.260 ;
        RECT 216.730 20.300 217.050 20.360 ;
        RECT 560.350 20.300 560.670 20.360 ;
        RECT 216.730 20.160 560.670 20.300 ;
        RECT 216.730 20.100 217.050 20.160 ;
        RECT 560.350 20.100 560.670 20.160 ;
      LAYER via ;
        RECT 559.000 386.280 559.260 386.540 ;
        RECT 560.380 386.280 560.640 386.540 ;
        RECT 559.000 330.860 559.260 331.120 ;
        RECT 559.460 282.920 559.720 283.180 ;
        RECT 559.000 144.880 559.260 145.140 ;
        RECT 560.380 144.880 560.640 145.140 ;
        RECT 559.460 110.200 559.720 110.460 ;
        RECT 560.380 110.200 560.640 110.460 ;
        RECT 560.380 96.260 560.640 96.520 ;
        RECT 560.380 59.200 560.640 59.460 ;
        RECT 216.760 20.100 217.020 20.360 ;
        RECT 560.380 20.100 560.640 20.360 ;
      LAYER met2 ;
        RECT 565.570 510.410 565.850 514.000 ;
        RECT 563.200 510.270 565.850 510.410 ;
        RECT 563.200 449.210 563.340 510.270 ;
        RECT 565.570 510.000 565.850 510.270 ;
        RECT 561.360 449.070 563.340 449.210 ;
        RECT 561.360 448.530 561.500 449.070 ;
        RECT 559.980 448.390 561.500 448.530 ;
        RECT 559.980 400.930 560.120 448.390 ;
        RECT 559.980 400.790 560.580 400.930 ;
        RECT 560.440 386.570 560.580 400.790 ;
        RECT 559.000 386.250 559.260 386.570 ;
        RECT 560.380 386.250 560.640 386.570 ;
        RECT 559.060 331.150 559.200 386.250 ;
        RECT 559.000 330.830 559.260 331.150 ;
        RECT 559.460 282.890 559.720 283.210 ;
        RECT 559.520 255.410 559.660 282.890 ;
        RECT 559.060 255.270 559.660 255.410 ;
        RECT 559.060 241.130 559.200 255.270 ;
        RECT 559.060 240.990 559.660 241.130 ;
        RECT 559.520 216.650 559.660 240.990 ;
        RECT 559.060 216.510 559.660 216.650 ;
        RECT 559.060 193.645 559.200 216.510 ;
        RECT 558.990 193.275 559.270 193.645 ;
        RECT 558.990 192.595 559.270 192.965 ;
        RECT 559.060 145.170 559.200 192.595 ;
        RECT 559.000 144.850 559.260 145.170 ;
        RECT 560.380 144.850 560.640 145.170 ;
        RECT 560.440 110.570 560.580 144.850 ;
        RECT 559.520 110.490 560.580 110.570 ;
        RECT 559.460 110.430 560.640 110.490 ;
        RECT 559.460 110.170 559.720 110.430 ;
        RECT 560.380 110.170 560.640 110.430 ;
        RECT 560.440 96.550 560.580 110.170 ;
        RECT 560.380 96.230 560.640 96.550 ;
        RECT 560.380 59.170 560.640 59.490 ;
        RECT 560.440 20.390 560.580 59.170 ;
        RECT 216.760 20.070 217.020 20.390 ;
        RECT 560.380 20.070 560.640 20.390 ;
        RECT 216.820 2.400 216.960 20.070 ;
        RECT 216.610 -4.800 217.170 2.400 ;
      LAYER via2 ;
        RECT 558.990 193.320 559.270 193.600 ;
        RECT 558.990 192.640 559.270 192.920 ;
      LAYER met3 ;
        RECT 558.965 193.610 559.295 193.625 ;
        RECT 558.965 193.310 559.970 193.610 ;
        RECT 558.965 193.295 559.295 193.310 ;
        RECT 558.965 192.930 559.295 192.945 ;
        RECT 559.670 192.930 559.970 193.310 ;
        RECT 558.965 192.630 559.970 192.930 ;
        RECT 558.965 192.615 559.295 192.630 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 572.770 472.840 573.090 472.900 ;
        RECT 575.990 472.840 576.310 472.900 ;
        RECT 572.770 472.700 576.310 472.840 ;
        RECT 572.770 472.640 573.090 472.700 ;
        RECT 575.990 472.640 576.310 472.700 ;
        RECT 234.670 20.640 234.990 20.700 ;
        RECT 234.670 20.500 561.040 20.640 ;
        RECT 234.670 20.440 234.990 20.500 ;
        RECT 560.900 20.300 561.040 20.500 ;
        RECT 572.770 20.300 573.090 20.360 ;
        RECT 560.900 20.160 573.090 20.300 ;
        RECT 572.770 20.100 573.090 20.160 ;
      LAYER via ;
        RECT 572.800 472.640 573.060 472.900 ;
        RECT 576.020 472.640 576.280 472.900 ;
        RECT 234.700 20.440 234.960 20.700 ;
        RECT 572.800 20.100 573.060 20.360 ;
      LAYER met2 ;
        RECT 577.990 510.410 578.270 514.000 ;
        RECT 576.080 510.270 578.270 510.410 ;
        RECT 576.080 472.930 576.220 510.270 ;
        RECT 577.990 510.000 578.270 510.270 ;
        RECT 572.800 472.610 573.060 472.930 ;
        RECT 576.020 472.610 576.280 472.930 ;
        RECT 234.700 20.410 234.960 20.730 ;
        RECT 234.760 2.400 234.900 20.410 ;
        RECT 572.860 20.390 573.000 472.610 ;
        RECT 572.800 20.070 573.060 20.390 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 56.190 17.780 448.890 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 448.570 17.720 448.890 17.780 ;
      LAYER via ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 448.600 17.720 448.860 17.980 ;
      LAYER met2 ;
        RECT 450.110 510.410 450.390 514.000 ;
        RECT 448.660 510.270 450.390 510.410 ;
        RECT 448.660 18.010 448.800 510.270 ;
        RECT 450.110 510.000 450.390 510.270 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 462.370 472.840 462.690 472.900 ;
        RECT 465.590 472.840 465.910 472.900 ;
        RECT 462.370 472.700 465.910 472.840 ;
        RECT 462.370 472.640 462.690 472.700 ;
        RECT 465.590 472.640 465.910 472.700 ;
        RECT 80.110 18.260 80.430 18.320 ;
        RECT 462.370 18.260 462.690 18.320 ;
        RECT 80.110 18.120 462.690 18.260 ;
        RECT 80.110 18.060 80.430 18.120 ;
        RECT 462.370 18.060 462.690 18.120 ;
      LAYER via ;
        RECT 462.400 472.640 462.660 472.900 ;
        RECT 465.620 472.640 465.880 472.900 ;
        RECT 80.140 18.060 80.400 18.320 ;
        RECT 462.400 18.060 462.660 18.320 ;
      LAYER met2 ;
        RECT 467.130 510.410 467.410 514.000 ;
        RECT 465.680 510.270 467.410 510.410 ;
        RECT 465.680 472.930 465.820 510.270 ;
        RECT 467.130 510.000 467.410 510.270 ;
        RECT 462.400 472.610 462.660 472.930 ;
        RECT 465.620 472.610 465.880 472.930 ;
        RECT 462.460 18.350 462.600 472.610 ;
        RECT 80.140 18.030 80.400 18.350 ;
        RECT 462.400 18.030 462.660 18.350 ;
        RECT 80.200 2.400 80.340 18.030 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 103.570 18.600 103.890 18.660 ;
        RECT 483.070 18.600 483.390 18.660 ;
        RECT 103.570 18.460 483.390 18.600 ;
        RECT 103.570 18.400 103.890 18.460 ;
        RECT 483.070 18.400 483.390 18.460 ;
      LAYER via ;
        RECT 103.600 18.400 103.860 18.660 ;
        RECT 483.100 18.400 483.360 18.660 ;
      LAYER met2 ;
        RECT 484.150 510.410 484.430 514.000 ;
        RECT 483.160 510.270 484.430 510.410 ;
        RECT 483.160 18.690 483.300 510.270 ;
        RECT 484.150 510.000 484.430 510.270 ;
        RECT 103.600 18.370 103.860 18.690 ;
        RECT 483.100 18.370 483.360 18.690 ;
        RECT 103.660 2.400 103.800 18.370 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.870 472.840 497.190 472.900 ;
        RECT 499.630 472.840 499.950 472.900 ;
        RECT 496.870 472.700 499.950 472.840 ;
        RECT 496.870 472.640 497.190 472.700 ;
        RECT 499.630 472.640 499.950 472.700 ;
        RECT 127.490 18.940 127.810 19.000 ;
        RECT 496.870 18.940 497.190 19.000 ;
        RECT 127.490 18.800 497.190 18.940 ;
        RECT 127.490 18.740 127.810 18.800 ;
        RECT 496.870 18.740 497.190 18.800 ;
      LAYER via ;
        RECT 496.900 472.640 497.160 472.900 ;
        RECT 499.660 472.640 499.920 472.900 ;
        RECT 127.520 18.740 127.780 19.000 ;
        RECT 496.900 18.740 497.160 19.000 ;
      LAYER met2 ;
        RECT 501.170 510.410 501.450 514.000 ;
        RECT 499.720 510.270 501.450 510.410 ;
        RECT 499.720 472.930 499.860 510.270 ;
        RECT 501.170 510.000 501.450 510.270 ;
        RECT 496.900 472.610 497.160 472.930 ;
        RECT 499.660 472.610 499.920 472.930 ;
        RECT 496.960 19.030 497.100 472.610 ;
        RECT 127.520 18.710 127.780 19.030 ;
        RECT 496.900 18.710 497.160 19.030 ;
        RECT 127.580 2.400 127.720 18.710 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 48.445 15.725 48.615 16.915 ;
        RECT 111.005 16.575 111.175 16.915 ;
        RECT 158.385 16.745 159.475 16.915 ;
        RECT 96.285 15.725 96.455 16.575 ;
        RECT 110.085 16.405 111.175 16.575 ;
      LAYER mcon ;
        RECT 48.445 16.745 48.615 16.915 ;
        RECT 111.005 16.745 111.175 16.915 ;
        RECT 159.305 16.745 159.475 16.915 ;
        RECT 96.285 16.405 96.455 16.575 ;
      LAYER met1 ;
        RECT 192.900 17.100 228.460 17.240 ;
        RECT 26.290 16.900 26.610 16.960 ;
        RECT 48.385 16.900 48.675 16.945 ;
        RECT 26.290 16.760 48.675 16.900 ;
        RECT 26.290 16.700 26.610 16.760 ;
        RECT 48.385 16.715 48.675 16.760 ;
        RECT 110.945 16.900 111.235 16.945 ;
        RECT 158.325 16.900 158.615 16.945 ;
        RECT 110.945 16.760 158.615 16.900 ;
        RECT 110.945 16.715 111.235 16.760 ;
        RECT 158.325 16.715 158.615 16.760 ;
        RECT 159.245 16.900 159.535 16.945 ;
        RECT 192.900 16.900 193.040 17.100 ;
        RECT 159.245 16.760 193.040 16.900 ;
        RECT 159.245 16.715 159.535 16.760 ;
        RECT 96.225 16.560 96.515 16.605 ;
        RECT 110.025 16.560 110.315 16.605 ;
        RECT 96.225 16.420 110.315 16.560 ;
        RECT 228.320 16.560 228.460 17.100 ;
        RECT 358.960 17.100 372.900 17.240 ;
        RECT 358.960 16.900 359.100 17.100 ;
        RECT 372.760 16.900 372.900 17.100 ;
        RECT 317.560 16.760 359.100 16.900 ;
        RECT 372.300 16.760 372.900 16.900 ;
        RECT 317.560 16.560 317.700 16.760 ;
        RECT 228.320 16.420 317.700 16.560 ;
        RECT 96.225 16.375 96.515 16.420 ;
        RECT 110.025 16.375 110.315 16.420 ;
        RECT 372.300 16.220 372.440 16.760 ;
        RECT 428.330 16.220 428.650 16.280 ;
        RECT 372.300 16.080 428.650 16.220 ;
        RECT 428.330 16.020 428.650 16.080 ;
        RECT 48.385 15.880 48.675 15.925 ;
        RECT 96.225 15.880 96.515 15.925 ;
        RECT 48.385 15.740 96.515 15.880 ;
        RECT 48.385 15.695 48.675 15.740 ;
        RECT 96.225 15.695 96.515 15.740 ;
      LAYER via ;
        RECT 26.320 16.700 26.580 16.960 ;
        RECT 428.360 16.020 428.620 16.280 ;
      LAYER met2 ;
        RECT 428.950 510.410 429.230 514.000 ;
        RECT 428.420 510.270 429.230 510.410 ;
        RECT 26.320 16.670 26.580 16.990 ;
        RECT 26.380 2.400 26.520 16.670 ;
        RECT 428.420 16.310 428.560 510.270 ;
        RECT 428.950 510.000 429.230 510.270 ;
        RECT 428.360 15.990 428.620 16.310 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 430.705 386.325 430.875 434.775 ;
        RECT 428.865 331.245 429.035 338.895 ;
        RECT 428.865 235.025 429.035 282.795 ;
        RECT 428.865 17.085 429.035 48.195 ;
      LAYER mcon ;
        RECT 430.705 434.605 430.875 434.775 ;
        RECT 428.865 338.725 429.035 338.895 ;
        RECT 428.865 282.625 429.035 282.795 ;
        RECT 428.865 48.025 429.035 48.195 ;
      LAYER met1 ;
        RECT 430.630 434.760 430.950 434.820 ;
        RECT 430.435 434.620 430.950 434.760 ;
        RECT 430.630 434.560 430.950 434.620 ;
        RECT 429.250 386.480 429.570 386.540 ;
        RECT 430.645 386.480 430.935 386.525 ;
        RECT 429.250 386.340 430.935 386.480 ;
        RECT 429.250 386.280 429.570 386.340 ;
        RECT 430.645 386.295 430.935 386.340 ;
        RECT 428.790 338.880 429.110 338.940 ;
        RECT 428.595 338.740 429.110 338.880 ;
        RECT 428.790 338.680 429.110 338.740 ;
        RECT 428.790 331.400 429.110 331.460 ;
        RECT 428.595 331.260 429.110 331.400 ;
        RECT 428.790 331.200 429.110 331.260 ;
        RECT 428.790 282.780 429.110 282.840 ;
        RECT 428.595 282.640 429.110 282.780 ;
        RECT 428.790 282.580 429.110 282.640 ;
        RECT 428.790 235.180 429.110 235.240 ;
        RECT 428.595 235.040 429.110 235.180 ;
        RECT 428.790 234.980 429.110 235.040 ;
        RECT 428.790 234.500 429.110 234.560 ;
        RECT 430.170 234.500 430.490 234.560 ;
        RECT 428.790 234.360 430.490 234.500 ;
        RECT 428.790 234.300 429.110 234.360 ;
        RECT 430.170 234.300 430.490 234.360 ;
        RECT 429.710 110.740 430.030 110.800 ;
        RECT 428.880 110.600 430.030 110.740 ;
        RECT 428.880 110.460 429.020 110.600 ;
        RECT 429.710 110.540 430.030 110.600 ;
        RECT 428.790 110.200 429.110 110.460 ;
        RECT 428.790 48.180 429.110 48.240 ;
        RECT 428.595 48.040 429.110 48.180 ;
        RECT 428.790 47.980 429.110 48.040 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 32.270 17.440 373.360 17.580 ;
        RECT 32.270 17.380 32.590 17.440 ;
        RECT 373.220 17.240 373.360 17.440 ;
        RECT 428.805 17.240 429.095 17.285 ;
        RECT 373.220 17.100 429.095 17.240 ;
        RECT 428.805 17.055 429.095 17.100 ;
      LAYER via ;
        RECT 430.660 434.560 430.920 434.820 ;
        RECT 429.280 386.280 429.540 386.540 ;
        RECT 428.820 338.680 429.080 338.940 ;
        RECT 428.820 331.200 429.080 331.460 ;
        RECT 428.820 282.580 429.080 282.840 ;
        RECT 428.820 234.980 429.080 235.240 ;
        RECT 428.820 234.300 429.080 234.560 ;
        RECT 430.200 234.300 430.460 234.560 ;
        RECT 429.740 110.540 430.000 110.800 ;
        RECT 428.820 110.200 429.080 110.460 ;
        RECT 428.820 47.980 429.080 48.240 ;
        RECT 32.300 17.380 32.560 17.640 ;
      LAYER met2 ;
        RECT 433.090 510.410 433.370 514.000 ;
        RECT 431.640 510.270 433.370 510.410 ;
        RECT 431.640 449.210 431.780 510.270 ;
        RECT 433.090 510.000 433.370 510.270 ;
        RECT 430.720 449.070 431.780 449.210 ;
        RECT 430.720 434.850 430.860 449.070 ;
        RECT 430.660 434.530 430.920 434.850 ;
        RECT 429.280 386.250 429.540 386.570 ;
        RECT 429.340 385.970 429.480 386.250 ;
        RECT 428.880 385.830 429.480 385.970 ;
        RECT 428.880 338.970 429.020 385.830 ;
        RECT 428.820 338.650 429.080 338.970 ;
        RECT 428.820 331.170 429.080 331.490 ;
        RECT 428.880 282.870 429.020 331.170 ;
        RECT 428.820 282.550 429.080 282.870 ;
        RECT 428.820 234.950 429.080 235.270 ;
        RECT 428.880 234.590 429.020 234.950 ;
        RECT 428.820 234.270 429.080 234.590 ;
        RECT 430.200 234.270 430.460 234.590 ;
        RECT 430.260 158.170 430.400 234.270 ;
        RECT 429.800 158.030 430.400 158.170 ;
        RECT 429.800 110.830 429.940 158.030 ;
        RECT 429.740 110.510 430.000 110.830 ;
        RECT 428.820 110.170 429.080 110.490 ;
        RECT 428.880 48.270 429.020 110.170 ;
        RECT 428.820 47.950 429.080 48.270 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 32.360 2.400 32.500 17.350 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 3010.000 547.020 3528.900 ;
        RECT 724.020 3010.000 727.020 3528.900 ;
        RECT 904.020 3010.000 907.020 3528.900 ;
        RECT 1084.020 3010.000 1087.020 3528.900 ;
        RECT 1264.020 3010.000 1267.020 3528.900 ;
        RECT 1444.020 3010.000 1447.020 3528.900 ;
        RECT 1624.020 3010.000 1627.020 3528.900 ;
        RECT 1804.020 3010.000 1807.020 3528.900 ;
        RECT 1984.020 3010.000 1987.020 3528.900 ;
        RECT 2164.020 3010.000 2167.020 3528.900 ;
        RECT 2344.020 3010.000 2347.020 3528.900 ;
        RECT 544.020 -9.220 547.020 510.000 ;
        RECT 724.020 -9.220 727.020 510.000 ;
        RECT 904.020 -9.220 907.020 510.000 ;
        RECT 1084.020 -9.220 1087.020 510.000 ;
        RECT 1264.020 -9.220 1267.020 510.000 ;
        RECT 1444.020 -9.220 1447.020 510.000 ;
        RECT 1624.020 -9.220 1627.020 510.000 ;
        RECT 1804.020 -9.220 1807.020 510.000 ;
        RECT 1984.020 -9.220 1987.020 510.000 ;
        RECT 2164.020 -9.220 2167.020 510.000 ;
        RECT 2344.020 -9.220 2347.020 510.000 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3010.000 457.020 3528.900 ;
        RECT 634.020 3010.000 637.020 3528.900 ;
        RECT 814.020 3010.000 817.020 3528.900 ;
        RECT 994.020 3010.000 997.020 3528.900 ;
        RECT 1174.020 3010.000 1177.020 3528.900 ;
        RECT 1354.020 3010.000 1357.020 3528.900 ;
        RECT 1534.020 3010.000 1537.020 3528.900 ;
        RECT 1714.020 3010.000 1717.020 3528.900 ;
        RECT 1894.020 3010.000 1897.020 3528.900 ;
        RECT 2074.020 3010.000 2077.020 3528.900 ;
        RECT 2254.020 3010.000 2257.020 3528.900 ;
        RECT 2434.020 3010.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 510.000 ;
        RECT 634.020 -9.220 637.020 510.000 ;
        RECT 814.020 -9.220 817.020 510.000 ;
        RECT 994.020 -9.220 997.020 510.000 ;
        RECT 1174.020 -9.220 1177.020 510.000 ;
        RECT 1354.020 -9.220 1357.020 510.000 ;
        RECT 1534.020 -9.220 1537.020 510.000 ;
        RECT 1714.020 -9.220 1717.020 510.000 ;
        RECT 1894.020 -9.220 1897.020 510.000 ;
        RECT 2074.020 -9.220 2077.020 510.000 ;
        RECT 2254.020 -9.220 2257.020 510.000 ;
        RECT 2434.020 -9.220 2437.020 510.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 3010.000 565.020 3538.100 ;
        RECT 742.020 3010.000 745.020 3538.100 ;
        RECT 922.020 3010.000 925.020 3538.100 ;
        RECT 1102.020 3010.000 1105.020 3538.100 ;
        RECT 1282.020 3010.000 1285.020 3538.100 ;
        RECT 1462.020 3010.000 1465.020 3538.100 ;
        RECT 1642.020 3010.000 1645.020 3538.100 ;
        RECT 1822.020 3010.000 1825.020 3538.100 ;
        RECT 2002.020 3010.000 2005.020 3538.100 ;
        RECT 2182.020 3010.000 2185.020 3538.100 ;
        RECT 2362.020 3010.000 2365.020 3538.100 ;
        RECT 562.020 -18.420 565.020 510.000 ;
        RECT 742.020 -18.420 745.020 510.000 ;
        RECT 922.020 -18.420 925.020 510.000 ;
        RECT 1102.020 -18.420 1105.020 510.000 ;
        RECT 1282.020 -18.420 1285.020 510.000 ;
        RECT 1462.020 -18.420 1465.020 510.000 ;
        RECT 1642.020 -18.420 1645.020 510.000 ;
        RECT 1822.020 -18.420 1825.020 510.000 ;
        RECT 2002.020 -18.420 2005.020 510.000 ;
        RECT 2182.020 -18.420 2185.020 510.000 ;
        RECT 2362.020 -18.420 2365.020 510.000 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3010.000 475.020 3538.100 ;
        RECT 652.020 3010.000 655.020 3538.100 ;
        RECT 832.020 3010.000 835.020 3538.100 ;
        RECT 1012.020 3010.000 1015.020 3538.100 ;
        RECT 1192.020 3010.000 1195.020 3538.100 ;
        RECT 1372.020 3010.000 1375.020 3538.100 ;
        RECT 1552.020 3010.000 1555.020 3538.100 ;
        RECT 1732.020 3010.000 1735.020 3538.100 ;
        RECT 1912.020 3010.000 1915.020 3538.100 ;
        RECT 2092.020 3010.000 2095.020 3538.100 ;
        RECT 2272.020 3010.000 2275.020 3538.100 ;
        RECT 2452.020 3010.000 2455.020 3538.100 ;
        RECT 472.020 -18.420 475.020 510.000 ;
        RECT 652.020 -18.420 655.020 510.000 ;
        RECT 832.020 -18.420 835.020 510.000 ;
        RECT 1012.020 -18.420 1015.020 510.000 ;
        RECT 1192.020 -18.420 1195.020 510.000 ;
        RECT 1372.020 -18.420 1375.020 510.000 ;
        RECT 1552.020 -18.420 1555.020 510.000 ;
        RECT 1732.020 -18.420 1735.020 510.000 ;
        RECT 1912.020 -18.420 1915.020 510.000 ;
        RECT 2092.020 -18.420 2095.020 510.000 ;
        RECT 2272.020 -18.420 2275.020 510.000 ;
        RECT 2452.020 -18.420 2455.020 510.000 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 3010.000 583.020 3547.300 ;
        RECT 760.020 3010.000 763.020 3547.300 ;
        RECT 940.020 3010.000 943.020 3547.300 ;
        RECT 1120.020 3010.000 1123.020 3547.300 ;
        RECT 1300.020 3010.000 1303.020 3547.300 ;
        RECT 1480.020 3010.000 1483.020 3547.300 ;
        RECT 1660.020 3010.000 1663.020 3547.300 ;
        RECT 1840.020 3010.000 1843.020 3547.300 ;
        RECT 2020.020 3010.000 2023.020 3547.300 ;
        RECT 2200.020 3010.000 2203.020 3547.300 ;
        RECT 2380.020 3010.000 2383.020 3547.300 ;
        RECT 580.020 -27.620 583.020 510.000 ;
        RECT 760.020 -27.620 763.020 510.000 ;
        RECT 940.020 -27.620 943.020 510.000 ;
        RECT 1120.020 -27.620 1123.020 510.000 ;
        RECT 1300.020 -27.620 1303.020 510.000 ;
        RECT 1480.020 -27.620 1483.020 510.000 ;
        RECT 1660.020 -27.620 1663.020 510.000 ;
        RECT 1840.020 -27.620 1843.020 510.000 ;
        RECT 2020.020 -27.620 2023.020 510.000 ;
        RECT 2200.020 -27.620 2203.020 510.000 ;
        RECT 2380.020 -27.620 2383.020 510.000 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 3010.000 493.020 3547.300 ;
        RECT 670.020 3010.000 673.020 3547.300 ;
        RECT 850.020 3010.000 853.020 3547.300 ;
        RECT 1030.020 3010.000 1033.020 3547.300 ;
        RECT 1210.020 3010.000 1213.020 3547.300 ;
        RECT 1390.020 3010.000 1393.020 3547.300 ;
        RECT 1570.020 3010.000 1573.020 3547.300 ;
        RECT 1750.020 3010.000 1753.020 3547.300 ;
        RECT 1930.020 3010.000 1933.020 3547.300 ;
        RECT 2110.020 3010.000 2113.020 3547.300 ;
        RECT 2290.020 3010.000 2293.020 3547.300 ;
        RECT 2470.020 3010.000 2473.020 3547.300 ;
        RECT 490.020 -27.620 493.020 510.000 ;
        RECT 670.020 -27.620 673.020 510.000 ;
        RECT 850.020 -27.620 853.020 510.000 ;
        RECT 1030.020 -27.620 1033.020 510.000 ;
        RECT 1210.020 -27.620 1213.020 510.000 ;
        RECT 1390.020 -27.620 1393.020 510.000 ;
        RECT 1570.020 -27.620 1573.020 510.000 ;
        RECT 1750.020 -27.620 1753.020 510.000 ;
        RECT 1930.020 -27.620 1933.020 510.000 ;
        RECT 2110.020 -27.620 2113.020 510.000 ;
        RECT 2290.020 -27.620 2293.020 510.000 ;
        RECT 2470.020 -27.620 2473.020 510.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3010.000 421.020 3556.500 ;
        RECT 598.020 3010.000 601.020 3556.500 ;
        RECT 778.020 3010.000 781.020 3556.500 ;
        RECT 958.020 3010.000 961.020 3556.500 ;
        RECT 1138.020 3010.000 1141.020 3556.500 ;
        RECT 1318.020 3010.000 1321.020 3556.500 ;
        RECT 1498.020 3010.000 1501.020 3556.500 ;
        RECT 1678.020 3010.000 1681.020 3556.500 ;
        RECT 1858.020 3010.000 1861.020 3556.500 ;
        RECT 2038.020 3010.000 2041.020 3556.500 ;
        RECT 2218.020 3010.000 2221.020 3556.500 ;
        RECT 2398.020 3010.000 2401.020 3556.500 ;
        RECT 418.020 -36.820 421.020 510.000 ;
        RECT 598.020 -36.820 601.020 510.000 ;
        RECT 778.020 -36.820 781.020 510.000 ;
        RECT 958.020 -36.820 961.020 510.000 ;
        RECT 1138.020 -36.820 1141.020 510.000 ;
        RECT 1318.020 -36.820 1321.020 510.000 ;
        RECT 1498.020 -36.820 1501.020 510.000 ;
        RECT 1678.020 -36.820 1681.020 510.000 ;
        RECT 1858.020 -36.820 1861.020 510.000 ;
        RECT 2038.020 -36.820 2041.020 510.000 ;
        RECT 2218.020 -36.820 2221.020 510.000 ;
        RECT 2398.020 -36.820 2401.020 510.000 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 3010.000 511.020 3556.500 ;
        RECT 688.020 3010.000 691.020 3556.500 ;
        RECT 868.020 3010.000 871.020 3556.500 ;
        RECT 1048.020 3010.000 1051.020 3556.500 ;
        RECT 1228.020 3010.000 1231.020 3556.500 ;
        RECT 1408.020 3010.000 1411.020 3556.500 ;
        RECT 1588.020 3010.000 1591.020 3556.500 ;
        RECT 1768.020 3010.000 1771.020 3556.500 ;
        RECT 1948.020 3010.000 1951.020 3556.500 ;
        RECT 2128.020 3010.000 2131.020 3556.500 ;
        RECT 2308.020 3010.000 2311.020 3556.500 ;
        RECT 2488.020 3010.000 2491.020 3556.500 ;
        RECT 508.020 -36.820 511.020 510.000 ;
        RECT 688.020 -36.820 691.020 510.000 ;
        RECT 868.020 -36.820 871.020 510.000 ;
        RECT 1048.020 -36.820 1051.020 510.000 ;
        RECT 1228.020 -36.820 1231.020 510.000 ;
        RECT 1408.020 -36.820 1411.020 510.000 ;
        RECT 1588.020 -36.820 1591.020 510.000 ;
        RECT 1768.020 -36.820 1771.020 510.000 ;
        RECT 1948.020 -36.820 1951.020 510.000 ;
        RECT 2128.020 -36.820 2131.020 510.000 ;
        RECT 2308.020 -36.820 2311.020 510.000 ;
        RECT 2488.020 -36.820 2491.020 510.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 415.520 520.795 2504.380 2998.885 ;
      LAYER met1 ;
        RECT 411.910 520.640 2504.380 2999.040 ;
      LAYER met2 ;
        RECT 411.940 3005.720 443.390 3006.010 ;
      LAYER met2 ;
        RECT 443.670 3006.000 443.950 3010.000 ;
      LAYER met2 ;
        RECT 444.230 3005.720 511.010 3006.010 ;
      LAYER met2 ;
        RECT 511.290 3006.000 511.570 3010.000 ;
      LAYER met2 ;
        RECT 511.850 3005.720 578.630 3006.010 ;
      LAYER met2 ;
        RECT 578.910 3006.000 579.190 3010.000 ;
      LAYER met2 ;
        RECT 579.470 3005.720 646.250 3006.010 ;
      LAYER met2 ;
        RECT 646.530 3006.000 646.810 3010.000 ;
      LAYER met2 ;
        RECT 647.090 3005.720 714.330 3006.010 ;
        RECT 715.170 3005.720 781.950 3006.010 ;
        RECT 782.790 3005.720 849.570 3006.010 ;
        RECT 850.410 3005.720 917.190 3006.010 ;
        RECT 918.030 3005.720 985.270 3006.010 ;
        RECT 986.110 3005.720 1052.890 3006.010 ;
        RECT 1053.730 3005.720 1120.510 3006.010 ;
        RECT 1121.350 3005.720 1188.130 3006.010 ;
        RECT 1188.970 3005.720 1256.210 3006.010 ;
        RECT 1257.050 3005.720 1323.830 3006.010 ;
        RECT 1324.670 3005.720 1391.450 3006.010 ;
        RECT 1392.290 3005.720 1459.070 3006.010 ;
        RECT 1459.910 3005.720 1527.150 3006.010 ;
        RECT 1527.990 3005.720 1594.770 3006.010 ;
        RECT 1595.610 3005.720 1662.390 3006.010 ;
        RECT 1663.230 3005.720 1730.010 3006.010 ;
        RECT 1730.850 3005.720 1798.090 3006.010 ;
        RECT 1798.930 3005.720 1865.710 3006.010 ;
        RECT 1866.550 3005.720 1933.330 3006.010 ;
        RECT 1934.170 3005.720 2000.950 3006.010 ;
        RECT 2001.790 3005.720 2069.030 3006.010 ;
        RECT 2069.870 3005.720 2136.650 3006.010 ;
        RECT 2137.490 3005.720 2204.270 3006.010 ;
        RECT 2205.110 3005.720 2271.890 3006.010 ;
        RECT 2272.730 3005.720 2339.970 3006.010 ;
        RECT 2340.810 3005.720 2407.590 3006.010 ;
        RECT 2408.430 3005.720 2475.210 3006.010 ;
        RECT 2476.050 3005.720 2498.770 3006.010 ;
        RECT 411.940 514.280 2498.770 3005.720 ;
        RECT 412.490 514.000 415.790 514.280 ;
        RECT 416.630 514.000 419.930 514.280 ;
        RECT 420.770 514.000 424.070 514.280 ;
        RECT 424.910 514.000 428.670 514.280 ;
        RECT 429.510 514.000 432.810 514.280 ;
        RECT 433.650 514.000 436.950 514.280 ;
        RECT 437.790 514.000 441.090 514.280 ;
        RECT 441.930 514.000 445.690 514.280 ;
        RECT 446.530 514.000 449.830 514.280 ;
        RECT 450.670 514.000 453.970 514.280 ;
        RECT 454.810 514.000 458.570 514.280 ;
        RECT 459.410 514.000 462.710 514.280 ;
        RECT 463.550 514.000 466.850 514.280 ;
        RECT 467.690 514.000 470.990 514.280 ;
        RECT 471.830 514.000 475.590 514.280 ;
        RECT 476.430 514.000 479.730 514.280 ;
        RECT 480.570 514.000 483.870 514.280 ;
        RECT 484.710 514.000 488.470 514.280 ;
        RECT 489.310 514.000 492.610 514.280 ;
        RECT 493.450 514.000 496.750 514.280 ;
        RECT 497.590 514.000 500.890 514.280 ;
        RECT 501.730 514.000 505.490 514.280 ;
        RECT 506.330 514.000 509.630 514.280 ;
        RECT 510.470 514.000 513.770 514.280 ;
        RECT 514.610 514.000 517.910 514.280 ;
        RECT 518.750 514.000 522.510 514.280 ;
        RECT 523.350 514.000 526.650 514.280 ;
        RECT 527.490 514.000 530.790 514.280 ;
        RECT 531.630 514.000 535.390 514.280 ;
        RECT 536.230 514.000 539.530 514.280 ;
        RECT 540.370 514.000 543.670 514.280 ;
        RECT 544.510 514.000 547.810 514.280 ;
        RECT 548.650 514.000 552.410 514.280 ;
        RECT 553.250 514.000 556.550 514.280 ;
        RECT 557.390 514.000 560.690 514.280 ;
        RECT 561.530 514.000 565.290 514.280 ;
        RECT 566.130 514.000 569.430 514.280 ;
        RECT 570.270 514.000 573.570 514.280 ;
        RECT 574.410 514.000 577.710 514.280 ;
        RECT 578.550 514.000 582.310 514.280 ;
        RECT 583.150 514.000 586.450 514.280 ;
        RECT 587.290 514.000 590.590 514.280 ;
        RECT 591.430 514.000 594.730 514.280 ;
        RECT 595.570 514.000 599.330 514.280 ;
        RECT 600.170 514.000 603.470 514.280 ;
        RECT 604.310 514.000 607.610 514.280 ;
        RECT 608.450 514.000 612.210 514.280 ;
        RECT 613.050 514.000 616.350 514.280 ;
        RECT 617.190 514.000 620.490 514.280 ;
        RECT 621.330 514.000 624.630 514.280 ;
        RECT 625.470 514.000 629.230 514.280 ;
        RECT 630.070 514.000 633.370 514.280 ;
        RECT 634.210 514.000 637.510 514.280 ;
        RECT 638.350 514.000 642.110 514.280 ;
        RECT 642.950 514.000 646.250 514.280 ;
        RECT 647.090 514.000 650.390 514.280 ;
        RECT 651.230 514.000 654.530 514.280 ;
        RECT 655.370 514.000 659.130 514.280 ;
        RECT 659.970 514.000 663.270 514.280 ;
        RECT 664.110 514.000 667.410 514.280 ;
        RECT 668.250 514.000 671.550 514.280 ;
        RECT 672.390 514.000 676.150 514.280 ;
        RECT 676.990 514.000 680.290 514.280 ;
        RECT 681.130 514.000 684.430 514.280 ;
        RECT 685.270 514.000 689.030 514.280 ;
        RECT 689.870 514.000 693.170 514.280 ;
        RECT 694.010 514.000 697.310 514.280 ;
        RECT 698.150 514.000 701.450 514.280 ;
        RECT 702.290 514.000 706.050 514.280 ;
        RECT 706.890 514.000 710.190 514.280 ;
        RECT 711.030 514.000 714.330 514.280 ;
        RECT 715.170 514.000 718.930 514.280 ;
        RECT 719.770 514.000 723.070 514.280 ;
        RECT 723.910 514.000 727.210 514.280 ;
        RECT 728.050 514.000 731.350 514.280 ;
        RECT 732.190 514.000 735.950 514.280 ;
        RECT 736.790 514.000 740.090 514.280 ;
        RECT 740.930 514.000 744.230 514.280 ;
        RECT 745.070 514.000 748.370 514.280 ;
        RECT 749.210 514.000 752.970 514.280 ;
        RECT 753.810 514.000 757.110 514.280 ;
        RECT 757.950 514.000 761.250 514.280 ;
        RECT 762.090 514.000 765.850 514.280 ;
        RECT 766.690 514.000 769.990 514.280 ;
        RECT 770.830 514.000 774.130 514.280 ;
        RECT 774.970 514.000 778.270 514.280 ;
        RECT 779.110 514.000 782.870 514.280 ;
        RECT 783.710 514.000 787.010 514.280 ;
        RECT 787.850 514.000 791.150 514.280 ;
        RECT 791.990 514.000 795.750 514.280 ;
        RECT 796.590 514.000 799.890 514.280 ;
        RECT 800.730 514.000 804.030 514.280 ;
        RECT 804.870 514.000 808.170 514.280 ;
        RECT 809.010 514.000 812.770 514.280 ;
        RECT 813.610 514.000 816.910 514.280 ;
        RECT 817.750 514.000 821.050 514.280 ;
        RECT 821.890 514.000 825.650 514.280 ;
        RECT 826.490 514.000 829.790 514.280 ;
        RECT 830.630 514.000 833.930 514.280 ;
        RECT 834.770 514.000 838.070 514.280 ;
        RECT 838.910 514.000 842.670 514.280 ;
        RECT 843.510 514.000 846.810 514.280 ;
        RECT 847.650 514.000 850.950 514.280 ;
        RECT 851.790 514.000 855.090 514.280 ;
        RECT 855.930 514.000 859.690 514.280 ;
        RECT 860.530 514.000 863.830 514.280 ;
        RECT 864.670 514.000 867.970 514.280 ;
        RECT 868.810 514.000 872.570 514.280 ;
        RECT 873.410 514.000 876.710 514.280 ;
        RECT 877.550 514.000 880.850 514.280 ;
        RECT 881.690 514.000 884.990 514.280 ;
        RECT 885.830 514.000 889.590 514.280 ;
        RECT 890.430 514.000 893.730 514.280 ;
        RECT 894.570 514.000 897.870 514.280 ;
        RECT 898.710 514.000 902.470 514.280 ;
        RECT 903.310 514.000 906.610 514.280 ;
        RECT 907.450 514.000 910.750 514.280 ;
        RECT 911.590 514.000 914.890 514.280 ;
        RECT 915.730 514.000 919.490 514.280 ;
        RECT 920.330 514.000 923.630 514.280 ;
        RECT 924.470 514.000 927.770 514.280 ;
        RECT 928.610 514.000 931.910 514.280 ;
        RECT 932.750 514.000 936.510 514.280 ;
        RECT 937.350 514.000 940.650 514.280 ;
        RECT 941.490 514.000 944.790 514.280 ;
        RECT 945.630 514.000 949.390 514.280 ;
        RECT 950.230 514.000 953.530 514.280 ;
        RECT 954.370 514.000 957.670 514.280 ;
        RECT 958.510 514.000 961.810 514.280 ;
        RECT 962.650 514.000 966.410 514.280 ;
        RECT 967.250 514.000 970.550 514.280 ;
        RECT 971.390 514.000 974.690 514.280 ;
        RECT 975.530 514.000 979.290 514.280 ;
        RECT 980.130 514.000 983.430 514.280 ;
        RECT 984.270 514.000 987.570 514.280 ;
        RECT 988.410 514.000 991.710 514.280 ;
        RECT 992.550 514.000 996.310 514.280 ;
        RECT 997.150 514.000 1000.450 514.280 ;
        RECT 1001.290 514.000 1004.590 514.280 ;
        RECT 1005.430 514.000 1008.730 514.280 ;
        RECT 1009.570 514.000 1013.330 514.280 ;
        RECT 1014.170 514.000 1017.470 514.280 ;
        RECT 1018.310 514.000 1021.610 514.280 ;
        RECT 1022.450 514.000 1026.210 514.280 ;
        RECT 1027.050 514.000 1030.350 514.280 ;
        RECT 1031.190 514.000 1034.490 514.280 ;
        RECT 1035.330 514.000 1038.630 514.280 ;
        RECT 1039.470 514.000 1043.230 514.280 ;
        RECT 1044.070 514.000 1047.370 514.280 ;
        RECT 1048.210 514.000 1051.510 514.280 ;
        RECT 1052.350 514.000 1056.110 514.280 ;
        RECT 1056.950 514.000 1060.250 514.280 ;
        RECT 1061.090 514.000 1064.390 514.280 ;
        RECT 1065.230 514.000 1068.530 514.280 ;
        RECT 1069.370 514.000 1073.130 514.280 ;
        RECT 1073.970 514.000 1077.270 514.280 ;
        RECT 1078.110 514.000 1081.410 514.280 ;
        RECT 1082.250 514.000 1085.550 514.280 ;
        RECT 1086.390 514.000 1090.150 514.280 ;
        RECT 1090.990 514.000 1094.290 514.280 ;
        RECT 1095.130 514.000 1098.430 514.280 ;
        RECT 1099.270 514.000 1103.030 514.280 ;
        RECT 1103.870 514.000 1107.170 514.280 ;
        RECT 1108.010 514.000 1111.310 514.280 ;
        RECT 1112.150 514.000 1115.450 514.280 ;
        RECT 1116.290 514.000 1120.050 514.280 ;
        RECT 1120.890 514.000 1124.190 514.280 ;
        RECT 1125.030 514.000 1128.330 514.280 ;
        RECT 1129.170 514.000 1132.930 514.280 ;
        RECT 1133.770 514.000 1137.070 514.280 ;
        RECT 1137.910 514.000 1141.210 514.280 ;
        RECT 1142.050 514.000 1145.350 514.280 ;
        RECT 1146.190 514.000 1149.950 514.280 ;
        RECT 1150.790 514.000 1154.090 514.280 ;
        RECT 1154.930 514.000 1158.230 514.280 ;
        RECT 1159.070 514.000 1162.830 514.280 ;
        RECT 1163.670 514.000 1166.970 514.280 ;
        RECT 1167.810 514.000 1171.110 514.280 ;
        RECT 1171.950 514.000 1175.250 514.280 ;
        RECT 1176.090 514.000 1179.850 514.280 ;
        RECT 1180.690 514.000 1183.990 514.280 ;
        RECT 1184.830 514.000 1188.130 514.280 ;
        RECT 1188.970 514.000 1192.270 514.280 ;
        RECT 1193.110 514.000 1196.870 514.280 ;
        RECT 1197.710 514.000 1201.010 514.280 ;
        RECT 1201.850 514.000 1205.150 514.280 ;
        RECT 1205.990 514.000 1209.750 514.280 ;
        RECT 1210.590 514.000 1213.890 514.280 ;
        RECT 1214.730 514.000 1218.030 514.280 ;
        RECT 1218.870 514.000 1222.170 514.280 ;
        RECT 1223.010 514.000 1226.770 514.280 ;
        RECT 1227.610 514.000 1230.910 514.280 ;
        RECT 1231.750 514.000 1235.050 514.280 ;
        RECT 1235.890 514.000 1239.650 514.280 ;
        RECT 1240.490 514.000 1243.790 514.280 ;
        RECT 1244.630 514.000 1247.930 514.280 ;
        RECT 1248.770 514.000 1252.070 514.280 ;
        RECT 1252.910 514.000 1256.670 514.280 ;
        RECT 1257.510 514.000 1260.810 514.280 ;
        RECT 1261.650 514.000 1264.950 514.280 ;
        RECT 1265.790 514.000 1269.090 514.280 ;
        RECT 1269.930 514.000 1273.690 514.280 ;
        RECT 1274.530 514.000 1277.830 514.280 ;
        RECT 1278.670 514.000 1281.970 514.280 ;
        RECT 1282.810 514.000 1286.570 514.280 ;
        RECT 1287.410 514.000 1290.710 514.280 ;
        RECT 1291.550 514.000 1294.850 514.280 ;
        RECT 1295.690 514.000 1298.990 514.280 ;
        RECT 1299.830 514.000 1303.590 514.280 ;
        RECT 1304.430 514.000 1307.730 514.280 ;
        RECT 1308.570 514.000 1311.870 514.280 ;
        RECT 1312.710 514.000 1316.470 514.280 ;
        RECT 1317.310 514.000 1320.610 514.280 ;
        RECT 1321.450 514.000 1324.750 514.280 ;
        RECT 1325.590 514.000 1328.890 514.280 ;
        RECT 1329.730 514.000 1333.490 514.280 ;
        RECT 1334.330 514.000 1337.630 514.280 ;
        RECT 1338.470 514.000 1341.770 514.280 ;
        RECT 1342.610 514.000 1345.910 514.280 ;
        RECT 1346.750 514.000 1350.510 514.280 ;
        RECT 1351.350 514.000 1354.650 514.280 ;
        RECT 1355.490 514.000 1358.790 514.280 ;
        RECT 1359.630 514.000 1363.390 514.280 ;
        RECT 1364.230 514.000 1367.530 514.280 ;
        RECT 1368.370 514.000 1371.670 514.280 ;
        RECT 1372.510 514.000 1375.810 514.280 ;
        RECT 1376.650 514.000 1380.410 514.280 ;
        RECT 1381.250 514.000 1384.550 514.280 ;
        RECT 1385.390 514.000 1388.690 514.280 ;
        RECT 1389.530 514.000 1393.290 514.280 ;
        RECT 1394.130 514.000 1397.430 514.280 ;
        RECT 1398.270 514.000 1401.570 514.280 ;
        RECT 1402.410 514.000 1405.710 514.280 ;
        RECT 1406.550 514.000 1410.310 514.280 ;
        RECT 1411.150 514.000 1414.450 514.280 ;
        RECT 1415.290 514.000 1418.590 514.280 ;
        RECT 1419.430 514.000 1422.730 514.280 ;
        RECT 1423.570 514.000 1427.330 514.280 ;
        RECT 1428.170 514.000 1431.470 514.280 ;
        RECT 1432.310 514.000 1435.610 514.280 ;
        RECT 1436.450 514.000 1440.210 514.280 ;
        RECT 1441.050 514.000 1444.350 514.280 ;
        RECT 1445.190 514.000 1448.490 514.280 ;
        RECT 1449.330 514.000 1452.630 514.280 ;
        RECT 1453.470 514.000 1457.230 514.280 ;
        RECT 1458.070 514.000 1461.370 514.280 ;
        RECT 1462.210 514.000 1465.510 514.280 ;
        RECT 1466.350 514.000 1470.110 514.280 ;
        RECT 1470.950 514.000 1474.250 514.280 ;
        RECT 1475.090 514.000 1478.390 514.280 ;
        RECT 1479.230 514.000 1482.530 514.280 ;
        RECT 1483.370 514.000 1487.130 514.280 ;
        RECT 1487.970 514.000 1491.270 514.280 ;
        RECT 1492.110 514.000 1495.410 514.280 ;
        RECT 1496.250 514.000 1500.010 514.280 ;
        RECT 1500.850 514.000 1504.150 514.280 ;
        RECT 1504.990 514.000 1508.290 514.280 ;
        RECT 1509.130 514.000 1512.430 514.280 ;
        RECT 1513.270 514.000 1517.030 514.280 ;
        RECT 1517.870 514.000 1521.170 514.280 ;
        RECT 1522.010 514.000 1525.310 514.280 ;
        RECT 1526.150 514.000 1529.450 514.280 ;
        RECT 1530.290 514.000 1534.050 514.280 ;
        RECT 1534.890 514.000 1538.190 514.280 ;
        RECT 1539.030 514.000 1542.330 514.280 ;
        RECT 1543.170 514.000 1546.930 514.280 ;
        RECT 1547.770 514.000 1551.070 514.280 ;
        RECT 1551.910 514.000 1555.210 514.280 ;
        RECT 1556.050 514.000 1559.350 514.280 ;
        RECT 1560.190 514.000 1563.950 514.280 ;
        RECT 1564.790 514.000 1568.090 514.280 ;
        RECT 1568.930 514.000 1572.230 514.280 ;
        RECT 1573.070 514.000 1576.830 514.280 ;
        RECT 1577.670 514.000 1580.970 514.280 ;
        RECT 1581.810 514.000 1585.110 514.280 ;
        RECT 1585.950 514.000 1589.250 514.280 ;
        RECT 1590.090 514.000 1593.850 514.280 ;
        RECT 1594.690 514.000 1597.990 514.280 ;
        RECT 1598.830 514.000 1602.130 514.280 ;
        RECT 1602.970 514.000 1606.270 514.280 ;
        RECT 1607.110 514.000 1610.870 514.280 ;
        RECT 1611.710 514.000 1615.010 514.280 ;
        RECT 1615.850 514.000 1619.150 514.280 ;
        RECT 1619.990 514.000 1623.750 514.280 ;
        RECT 1624.590 514.000 1627.890 514.280 ;
        RECT 1628.730 514.000 1632.030 514.280 ;
        RECT 1632.870 514.000 1636.170 514.280 ;
        RECT 1637.010 514.000 1640.770 514.280 ;
        RECT 1641.610 514.000 1644.910 514.280 ;
        RECT 1645.750 514.000 1649.050 514.280 ;
        RECT 1649.890 514.000 1653.650 514.280 ;
        RECT 1654.490 514.000 1657.790 514.280 ;
        RECT 1658.630 514.000 1661.930 514.280 ;
        RECT 1662.770 514.000 1666.070 514.280 ;
        RECT 1666.910 514.000 1670.670 514.280 ;
        RECT 1671.510 514.000 1674.810 514.280 ;
        RECT 1675.650 514.000 1678.950 514.280 ;
        RECT 1679.790 514.000 1683.090 514.280 ;
        RECT 1683.930 514.000 1687.690 514.280 ;
        RECT 1688.530 514.000 1691.830 514.280 ;
        RECT 1692.670 514.000 1695.970 514.280 ;
        RECT 1696.810 514.000 1700.570 514.280 ;
        RECT 1701.410 514.000 1704.710 514.280 ;
        RECT 1705.550 514.000 1708.850 514.280 ;
        RECT 1709.690 514.000 1712.990 514.280 ;
        RECT 1713.830 514.000 1717.590 514.280 ;
        RECT 1718.430 514.000 1721.730 514.280 ;
        RECT 1722.570 514.000 1725.870 514.280 ;
        RECT 1726.710 514.000 1730.470 514.280 ;
        RECT 1731.310 514.000 1734.610 514.280 ;
        RECT 1735.450 514.000 1738.750 514.280 ;
        RECT 1739.590 514.000 1742.890 514.280 ;
        RECT 1743.730 514.000 1747.490 514.280 ;
        RECT 1748.330 514.000 1751.630 514.280 ;
        RECT 1752.470 514.000 1755.770 514.280 ;
        RECT 1756.610 514.000 1759.910 514.280 ;
        RECT 1760.750 514.000 1764.510 514.280 ;
        RECT 1765.350 514.000 1768.650 514.280 ;
        RECT 1769.490 514.000 1772.790 514.280 ;
        RECT 1773.630 514.000 1777.390 514.280 ;
        RECT 1778.230 514.000 1781.530 514.280 ;
        RECT 1782.370 514.000 1785.670 514.280 ;
        RECT 1786.510 514.000 1789.810 514.280 ;
        RECT 1790.650 514.000 1794.410 514.280 ;
        RECT 1795.250 514.000 1798.550 514.280 ;
        RECT 1799.390 514.000 1802.690 514.280 ;
        RECT 1803.530 514.000 1807.290 514.280 ;
        RECT 1808.130 514.000 1811.430 514.280 ;
        RECT 1812.270 514.000 1815.570 514.280 ;
        RECT 1816.410 514.000 1819.710 514.280 ;
        RECT 1820.550 514.000 1824.310 514.280 ;
        RECT 1825.150 514.000 1828.450 514.280 ;
        RECT 1829.290 514.000 1832.590 514.280 ;
        RECT 1833.430 514.000 1837.190 514.280 ;
        RECT 1838.030 514.000 1841.330 514.280 ;
        RECT 1842.170 514.000 1845.470 514.280 ;
        RECT 1846.310 514.000 1849.610 514.280 ;
        RECT 1850.450 514.000 1854.210 514.280 ;
        RECT 1855.050 514.000 1858.350 514.280 ;
        RECT 1859.190 514.000 1862.490 514.280 ;
        RECT 1863.330 514.000 1866.630 514.280 ;
        RECT 1867.470 514.000 1871.230 514.280 ;
        RECT 1872.070 514.000 1875.370 514.280 ;
        RECT 1876.210 514.000 1879.510 514.280 ;
        RECT 1880.350 514.000 1884.110 514.280 ;
        RECT 1884.950 514.000 1888.250 514.280 ;
        RECT 1889.090 514.000 1892.390 514.280 ;
        RECT 1893.230 514.000 1896.530 514.280 ;
        RECT 1897.370 514.000 1901.130 514.280 ;
        RECT 1901.970 514.000 1905.270 514.280 ;
        RECT 1906.110 514.000 1909.410 514.280 ;
        RECT 1910.250 514.000 1914.010 514.280 ;
        RECT 1914.850 514.000 1918.150 514.280 ;
        RECT 1918.990 514.000 1922.290 514.280 ;
        RECT 1923.130 514.000 1926.430 514.280 ;
        RECT 1927.270 514.000 1931.030 514.280 ;
        RECT 1931.870 514.000 1935.170 514.280 ;
        RECT 1936.010 514.000 1939.310 514.280 ;
        RECT 1940.150 514.000 1943.450 514.280 ;
        RECT 1944.290 514.000 1948.050 514.280 ;
        RECT 1948.890 514.000 1952.190 514.280 ;
        RECT 1953.030 514.000 1956.330 514.280 ;
        RECT 1957.170 514.000 1960.930 514.280 ;
        RECT 1961.770 514.000 1965.070 514.280 ;
        RECT 1965.910 514.000 1969.210 514.280 ;
        RECT 1970.050 514.000 1973.350 514.280 ;
        RECT 1974.190 514.000 1977.950 514.280 ;
        RECT 1978.790 514.000 1982.090 514.280 ;
        RECT 1982.930 514.000 1986.230 514.280 ;
        RECT 1987.070 514.000 1990.830 514.280 ;
        RECT 1991.670 514.000 1994.970 514.280 ;
        RECT 1995.810 514.000 1999.110 514.280 ;
        RECT 1999.950 514.000 2003.250 514.280 ;
        RECT 2004.090 514.000 2007.850 514.280 ;
        RECT 2008.690 514.000 2011.990 514.280 ;
        RECT 2012.830 514.000 2016.130 514.280 ;
        RECT 2016.970 514.000 2020.270 514.280 ;
        RECT 2021.110 514.000 2024.870 514.280 ;
        RECT 2025.710 514.000 2029.010 514.280 ;
        RECT 2029.850 514.000 2033.150 514.280 ;
        RECT 2033.990 514.000 2037.750 514.280 ;
        RECT 2038.590 514.000 2041.890 514.280 ;
        RECT 2042.730 514.000 2046.030 514.280 ;
        RECT 2046.870 514.000 2050.170 514.280 ;
        RECT 2051.010 514.000 2054.770 514.280 ;
        RECT 2055.610 514.000 2058.910 514.280 ;
        RECT 2059.750 514.000 2063.050 514.280 ;
        RECT 2063.890 514.000 2067.650 514.280 ;
        RECT 2068.490 514.000 2071.790 514.280 ;
        RECT 2072.630 514.000 2075.930 514.280 ;
        RECT 2076.770 514.000 2080.070 514.280 ;
        RECT 2080.910 514.000 2084.670 514.280 ;
        RECT 2085.510 514.000 2088.810 514.280 ;
        RECT 2089.650 514.000 2092.950 514.280 ;
        RECT 2093.790 514.000 2097.090 514.280 ;
        RECT 2097.930 514.000 2101.690 514.280 ;
        RECT 2102.530 514.000 2105.830 514.280 ;
        RECT 2106.670 514.000 2109.970 514.280 ;
        RECT 2110.810 514.000 2114.570 514.280 ;
        RECT 2115.410 514.000 2118.710 514.280 ;
        RECT 2119.550 514.000 2122.850 514.280 ;
        RECT 2123.690 514.000 2126.990 514.280 ;
        RECT 2127.830 514.000 2131.590 514.280 ;
        RECT 2132.430 514.000 2135.730 514.280 ;
        RECT 2136.570 514.000 2139.870 514.280 ;
        RECT 2140.710 514.000 2144.470 514.280 ;
        RECT 2145.310 514.000 2148.610 514.280 ;
        RECT 2149.450 514.000 2152.750 514.280 ;
        RECT 2153.590 514.000 2156.890 514.280 ;
        RECT 2157.730 514.000 2161.490 514.280 ;
        RECT 2162.330 514.000 2165.630 514.280 ;
        RECT 2166.470 514.000 2169.770 514.280 ;
        RECT 2170.610 514.000 2174.370 514.280 ;
        RECT 2175.210 514.000 2178.510 514.280 ;
        RECT 2179.350 514.000 2182.650 514.280 ;
        RECT 2183.490 514.000 2186.790 514.280 ;
        RECT 2187.630 514.000 2191.390 514.280 ;
        RECT 2192.230 514.000 2195.530 514.280 ;
        RECT 2196.370 514.000 2199.670 514.280 ;
        RECT 2200.510 514.000 2203.810 514.280 ;
        RECT 2204.650 514.000 2208.410 514.280 ;
        RECT 2209.250 514.000 2212.550 514.280 ;
        RECT 2213.390 514.000 2216.690 514.280 ;
        RECT 2217.530 514.000 2221.290 514.280 ;
        RECT 2222.130 514.000 2225.430 514.280 ;
        RECT 2226.270 514.000 2229.570 514.280 ;
        RECT 2230.410 514.000 2233.710 514.280 ;
        RECT 2234.550 514.000 2238.310 514.280 ;
        RECT 2239.150 514.000 2242.450 514.280 ;
        RECT 2243.290 514.000 2246.590 514.280 ;
        RECT 2247.430 514.000 2251.190 514.280 ;
        RECT 2252.030 514.000 2255.330 514.280 ;
        RECT 2256.170 514.000 2259.470 514.280 ;
        RECT 2260.310 514.000 2263.610 514.280 ;
        RECT 2264.450 514.000 2268.210 514.280 ;
        RECT 2269.050 514.000 2272.350 514.280 ;
        RECT 2273.190 514.000 2276.490 514.280 ;
        RECT 2277.330 514.000 2280.630 514.280 ;
        RECT 2281.470 514.000 2285.230 514.280 ;
        RECT 2286.070 514.000 2289.370 514.280 ;
        RECT 2290.210 514.000 2293.510 514.280 ;
        RECT 2294.350 514.000 2298.110 514.280 ;
        RECT 2298.950 514.000 2302.250 514.280 ;
        RECT 2303.090 514.000 2306.390 514.280 ;
        RECT 2307.230 514.000 2310.530 514.280 ;
        RECT 2311.370 514.000 2315.130 514.280 ;
        RECT 2315.970 514.000 2319.270 514.280 ;
        RECT 2320.110 514.000 2323.410 514.280 ;
        RECT 2324.250 514.000 2328.010 514.280 ;
        RECT 2328.850 514.000 2332.150 514.280 ;
        RECT 2332.990 514.000 2336.290 514.280 ;
        RECT 2337.130 514.000 2340.430 514.280 ;
        RECT 2341.270 514.000 2345.030 514.280 ;
        RECT 2345.870 514.000 2349.170 514.280 ;
        RECT 2350.010 514.000 2353.310 514.280 ;
        RECT 2354.150 514.000 2357.450 514.280 ;
        RECT 2358.290 514.000 2362.050 514.280 ;
        RECT 2362.890 514.000 2366.190 514.280 ;
        RECT 2367.030 514.000 2370.330 514.280 ;
        RECT 2371.170 514.000 2374.930 514.280 ;
        RECT 2375.770 514.000 2379.070 514.280 ;
        RECT 2379.910 514.000 2383.210 514.280 ;
        RECT 2384.050 514.000 2387.350 514.280 ;
        RECT 2388.190 514.000 2391.950 514.280 ;
        RECT 2392.790 514.000 2396.090 514.280 ;
        RECT 2396.930 514.000 2400.230 514.280 ;
        RECT 2401.070 514.000 2404.830 514.280 ;
        RECT 2405.670 514.000 2408.970 514.280 ;
        RECT 2409.810 514.000 2413.110 514.280 ;
        RECT 2413.950 514.000 2417.250 514.280 ;
        RECT 2418.090 514.000 2421.850 514.280 ;
        RECT 2422.690 514.000 2425.990 514.280 ;
        RECT 2426.830 514.000 2430.130 514.280 ;
        RECT 2430.970 514.000 2434.270 514.280 ;
        RECT 2435.110 514.000 2438.870 514.280 ;
        RECT 2439.710 514.000 2443.010 514.280 ;
        RECT 2443.850 514.000 2447.150 514.280 ;
        RECT 2447.990 514.000 2451.750 514.280 ;
        RECT 2452.590 514.000 2455.890 514.280 ;
        RECT 2456.730 514.000 2460.030 514.280 ;
        RECT 2460.870 514.000 2464.170 514.280 ;
        RECT 2465.010 514.000 2468.770 514.280 ;
        RECT 2469.610 514.000 2472.910 514.280 ;
        RECT 2473.750 514.000 2477.050 514.280 ;
        RECT 2477.890 514.000 2481.650 514.280 ;
        RECT 2482.490 514.000 2485.790 514.280 ;
        RECT 2486.630 514.000 2489.930 514.280 ;
        RECT 2490.770 514.000 2494.070 514.280 ;
        RECT 2494.910 514.000 2498.670 514.280 ;
      LAYER met2 ;
        RECT 2503.090 510.000 2503.370 514.000 ;
        RECT 2507.230 510.000 2507.510 514.000 ;
      LAYER met3 ;
        RECT 414.000 2982.840 2506.000 2998.965 ;
        RECT 414.000 2981.440 2505.600 2982.840 ;
      LAYER met3 ;
        RECT 2506.000 2981.840 2510.000 2982.440 ;
      LAYER met3 ;
        RECT 414.000 2980.800 2506.000 2981.440 ;
        RECT 414.400 2979.400 2506.000 2980.800 ;
        RECT 414.000 2928.440 2506.000 2979.400 ;
        RECT 414.000 2927.040 2505.600 2928.440 ;
        RECT 414.000 2923.000 2506.000 2927.040 ;
        RECT 414.400 2921.600 2506.000 2923.000 ;
        RECT 414.000 2874.040 2506.000 2921.600 ;
        RECT 414.000 2872.640 2505.600 2874.040 ;
        RECT 414.000 2864.520 2506.000 2872.640 ;
        RECT 414.400 2863.120 2506.000 2864.520 ;
        RECT 414.000 2819.640 2506.000 2863.120 ;
        RECT 414.000 2818.240 2505.600 2819.640 ;
        RECT 414.000 2806.720 2506.000 2818.240 ;
        RECT 414.400 2805.320 2506.000 2806.720 ;
        RECT 414.000 2765.240 2506.000 2805.320 ;
        RECT 414.000 2763.840 2505.600 2765.240 ;
        RECT 414.000 2748.240 2506.000 2763.840 ;
        RECT 414.400 2746.840 2506.000 2748.240 ;
        RECT 414.000 2710.840 2506.000 2746.840 ;
        RECT 414.000 2709.440 2505.600 2710.840 ;
        RECT 414.000 2690.440 2506.000 2709.440 ;
        RECT 414.400 2689.040 2506.000 2690.440 ;
        RECT 414.000 2656.440 2506.000 2689.040 ;
        RECT 414.000 2655.040 2505.600 2656.440 ;
        RECT 414.000 2631.960 2506.000 2655.040 ;
        RECT 414.400 2630.560 2506.000 2631.960 ;
        RECT 414.000 2602.040 2506.000 2630.560 ;
        RECT 414.000 2600.640 2505.600 2602.040 ;
        RECT 414.000 2574.160 2506.000 2600.640 ;
        RECT 414.400 2572.760 2506.000 2574.160 ;
        RECT 414.000 2547.640 2506.000 2572.760 ;
        RECT 414.000 2546.240 2505.600 2547.640 ;
        RECT 414.000 2515.680 2506.000 2546.240 ;
        RECT 414.400 2514.280 2506.000 2515.680 ;
        RECT 414.000 2493.240 2506.000 2514.280 ;
        RECT 414.000 2491.840 2505.600 2493.240 ;
        RECT 414.000 2457.880 2506.000 2491.840 ;
        RECT 414.400 2456.480 2506.000 2457.880 ;
        RECT 414.000 2438.840 2506.000 2456.480 ;
        RECT 414.000 2437.440 2505.600 2438.840 ;
        RECT 414.000 2399.400 2506.000 2437.440 ;
        RECT 414.400 2398.000 2506.000 2399.400 ;
        RECT 414.000 2385.120 2506.000 2398.000 ;
        RECT 414.000 2383.720 2505.600 2385.120 ;
        RECT 414.000 2341.600 2506.000 2383.720 ;
        RECT 414.400 2340.200 2506.000 2341.600 ;
        RECT 414.000 2330.720 2506.000 2340.200 ;
        RECT 414.000 2329.320 2505.600 2330.720 ;
        RECT 414.000 2283.120 2506.000 2329.320 ;
        RECT 414.400 2281.720 2506.000 2283.120 ;
        RECT 414.000 2276.320 2506.000 2281.720 ;
        RECT 414.000 2274.920 2505.600 2276.320 ;
        RECT 414.000 2225.320 2506.000 2274.920 ;
        RECT 414.400 2223.920 2506.000 2225.320 ;
        RECT 414.000 2221.920 2506.000 2223.920 ;
        RECT 414.000 2220.520 2505.600 2221.920 ;
        RECT 414.000 2167.520 2506.000 2220.520 ;
        RECT 414.000 2166.840 2505.600 2167.520 ;
        RECT 414.400 2166.120 2505.600 2166.840 ;
        RECT 414.400 2165.440 2506.000 2166.120 ;
        RECT 414.000 2113.120 2506.000 2165.440 ;
        RECT 414.000 2111.720 2505.600 2113.120 ;
        RECT 414.000 2109.040 2506.000 2111.720 ;
        RECT 414.400 2107.640 2506.000 2109.040 ;
        RECT 414.000 2058.720 2506.000 2107.640 ;
        RECT 414.000 2057.320 2505.600 2058.720 ;
        RECT 414.000 2050.560 2506.000 2057.320 ;
        RECT 414.400 2049.160 2506.000 2050.560 ;
        RECT 414.000 2004.320 2506.000 2049.160 ;
        RECT 414.000 2002.920 2505.600 2004.320 ;
        RECT 414.000 1992.760 2506.000 2002.920 ;
        RECT 414.400 1991.360 2506.000 1992.760 ;
        RECT 414.000 1949.920 2506.000 1991.360 ;
        RECT 414.000 1948.520 2505.600 1949.920 ;
        RECT 414.000 1934.280 2506.000 1948.520 ;
        RECT 414.400 1932.880 2506.000 1934.280 ;
        RECT 414.000 1895.520 2506.000 1932.880 ;
        RECT 414.000 1894.120 2505.600 1895.520 ;
        RECT 414.000 1876.480 2506.000 1894.120 ;
        RECT 414.400 1875.080 2506.000 1876.480 ;
        RECT 414.000 1841.120 2506.000 1875.080 ;
        RECT 414.000 1839.720 2505.600 1841.120 ;
        RECT 414.000 1818.000 2506.000 1839.720 ;
        RECT 414.400 1816.600 2506.000 1818.000 ;
        RECT 414.000 1787.400 2506.000 1816.600 ;
        RECT 414.000 1786.000 2505.600 1787.400 ;
        RECT 414.000 1760.200 2506.000 1786.000 ;
        RECT 414.400 1758.800 2506.000 1760.200 ;
        RECT 414.000 1733.000 2506.000 1758.800 ;
        RECT 414.000 1731.600 2505.600 1733.000 ;
        RECT 414.000 1701.720 2506.000 1731.600 ;
        RECT 414.400 1700.320 2506.000 1701.720 ;
        RECT 414.000 1678.600 2506.000 1700.320 ;
        RECT 414.000 1677.200 2505.600 1678.600 ;
        RECT 414.000 1643.920 2506.000 1677.200 ;
        RECT 414.400 1642.520 2506.000 1643.920 ;
        RECT 414.000 1624.200 2506.000 1642.520 ;
        RECT 414.000 1622.800 2505.600 1624.200 ;
        RECT 414.000 1585.440 2506.000 1622.800 ;
        RECT 414.400 1584.040 2506.000 1585.440 ;
        RECT 414.000 1569.800 2506.000 1584.040 ;
        RECT 414.000 1568.400 2505.600 1569.800 ;
        RECT 414.000 1527.640 2506.000 1568.400 ;
        RECT 414.400 1526.240 2506.000 1527.640 ;
        RECT 414.000 1515.400 2506.000 1526.240 ;
        RECT 414.000 1514.000 2505.600 1515.400 ;
        RECT 414.000 1469.160 2506.000 1514.000 ;
        RECT 414.400 1467.760 2506.000 1469.160 ;
        RECT 414.000 1461.000 2506.000 1467.760 ;
        RECT 414.000 1459.600 2505.600 1461.000 ;
        RECT 414.000 1411.360 2506.000 1459.600 ;
        RECT 414.400 1409.960 2506.000 1411.360 ;
        RECT 414.000 1406.600 2506.000 1409.960 ;
        RECT 414.000 1405.200 2505.600 1406.600 ;
        RECT 414.000 1352.880 2506.000 1405.200 ;
        RECT 414.400 1352.200 2506.000 1352.880 ;
        RECT 414.400 1351.480 2505.600 1352.200 ;
        RECT 414.000 1350.800 2505.600 1351.480 ;
        RECT 414.000 1297.800 2506.000 1350.800 ;
        RECT 414.000 1296.400 2505.600 1297.800 ;
        RECT 414.000 1295.080 2506.000 1296.400 ;
        RECT 414.400 1293.680 2506.000 1295.080 ;
        RECT 414.000 1243.400 2506.000 1293.680 ;
        RECT 414.000 1242.000 2505.600 1243.400 ;
        RECT 414.000 1236.600 2506.000 1242.000 ;
        RECT 414.400 1235.200 2506.000 1236.600 ;
        RECT 414.000 1189.000 2506.000 1235.200 ;
        RECT 414.000 1187.600 2505.600 1189.000 ;
        RECT 414.000 1178.800 2506.000 1187.600 ;
        RECT 414.400 1177.400 2506.000 1178.800 ;
        RECT 414.000 1135.280 2506.000 1177.400 ;
        RECT 414.000 1133.880 2505.600 1135.280 ;
        RECT 414.000 1120.320 2506.000 1133.880 ;
        RECT 414.400 1118.920 2506.000 1120.320 ;
        RECT 414.000 1080.880 2506.000 1118.920 ;
        RECT 414.000 1079.480 2505.600 1080.880 ;
        RECT 414.000 1062.520 2506.000 1079.480 ;
        RECT 414.400 1061.120 2506.000 1062.520 ;
        RECT 414.000 1026.480 2506.000 1061.120 ;
        RECT 414.000 1025.080 2505.600 1026.480 ;
        RECT 414.000 1004.040 2506.000 1025.080 ;
        RECT 414.400 1002.640 2506.000 1004.040 ;
        RECT 414.000 972.080 2506.000 1002.640 ;
        RECT 414.000 970.680 2505.600 972.080 ;
        RECT 414.000 946.240 2506.000 970.680 ;
        RECT 414.400 944.840 2506.000 946.240 ;
        RECT 414.000 917.680 2506.000 944.840 ;
        RECT 414.000 916.280 2505.600 917.680 ;
        RECT 414.000 887.760 2506.000 916.280 ;
        RECT 414.400 886.360 2506.000 887.760 ;
        RECT 414.000 863.280 2506.000 886.360 ;
        RECT 414.000 861.880 2505.600 863.280 ;
        RECT 414.000 829.960 2506.000 861.880 ;
        RECT 414.400 828.560 2506.000 829.960 ;
        RECT 414.000 808.880 2506.000 828.560 ;
        RECT 414.000 807.480 2505.600 808.880 ;
        RECT 414.000 771.480 2506.000 807.480 ;
        RECT 414.400 770.080 2506.000 771.480 ;
        RECT 414.000 754.480 2506.000 770.080 ;
        RECT 414.000 753.080 2505.600 754.480 ;
        RECT 414.000 713.680 2506.000 753.080 ;
        RECT 414.400 712.280 2506.000 713.680 ;
        RECT 414.000 700.080 2506.000 712.280 ;
        RECT 414.000 698.680 2505.600 700.080 ;
        RECT 414.000 655.200 2506.000 698.680 ;
        RECT 414.400 653.800 2506.000 655.200 ;
        RECT 414.000 645.680 2506.000 653.800 ;
        RECT 414.000 644.280 2505.600 645.680 ;
        RECT 414.000 597.400 2506.000 644.280 ;
        RECT 414.400 596.000 2506.000 597.400 ;
        RECT 414.000 591.280 2506.000 596.000 ;
        RECT 414.000 589.880 2505.600 591.280 ;
        RECT 414.000 539.600 2506.000 589.880 ;
      LAYER met3 ;
        RECT 410.000 538.600 414.000 539.200 ;
      LAYER met3 ;
        RECT 414.400 538.200 2506.000 539.600 ;
        RECT 414.000 537.560 2506.000 538.200 ;
        RECT 414.000 536.160 2505.600 537.560 ;
        RECT 414.000 520.715 2506.000 536.160 ;
      LAYER met4 ;
        RECT 431.040 520.640 432.640 2999.040 ;
        RECT 507.840 520.640 509.440 2999.040 ;
      LAYER met4 ;
        RECT 584.640 520.640 2429.440 2999.040 ;
  END
END user_project_wrapper
END LIBRARY

