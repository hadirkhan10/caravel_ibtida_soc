magic
tech sky130A
magscale 1 2
timestamp 1607298761
<< checkpaint >>
rect -9696 -8626 593620 712562
<< locali >>
rect 412649 683247 412683 692733
rect 413017 666587 413051 683077
rect 412833 601715 412867 608549
rect 412925 589339 412959 598893
rect 89729 584103 89763 584749
rect 96445 584035 96479 584749
rect 498117 584443 498151 584613
rect 500233 584239 500267 584409
rect 106473 583695 106507 584069
rect 124137 583695 124171 584069
rect 500325 583763 500359 584205
rect 99941 582335 99975 582573
rect 134349 581247 134383 581621
rect 144377 581247 144411 581621
rect 524429 550647 524463 568497
rect 82829 520319 82863 529873
rect 82829 491351 82863 500905
rect 524429 462451 524463 471937
rect 82737 438175 82771 442901
rect 82829 439535 82863 447797
rect 524429 443003 524463 452557
rect 524429 423691 524463 433245
rect 82829 414035 82863 423589
rect 82921 418999 82955 422977
rect 82737 400231 82771 400673
rect 82829 399551 82863 400333
rect 82921 387991 82955 406249
rect 524429 404379 524463 413933
rect 524429 385067 524463 394621
rect 82829 375479 82863 384965
rect 82277 365279 82311 370821
rect 82921 369359 82955 372589
rect 524429 365755 524463 375309
rect 524429 346443 524463 355997
rect 524429 327131 524463 336685
rect 79609 309859 79643 319073
rect 82921 317475 82955 326961
rect 79517 309825 79643 309859
rect 79517 296123 79551 309825
rect 82737 309111 82771 313293
rect 82737 302923 82771 303297
rect 82829 298299 82863 311321
rect 82921 310607 82955 310845
rect 524429 307819 524463 317373
rect 79333 280823 79367 287317
rect 79793 280823 79827 287317
rect 82737 286399 82771 298061
rect 82829 288847 82863 293369
rect 82921 291907 82955 303025
rect 82921 287759 82955 291737
rect 82921 277423 82955 282217
rect 82645 265455 82679 269569
rect 82737 265863 82771 269433
rect 82829 263551 82863 269773
rect 82921 263143 82955 273785
rect 501797 272391 501831 278409
rect 501889 272663 501923 282217
rect 501981 272527 502015 290241
rect 524429 288439 524463 298061
rect 502073 270895 502107 272765
rect 501521 253215 501555 270385
rect 501613 254643 501647 266985
rect 506213 264843 506247 277865
rect 82645 243695 82679 245905
rect 82737 244987 82771 246177
rect 82829 243559 82863 246313
rect 82921 245055 82955 248421
rect 504649 246415 504683 252977
rect 505845 251311 505879 254813
rect 81449 230639 81483 233665
rect 81541 229279 81575 238085
rect 82645 227919 82679 232577
rect 82737 228871 82771 232985
rect 82829 225675 82863 233053
rect 82921 226559 82955 238697
rect 82921 219487 82955 220813
rect 501521 210783 501555 220201
rect 501613 220031 501647 233597
rect 503637 227443 503671 241553
rect 503545 219691 503579 225505
rect 503637 221255 503671 221493
rect 506213 212211 506247 217957
rect 81541 200175 81575 202453
rect 81541 190519 81575 192389
rect 81633 187255 81667 191777
rect 82093 188615 82127 194769
rect 82185 190791 82219 195041
rect 82277 188411 82311 201773
rect 82645 201263 82679 209457
rect 82369 186983 82403 191233
rect 82461 190995 82495 194905
rect 82553 191199 82587 200277
rect 82553 189091 82587 190825
rect 82553 178619 82587 188921
rect 82645 182427 82679 191097
rect 82737 185691 82771 195245
rect 82829 195143 82863 195313
rect 82955 195177 83047 195211
rect 82829 187119 82863 194905
rect 82921 187051 82955 194769
rect 82829 187017 82955 187051
rect 82829 186779 82863 187017
rect 83013 186983 83047 195177
rect 82955 186949 83047 186983
rect 82955 186813 83047 186847
rect 82829 186745 82955 186779
rect 82921 184195 82955 186745
rect 82829 184161 82955 184195
rect 82829 178755 82863 184161
rect 82829 178721 82955 178755
rect 79609 175559 79643 176545
rect 82645 170255 82679 178721
rect 82737 173179 82771 177089
rect 82829 173179 82863 177225
rect 82921 176987 82955 178721
rect 83013 176647 83047 186813
rect 82955 176613 83047 176647
rect 82829 173145 82955 173179
rect 82737 166719 82771 167229
rect 82829 167127 82863 168385
rect 82921 166039 82955 173145
rect 501521 165631 501555 178177
rect 81541 157199 81575 157437
rect 81633 157335 81667 162129
rect 82645 156247 82679 162809
rect 82737 152167 82771 157573
rect 82829 152371 82863 157505
rect 501521 157471 501555 163761
rect 501613 160803 501647 207825
rect 502165 197727 502199 209321
rect 503545 199359 503579 204833
rect 503637 196231 503671 199461
rect 503085 189703 503119 194361
rect 505937 190791 505971 199597
rect 503637 180183 503671 186949
rect 501613 160769 501831 160803
rect 501705 155091 501739 159069
rect 501797 154887 501831 160769
rect 78781 150331 78815 150977
rect 82829 145503 82863 145877
rect 82921 145775 82955 152473
rect 501521 147271 501555 151793
rect 80161 137071 80195 140369
rect 80437 137207 80471 144041
rect 80989 136527 81023 136833
rect 79609 121499 79643 133297
rect 82645 132311 82679 137173
rect 82737 136935 82771 137309
rect 82829 133059 82863 138465
rect 82921 137071 82955 138669
rect 80437 122723 80471 123437
rect 81909 121499 81943 122689
rect 82093 122383 82127 123641
rect 82461 121771 82495 123573
rect 82093 121091 82127 121737
rect 82829 120615 82863 123641
rect 82921 120479 82955 133161
rect 501521 131087 501555 144449
rect 501613 136187 501647 138057
rect 501613 129591 501647 133297
rect 501705 133195 501739 149005
rect 501889 143667 501923 166345
rect 501981 154751 502015 162129
rect 502901 158695 502935 162401
rect 502993 155431 503027 164917
rect 503637 154615 503671 169201
rect 501521 129557 501647 129591
rect 501521 127143 501555 129557
rect 103529 122043 103563 122757
rect 84117 120615 84151 121737
rect 82461 119255 82495 119357
rect 82737 113203 82771 119425
rect 83473 119255 83507 119357
rect 86325 118099 86359 119561
rect 107577 119255 107611 119561
rect 110429 114563 110463 120513
rect 114569 118847 114603 119221
rect 156061 118643 156095 122553
rect 326997 122043 327031 122757
rect 338129 121703 338163 122485
rect 393973 121975 394007 122077
rect 498209 121873 498427 121907
rect 498209 121839 498243 121873
rect 498301 121703 498335 121805
rect 498243 121669 498335 121703
rect 498393 121635 498427 121873
rect 498485 121669 499405 121703
rect 498301 121567 498335 121601
rect 498485 121567 498519 121669
rect 498301 121533 498519 121567
rect 501521 121431 501555 124729
rect 501613 123335 501647 127313
rect 501705 123471 501739 133025
rect 501797 127211 501831 140097
rect 501889 135507 501923 141797
rect 501981 137479 502015 139961
rect 501613 121091 501647 123165
rect 501889 121499 501923 127313
rect 501981 123879 502015 132481
rect 499037 120683 499071 121057
rect 496829 120615 496863 120649
rect 496829 120581 497013 120615
rect 501613 120343 501647 120445
rect 161305 116059 161339 119289
rect 212457 119187 212491 119493
rect 489193 119391 489227 119629
rect 248981 119289 249199 119323
rect 248981 118915 249015 119289
rect 249165 119255 249199 119289
rect 492781 119255 492815 119357
rect 249073 118915 249107 119221
rect 501705 119187 501739 121057
rect 226349 118711 226383 118813
rect 350549 118711 350583 118813
rect 502073 118575 502107 137785
rect 502165 137071 502199 140369
rect 502257 133059 502291 148801
rect 503729 148087 503763 162809
rect 503729 148053 503855 148087
rect 502349 136323 502383 147441
rect 503729 146999 503763 147985
rect 503821 146931 503855 148053
rect 503729 146897 503855 146931
rect 502441 136935 502475 140233
rect 502165 123743 502199 127313
rect 502349 123199 502383 130577
rect 502533 129999 502567 140505
rect 502625 121771 502659 124729
rect 503453 117827 503487 131053
rect 503545 124831 503579 127789
rect 503637 127687 503671 143361
rect 503729 133943 503763 146897
rect 504557 146183 504591 152541
rect 505569 151895 505603 155533
rect 505753 147407 505787 152065
rect 505845 151283 505879 162945
rect 524429 153255 524463 162809
rect 532709 153255 532743 162809
rect 504097 138295 504131 145945
rect 505845 131835 505879 143633
rect 506397 131835 506431 148869
rect 524429 133943 524463 143497
rect 532709 133943 532743 143497
rect 503729 122383 503763 131053
rect 80069 102187 80103 111741
rect 110429 104907 110463 114393
rect 117513 100827 117547 110381
rect 131221 106335 131255 115889
rect 153025 108919 153059 115821
rect 155877 104907 155911 114461
rect 161305 108919 161339 115889
rect 179337 106403 179371 115889
rect 186237 114563 186271 115345
rect 244289 106335 244323 115889
rect 110429 85663 110463 95149
rect 117513 89743 117547 99297
rect 131221 87023 131255 96577
rect 156245 95251 156279 104737
rect 179337 87091 179371 104805
rect 186237 95251 186271 104805
rect 220737 95251 220771 104805
rect 223589 95251 223623 104805
rect 258089 102935 258123 115889
rect 272901 108919 272935 109157
rect 304917 105519 304951 111265
rect 220553 85595 220587 95149
rect 244289 87023 244323 96577
rect 258089 87023 258123 96577
rect 272993 87023 273027 96577
rect 299305 87023 299339 96577
rect 351745 89675 351779 104805
rect 378149 95251 378183 110993
rect 436109 96747 436143 111061
rect 445861 106335 445895 115889
rect 511641 115855 511675 119969
rect 524429 114563 524463 124049
rect 532709 114563 532743 124049
rect 511549 104907 511583 114461
rect 445861 87023 445895 96577
rect 511733 96543 511767 104737
rect 524429 95251 524463 104805
rect 532709 95251 532743 104805
rect 80069 73219 80103 82773
rect 120365 81447 120399 82841
rect 179337 75939 179371 85493
rect 186237 75939 186271 85493
rect 220645 75939 220679 85493
rect 223589 75939 223623 85493
rect 110429 66283 110463 75837
rect 244289 67643 244323 77129
rect 258089 67643 258123 77129
rect 378149 75939 378183 85493
rect 436109 77299 436143 86921
rect 500233 77299 500267 93857
rect 445861 67643 445895 77129
rect 511549 75939 511583 85493
rect 524429 75939 524463 85493
rect 532709 75939 532743 85493
rect 155969 56627 156003 66181
rect 110429 46971 110463 56457
rect 161029 55267 161063 64821
rect 179337 56627 179371 66181
rect 186237 56627 186271 66181
rect 220737 56627 220771 66181
rect 223589 56627 223623 66181
rect 244289 48331 244323 57885
rect 258089 48331 258123 57885
rect 378149 56627 378183 66181
rect 436109 57987 436143 67541
rect 436109 48331 436143 57817
rect 445861 48331 445895 57885
rect 511549 56627 511583 66181
rect 524429 56627 524463 66181
rect 532709 56627 532743 66181
rect 82645 44183 82679 45577
rect 156061 41395 156095 46869
rect 110429 27659 110463 37145
rect 117513 27659 117547 39321
rect 120273 27659 120307 39321
rect 161121 37315 161155 46869
rect 179245 37315 179279 46869
rect 186237 37315 186271 46869
rect 220645 37315 220679 46869
rect 223589 37315 223623 46869
rect 272993 38675 273027 48229
rect 152933 29019 152967 31773
rect 117421 15215 117455 22117
rect 131221 9707 131255 19261
rect 152933 18003 152967 27557
rect 156153 19363 156187 28917
rect 161213 27659 161247 32453
rect 161489 18003 161523 28917
rect 220461 27659 220495 37213
rect 244289 29019 244323 38573
rect 258089 29019 258123 38573
rect 289737 37315 289771 46869
rect 299397 38675 299431 48229
rect 351745 38675 351779 48229
rect 378149 37315 378183 46869
rect 505845 41259 505879 46869
rect 436109 29087 436143 38573
rect 445861 29019 445895 38573
rect 156153 9707 156187 14569
rect 178969 9707 179003 27557
rect 186053 9775 186087 27557
rect 220737 18003 220771 27557
rect 223589 18003 223623 27557
rect 220553 9707 220587 12529
rect 221749 9707 221783 12461
rect 244289 9707 244323 19261
rect 245485 11543 245519 13413
rect 289737 12495 289771 27557
rect 299121 18003 299155 27557
rect 341901 9707 341935 14705
rect 351745 9775 351779 19261
rect 378149 18003 378183 27557
rect 393053 9707 393087 12529
rect 436109 9775 436143 19261
rect 445861 9707 445895 19261
rect 505753 19227 505787 29665
rect 511549 29087 511583 46869
rect 524429 37315 524463 46869
rect 532709 37315 532743 46869
rect 511549 18003 511583 27557
rect 524429 18003 524463 27557
rect 527465 12359 527499 13549
rect 532709 9707 532743 27557
rect 541725 9707 541759 13345
rect 69305 3519 69339 3689
rect 88349 3043 88383 4097
rect 94421 3043 94455 4165
rect 94513 3043 94547 4097
rect 99205 3723 99239 4097
rect 99297 3111 99331 4165
rect 100493 595 100527 9605
rect 109049 2771 109083 3689
rect 111165 595 111199 6817
rect 112269 3723 112303 4165
rect 118341 3723 118375 4165
rect 118743 3077 118835 3111
rect 118801 2975 118835 3077
rect 128219 3009 128403 3043
rect 122849 2771 122883 3009
rect 128369 2975 128403 3009
rect 128277 2907 128311 2941
rect 128461 2907 128495 3009
rect 128277 2873 128495 2907
rect 132417 2771 132451 3077
rect 133889 2839 133923 3077
rect 134901 595 134935 9605
rect 154037 3077 154255 3111
rect 154037 3043 154071 3077
rect 136741 2839 136775 3009
rect 142813 2839 142847 2941
rect 154129 2839 154163 3009
rect 154221 2839 154255 3077
rect 157257 2839 157291 3077
rect 157349 2839 157383 3077
rect 166917 2839 166951 3077
rect 186053 595 186087 9605
rect 208593 3179 208627 3825
rect 201509 2839 201543 2941
rect 208501 2907 208535 3145
rect 209513 3111 209547 3349
rect 219541 3111 219575 3349
rect 211077 2839 211111 3009
rect 220093 2907 220127 3145
rect 220829 3043 220863 3145
rect 248981 3043 249015 3213
rect 229109 2907 229143 3009
rect 234905 2907 234939 3009
rect 249073 2975 249107 3349
rect 258641 595 258675 9605
rect 351745 4675 351779 9605
rect 305009 3383 305043 3961
rect 258733 2975 258767 3349
rect 326353 3383 326387 3961
rect 349077 3383 349111 4029
rect 283573 3111 283607 3349
rect 297373 3111 297407 3281
rect 370421 595 370455 9605
rect 371617 595 371651 9605
rect 372813 595 372847 9605
rect 374653 4675 374687 4913
rect 377597 595 377631 9605
rect 378793 595 378827 9605
rect 393973 3111 394007 3621
rect 415593 3111 415627 3621
rect 428749 595 428783 9605
rect 430129 3111 430163 3621
rect 437029 595 437063 9605
rect 490573 2839 490607 3213
rect 490665 2839 490699 3349
rect 494989 2839 495023 4301
rect 498853 3179 498887 3825
rect 500233 3383 500267 3621
rect 503027 3213 503269 3247
rect 496737 2839 496771 3077
rect 499531 2805 499623 2839
rect 499589 2771 499623 2805
<< viali >>
rect 412649 692733 412683 692767
rect 412649 683213 412683 683247
rect 413017 683077 413051 683111
rect 413017 666553 413051 666587
rect 412833 608549 412867 608583
rect 412833 601681 412867 601715
rect 412925 598893 412959 598927
rect 412925 589305 412959 589339
rect 89729 584749 89763 584783
rect 89729 584069 89763 584103
rect 96445 584749 96479 584783
rect 498117 584613 498151 584647
rect 498117 584409 498151 584443
rect 500233 584409 500267 584443
rect 500233 584205 500267 584239
rect 500325 584205 500359 584239
rect 96445 584001 96479 584035
rect 106473 584069 106507 584103
rect 106473 583661 106507 583695
rect 124137 584069 124171 584103
rect 500325 583729 500359 583763
rect 124137 583661 124171 583695
rect 99941 582573 99975 582607
rect 99941 582301 99975 582335
rect 134349 581621 134383 581655
rect 134349 581213 134383 581247
rect 144377 581621 144411 581655
rect 144377 581213 144411 581247
rect 524429 568497 524463 568531
rect 524429 550613 524463 550647
rect 82829 529873 82863 529907
rect 82829 520285 82863 520319
rect 82829 500905 82863 500939
rect 82829 491317 82863 491351
rect 524429 471937 524463 471971
rect 524429 462417 524463 462451
rect 524429 452557 524463 452591
rect 82829 447797 82863 447831
rect 82737 442901 82771 442935
rect 524429 442969 524463 443003
rect 82829 439501 82863 439535
rect 82737 438141 82771 438175
rect 524429 433245 524463 433279
rect 524429 423657 524463 423691
rect 82829 423589 82863 423623
rect 82921 422977 82955 423011
rect 82921 418965 82955 418999
rect 82829 414001 82863 414035
rect 524429 413933 524463 413967
rect 82921 406249 82955 406283
rect 82737 400673 82771 400707
rect 82737 400197 82771 400231
rect 82829 400333 82863 400367
rect 82829 399517 82863 399551
rect 524429 404345 524463 404379
rect 82921 387957 82955 387991
rect 524429 394621 524463 394655
rect 524429 385033 524463 385067
rect 82829 384965 82863 384999
rect 82829 375445 82863 375479
rect 524429 375309 524463 375343
rect 82921 372589 82955 372623
rect 82277 370821 82311 370855
rect 82921 369325 82955 369359
rect 524429 365721 524463 365755
rect 82277 365245 82311 365279
rect 524429 355997 524463 356031
rect 524429 346409 524463 346443
rect 524429 336685 524463 336719
rect 524429 327097 524463 327131
rect 82921 326961 82955 326995
rect 79609 319073 79643 319107
rect 82921 317441 82955 317475
rect 524429 317373 524463 317407
rect 82737 313293 82771 313327
rect 82737 309077 82771 309111
rect 82829 311321 82863 311355
rect 82737 303297 82771 303331
rect 82737 302889 82771 302923
rect 82921 310845 82955 310879
rect 82921 310573 82955 310607
rect 524429 307785 524463 307819
rect 82829 298265 82863 298299
rect 82921 303025 82955 303059
rect 79517 296089 79551 296123
rect 82737 298061 82771 298095
rect 79333 287317 79367 287351
rect 79333 280789 79367 280823
rect 79793 287317 79827 287351
rect 82829 293369 82863 293403
rect 82921 291873 82955 291907
rect 524429 298061 524463 298095
rect 82829 288813 82863 288847
rect 82921 291737 82955 291771
rect 82921 287725 82955 287759
rect 501981 290241 502015 290275
rect 82737 286365 82771 286399
rect 79793 280789 79827 280823
rect 82921 282217 82955 282251
rect 501889 282217 501923 282251
rect 82921 277389 82955 277423
rect 501797 278409 501831 278443
rect 82921 273785 82955 273819
rect 82829 269773 82863 269807
rect 82645 269569 82679 269603
rect 82737 269433 82771 269467
rect 82737 265829 82771 265863
rect 82645 265421 82679 265455
rect 82829 263517 82863 263551
rect 501889 272629 501923 272663
rect 524429 288405 524463 288439
rect 506213 277865 506247 277899
rect 501981 272493 502015 272527
rect 502073 272765 502107 272799
rect 501797 272357 501831 272391
rect 502073 270861 502107 270895
rect 82921 263109 82955 263143
rect 501521 270385 501555 270419
rect 501613 266985 501647 267019
rect 506213 264809 506247 264843
rect 501613 254609 501647 254643
rect 505845 254813 505879 254847
rect 501521 253181 501555 253215
rect 504649 252977 504683 253011
rect 82921 248421 82955 248455
rect 82829 246313 82863 246347
rect 82737 246177 82771 246211
rect 82645 245905 82679 245939
rect 82737 244953 82771 244987
rect 82645 243661 82679 243695
rect 505845 251277 505879 251311
rect 504649 246381 504683 246415
rect 82921 245021 82955 245055
rect 82829 243525 82863 243559
rect 503637 241553 503671 241587
rect 82921 238697 82955 238731
rect 81541 238085 81575 238119
rect 81449 233665 81483 233699
rect 81449 230605 81483 230639
rect 82829 233053 82863 233087
rect 82737 232985 82771 233019
rect 81541 229245 81575 229279
rect 82645 232577 82679 232611
rect 82737 228837 82771 228871
rect 82645 227885 82679 227919
rect 82921 226525 82955 226559
rect 501613 233597 501647 233631
rect 82829 225641 82863 225675
rect 82921 220813 82955 220847
rect 82921 219453 82955 219487
rect 501521 220201 501555 220235
rect 503637 227409 503671 227443
rect 501613 219997 501647 220031
rect 503545 225505 503579 225539
rect 503637 221493 503671 221527
rect 503637 221221 503671 221255
rect 503545 219657 503579 219691
rect 506213 217957 506247 217991
rect 506213 212177 506247 212211
rect 501521 210749 501555 210783
rect 82645 209457 82679 209491
rect 81541 202453 81575 202487
rect 81541 200141 81575 200175
rect 82277 201773 82311 201807
rect 82185 195041 82219 195075
rect 82093 194769 82127 194803
rect 81541 192389 81575 192423
rect 81541 190485 81575 190519
rect 81633 191777 81667 191811
rect 82185 190757 82219 190791
rect 82093 188581 82127 188615
rect 502165 209321 502199 209355
rect 82645 201229 82679 201263
rect 501613 207825 501647 207859
rect 82553 200277 82587 200311
rect 82461 194905 82495 194939
rect 82277 188377 82311 188411
rect 82369 191233 82403 191267
rect 81633 187221 81667 187255
rect 82829 195313 82863 195347
rect 82553 191165 82587 191199
rect 82737 195245 82771 195279
rect 82461 190961 82495 190995
rect 82645 191097 82679 191131
rect 82553 190825 82587 190859
rect 82553 189057 82587 189091
rect 82369 186949 82403 186983
rect 82553 188921 82587 188955
rect 82921 195177 82955 195211
rect 82829 195109 82863 195143
rect 82829 194905 82863 194939
rect 82829 187085 82863 187119
rect 82921 194769 82955 194803
rect 82921 186949 82955 186983
rect 82921 186813 82955 186847
rect 82737 185657 82771 185691
rect 82645 182393 82679 182427
rect 82553 178585 82587 178619
rect 82645 178721 82679 178755
rect 79609 176545 79643 176579
rect 79609 175525 79643 175559
rect 82829 177225 82863 177259
rect 82737 177089 82771 177123
rect 82737 173145 82771 173179
rect 82921 176953 82955 176987
rect 82921 176613 82955 176647
rect 501521 178177 501555 178211
rect 82645 170221 82679 170255
rect 82829 168385 82863 168419
rect 82737 167229 82771 167263
rect 82829 167093 82863 167127
rect 82737 166685 82771 166719
rect 82921 166005 82955 166039
rect 501521 165597 501555 165631
rect 501521 163761 501555 163795
rect 82645 162809 82679 162843
rect 81633 162129 81667 162163
rect 81541 157437 81575 157471
rect 81633 157301 81667 157335
rect 81541 157165 81575 157199
rect 82645 156213 82679 156247
rect 82737 157573 82771 157607
rect 82829 157505 82863 157539
rect 503545 204833 503579 204867
rect 505937 199597 505971 199631
rect 503545 199325 503579 199359
rect 503637 199461 503671 199495
rect 502165 197693 502199 197727
rect 503637 196197 503671 196231
rect 503085 194361 503119 194395
rect 505937 190757 505971 190791
rect 503085 189669 503119 189703
rect 503637 186949 503671 186983
rect 503637 180149 503671 180183
rect 503637 169201 503671 169235
rect 501889 166345 501923 166379
rect 501521 157437 501555 157471
rect 501705 159069 501739 159103
rect 501705 155057 501739 155091
rect 501797 154853 501831 154887
rect 82829 152337 82863 152371
rect 82921 152473 82955 152507
rect 82737 152133 82771 152167
rect 78781 150977 78815 151011
rect 78781 150297 78815 150331
rect 82829 145877 82863 145911
rect 501521 151793 501555 151827
rect 501521 147237 501555 147271
rect 501705 149005 501739 149039
rect 82921 145741 82955 145775
rect 82829 145469 82863 145503
rect 501521 144449 501555 144483
rect 80437 144041 80471 144075
rect 80161 140369 80195 140403
rect 82921 138669 82955 138703
rect 82829 138465 82863 138499
rect 82737 137309 82771 137343
rect 80437 137173 80471 137207
rect 82645 137173 82679 137207
rect 80161 137037 80195 137071
rect 80989 136833 81023 136867
rect 80989 136493 81023 136527
rect 79609 133297 79643 133331
rect 82737 136901 82771 136935
rect 82921 137037 82955 137071
rect 82829 133025 82863 133059
rect 82921 133161 82955 133195
rect 82645 132277 82679 132311
rect 82093 123641 82127 123675
rect 80437 123437 80471 123471
rect 80437 122689 80471 122723
rect 81909 122689 81943 122723
rect 79609 121465 79643 121499
rect 82829 123641 82863 123675
rect 82093 122349 82127 122383
rect 82461 123573 82495 123607
rect 81909 121465 81943 121499
rect 82093 121737 82127 121771
rect 82461 121737 82495 121771
rect 82093 121057 82127 121091
rect 82829 120581 82863 120615
rect 501613 138057 501647 138091
rect 501613 136153 501647 136187
rect 501521 131053 501555 131087
rect 501613 133297 501647 133331
rect 502993 164917 503027 164951
rect 502901 162401 502935 162435
rect 501981 162129 502015 162163
rect 502901 158661 502935 158695
rect 502993 155397 503027 155431
rect 501981 154717 502015 154751
rect 505845 162945 505879 162979
rect 503637 154581 503671 154615
rect 503729 162809 503763 162843
rect 501889 143633 501923 143667
rect 502257 148801 502291 148835
rect 501889 141797 501923 141831
rect 501705 133161 501739 133195
rect 501797 140097 501831 140131
rect 501705 133025 501739 133059
rect 501521 127109 501555 127143
rect 501613 127313 501647 127347
rect 501521 124729 501555 124763
rect 103529 122757 103563 122791
rect 326997 122757 327031 122791
rect 103529 122009 103563 122043
rect 156061 122553 156095 122587
rect 84117 121737 84151 121771
rect 84117 120581 84151 120615
rect 82921 120445 82955 120479
rect 110429 120513 110463 120547
rect 86325 119561 86359 119595
rect 82737 119425 82771 119459
rect 82461 119357 82495 119391
rect 82461 119221 82495 119255
rect 83473 119357 83507 119391
rect 83473 119221 83507 119255
rect 107577 119561 107611 119595
rect 107577 119221 107611 119255
rect 86325 118065 86359 118099
rect 114569 119221 114603 119255
rect 114569 118813 114603 118847
rect 326997 122009 327031 122043
rect 338129 122485 338163 122519
rect 393973 122077 394007 122111
rect 393973 121941 394007 121975
rect 498209 121805 498243 121839
rect 498301 121805 498335 121839
rect 338129 121669 338163 121703
rect 498209 121669 498243 121703
rect 498301 121601 498335 121635
rect 498393 121601 498427 121635
rect 499405 121669 499439 121703
rect 502165 140369 502199 140403
rect 501981 139961 502015 139995
rect 501981 137445 502015 137479
rect 502073 137785 502107 137819
rect 501889 135473 501923 135507
rect 501981 132481 502015 132515
rect 501797 127177 501831 127211
rect 501889 127313 501923 127347
rect 501705 123437 501739 123471
rect 501613 123301 501647 123335
rect 501521 121397 501555 121431
rect 501613 123165 501647 123199
rect 501981 123845 502015 123879
rect 501889 121465 501923 121499
rect 499037 121057 499071 121091
rect 501613 121057 501647 121091
rect 501705 121057 501739 121091
rect 496829 120649 496863 120683
rect 499037 120649 499071 120683
rect 497013 120581 497047 120615
rect 501613 120445 501647 120479
rect 501613 120309 501647 120343
rect 489193 119629 489227 119663
rect 212457 119493 212491 119527
rect 156061 118609 156095 118643
rect 161305 119289 161339 119323
rect 489193 119357 489227 119391
rect 492781 119357 492815 119391
rect 212457 119153 212491 119187
rect 248981 118881 249015 118915
rect 249073 119221 249107 119255
rect 249165 119221 249199 119255
rect 492781 119221 492815 119255
rect 501705 119153 501739 119187
rect 249073 118881 249107 118915
rect 226349 118813 226383 118847
rect 226349 118677 226383 118711
rect 350549 118813 350583 118847
rect 350549 118677 350583 118711
rect 502165 137037 502199 137071
rect 505569 155533 505603 155567
rect 504557 152541 504591 152575
rect 503729 147985 503763 148019
rect 502349 147441 502383 147475
rect 503729 146965 503763 146999
rect 503637 143361 503671 143395
rect 502533 140505 502567 140539
rect 502441 140233 502475 140267
rect 502441 136901 502475 136935
rect 502349 136289 502383 136323
rect 502257 133025 502291 133059
rect 502349 130577 502383 130611
rect 502165 127313 502199 127347
rect 502165 123709 502199 123743
rect 502533 129965 502567 129999
rect 503453 131053 503487 131087
rect 502349 123165 502383 123199
rect 502625 124729 502659 124763
rect 502625 121737 502659 121771
rect 502073 118541 502107 118575
rect 503545 127789 503579 127823
rect 505569 151861 505603 151895
rect 505753 152065 505787 152099
rect 524429 162809 524463 162843
rect 524429 153221 524463 153255
rect 532709 162809 532743 162843
rect 532709 153221 532743 153255
rect 505845 151249 505879 151283
rect 505753 147373 505787 147407
rect 506397 148869 506431 148903
rect 504557 146149 504591 146183
rect 504097 145945 504131 145979
rect 504097 138261 504131 138295
rect 505845 143633 505879 143667
rect 503729 133909 503763 133943
rect 505845 131801 505879 131835
rect 524429 143497 524463 143531
rect 524429 133909 524463 133943
rect 532709 143497 532743 143531
rect 532709 133909 532743 133943
rect 506397 131801 506431 131835
rect 503637 127653 503671 127687
rect 503729 131053 503763 131087
rect 503545 124797 503579 124831
rect 503729 122349 503763 122383
rect 524429 124049 524463 124083
rect 503453 117793 503487 117827
rect 511641 119969 511675 120003
rect 161305 116025 161339 116059
rect 110429 114529 110463 114563
rect 131221 115889 131255 115923
rect 82737 113169 82771 113203
rect 110429 114393 110463 114427
rect 80069 111741 80103 111775
rect 110429 104873 110463 104907
rect 117513 110381 117547 110415
rect 80069 102153 80103 102187
rect 161305 115889 161339 115923
rect 153025 115821 153059 115855
rect 153025 108885 153059 108919
rect 155877 114461 155911 114495
rect 131221 106301 131255 106335
rect 161305 108885 161339 108919
rect 179337 115889 179371 115923
rect 244289 115889 244323 115923
rect 186237 115345 186271 115379
rect 186237 114529 186271 114563
rect 179337 106369 179371 106403
rect 244289 106301 244323 106335
rect 258089 115889 258123 115923
rect 155877 104873 155911 104907
rect 179337 104805 179371 104839
rect 117513 100793 117547 100827
rect 156245 104737 156279 104771
rect 117513 99297 117547 99331
rect 110429 95149 110463 95183
rect 117513 89709 117547 89743
rect 131221 96577 131255 96611
rect 156245 95217 156279 95251
rect 186237 104805 186271 104839
rect 186237 95217 186271 95251
rect 220737 104805 220771 104839
rect 220737 95217 220771 95251
rect 223589 104805 223623 104839
rect 445861 115889 445895 115923
rect 304917 111265 304951 111299
rect 272901 109157 272935 109191
rect 272901 108885 272935 108919
rect 436109 111061 436143 111095
rect 304917 105485 304951 105519
rect 378149 110993 378183 111027
rect 258089 102901 258123 102935
rect 351745 104805 351779 104839
rect 223589 95217 223623 95251
rect 244289 96577 244323 96611
rect 179337 87057 179371 87091
rect 220553 95149 220587 95183
rect 131221 86989 131255 87023
rect 110429 85629 110463 85663
rect 244289 86989 244323 87023
rect 258089 96577 258123 96611
rect 258089 86989 258123 87023
rect 272993 96577 273027 96611
rect 272993 86989 273027 87023
rect 299305 96577 299339 96611
rect 511641 115821 511675 115855
rect 524429 114529 524463 114563
rect 532709 124049 532743 124083
rect 532709 114529 532743 114563
rect 445861 106301 445895 106335
rect 511549 114461 511583 114495
rect 511549 104873 511583 104907
rect 524429 104805 524463 104839
rect 436109 96713 436143 96747
rect 511733 104737 511767 104771
rect 378149 95217 378183 95251
rect 445861 96577 445895 96611
rect 351745 89641 351779 89675
rect 299305 86989 299339 87023
rect 511733 96509 511767 96543
rect 524429 95217 524463 95251
rect 532709 104805 532743 104839
rect 532709 95217 532743 95251
rect 445861 86989 445895 87023
rect 500233 93857 500267 93891
rect 220553 85561 220587 85595
rect 436109 86921 436143 86955
rect 179337 85493 179371 85527
rect 120365 82841 120399 82875
rect 80069 82773 80103 82807
rect 120365 81413 120399 81447
rect 179337 75905 179371 75939
rect 186237 85493 186271 85527
rect 186237 75905 186271 75939
rect 220645 85493 220679 85527
rect 220645 75905 220679 75939
rect 223589 85493 223623 85527
rect 378149 85493 378183 85527
rect 223589 75905 223623 75939
rect 244289 77129 244323 77163
rect 80069 73185 80103 73219
rect 110429 75837 110463 75871
rect 244289 67609 244323 67643
rect 258089 77129 258123 77163
rect 436109 77265 436143 77299
rect 500233 77265 500267 77299
rect 511549 85493 511583 85527
rect 378149 75905 378183 75939
rect 445861 77129 445895 77163
rect 258089 67609 258123 67643
rect 511549 75905 511583 75939
rect 524429 85493 524463 85527
rect 524429 75905 524463 75939
rect 532709 85493 532743 85527
rect 532709 75905 532743 75939
rect 445861 67609 445895 67643
rect 110429 66249 110463 66283
rect 436109 67541 436143 67575
rect 155969 66181 156003 66215
rect 179337 66181 179371 66215
rect 155969 56593 156003 56627
rect 161029 64821 161063 64855
rect 110429 56457 110463 56491
rect 179337 56593 179371 56627
rect 186237 66181 186271 66215
rect 186237 56593 186271 56627
rect 220737 66181 220771 66215
rect 220737 56593 220771 56627
rect 223589 66181 223623 66215
rect 378149 66181 378183 66215
rect 223589 56593 223623 56627
rect 244289 57885 244323 57919
rect 161029 55233 161063 55267
rect 244289 48297 244323 48331
rect 258089 57885 258123 57919
rect 436109 57953 436143 57987
rect 511549 66181 511583 66215
rect 445861 57885 445895 57919
rect 378149 56593 378183 56627
rect 436109 57817 436143 57851
rect 258089 48297 258123 48331
rect 436109 48297 436143 48331
rect 511549 56593 511583 56627
rect 524429 66181 524463 66215
rect 524429 56593 524463 56627
rect 532709 66181 532743 66215
rect 532709 56593 532743 56627
rect 445861 48297 445895 48331
rect 110429 46937 110463 46971
rect 272993 48229 273027 48263
rect 156061 46869 156095 46903
rect 82645 45577 82679 45611
rect 82645 44149 82679 44183
rect 156061 41361 156095 41395
rect 161121 46869 161155 46903
rect 117513 39321 117547 39355
rect 110429 37145 110463 37179
rect 110429 27625 110463 27659
rect 117513 27625 117547 27659
rect 120273 39321 120307 39355
rect 161121 37281 161155 37315
rect 179245 46869 179279 46903
rect 179245 37281 179279 37315
rect 186237 46869 186271 46903
rect 186237 37281 186271 37315
rect 220645 46869 220679 46903
rect 220645 37281 220679 37315
rect 223589 46869 223623 46903
rect 299397 48229 299431 48263
rect 272993 38641 273027 38675
rect 289737 46869 289771 46903
rect 223589 37281 223623 37315
rect 244289 38573 244323 38607
rect 220461 37213 220495 37247
rect 161213 32453 161247 32487
rect 152933 31773 152967 31807
rect 152933 28985 152967 29019
rect 120273 27625 120307 27659
rect 156153 28917 156187 28951
rect 152933 27557 152967 27591
rect 117421 22117 117455 22151
rect 117421 15181 117455 15215
rect 131221 19261 131255 19295
rect 161213 27625 161247 27659
rect 161489 28917 161523 28951
rect 156153 19329 156187 19363
rect 152933 17969 152967 18003
rect 244289 28985 244323 29019
rect 258089 38573 258123 38607
rect 299397 38641 299431 38675
rect 351745 48229 351779 48263
rect 351745 38641 351779 38675
rect 378149 46869 378183 46903
rect 289737 37281 289771 37315
rect 505845 46869 505879 46903
rect 505845 41225 505879 41259
rect 511549 46869 511583 46903
rect 378149 37281 378183 37315
rect 436109 38573 436143 38607
rect 436109 29053 436143 29087
rect 445861 38573 445895 38607
rect 258089 28985 258123 29019
rect 445861 28985 445895 29019
rect 505753 29665 505787 29699
rect 220461 27625 220495 27659
rect 161489 17969 161523 18003
rect 178969 27557 179003 27591
rect 131221 9673 131255 9707
rect 156153 14569 156187 14603
rect 156153 9673 156187 9707
rect 186053 27557 186087 27591
rect 220737 27557 220771 27591
rect 220737 17969 220771 18003
rect 223589 27557 223623 27591
rect 289737 27557 289771 27591
rect 223589 17969 223623 18003
rect 244289 19261 244323 19295
rect 186053 9741 186087 9775
rect 220553 12529 220587 12563
rect 178969 9673 179003 9707
rect 220553 9673 220587 9707
rect 221749 12461 221783 12495
rect 221749 9673 221783 9707
rect 245485 13413 245519 13447
rect 299121 27557 299155 27591
rect 378149 27557 378183 27591
rect 299121 17969 299155 18003
rect 351745 19261 351779 19295
rect 289737 12461 289771 12495
rect 341901 14705 341935 14739
rect 245485 11509 245519 11543
rect 244289 9673 244323 9707
rect 378149 17969 378183 18003
rect 436109 19261 436143 19295
rect 351745 9741 351779 9775
rect 393053 12529 393087 12563
rect 341901 9673 341935 9707
rect 436109 9741 436143 9775
rect 445861 19261 445895 19295
rect 393053 9673 393087 9707
rect 524429 46869 524463 46903
rect 524429 37281 524463 37315
rect 532709 46869 532743 46903
rect 532709 37281 532743 37315
rect 511549 29053 511583 29087
rect 505753 19193 505787 19227
rect 511549 27557 511583 27591
rect 511549 17969 511583 18003
rect 524429 27557 524463 27591
rect 524429 17969 524463 18003
rect 532709 27557 532743 27591
rect 527465 13549 527499 13583
rect 527465 12325 527499 12359
rect 445861 9673 445895 9707
rect 532709 9673 532743 9707
rect 541725 13345 541759 13379
rect 541725 9673 541759 9707
rect 100493 9605 100527 9639
rect 94421 4165 94455 4199
rect 88349 4097 88383 4131
rect 69305 3689 69339 3723
rect 69305 3485 69339 3519
rect 88349 3009 88383 3043
rect 99297 4165 99331 4199
rect 94421 3009 94455 3043
rect 94513 4097 94547 4131
rect 99205 4097 99239 4131
rect 99205 3689 99239 3723
rect 99297 3077 99331 3111
rect 94513 3009 94547 3043
rect 134901 9605 134935 9639
rect 111165 6817 111199 6851
rect 109049 3689 109083 3723
rect 109049 2737 109083 2771
rect 100493 561 100527 595
rect 112269 4165 112303 4199
rect 112269 3689 112303 3723
rect 118341 4165 118375 4199
rect 118341 3689 118375 3723
rect 118709 3077 118743 3111
rect 132417 3077 132451 3111
rect 118801 2941 118835 2975
rect 122849 3009 122883 3043
rect 128185 3009 128219 3043
rect 128277 2941 128311 2975
rect 128369 2941 128403 2975
rect 128461 3009 128495 3043
rect 122849 2737 122883 2771
rect 133889 3077 133923 3111
rect 133889 2805 133923 2839
rect 132417 2737 132451 2771
rect 111165 561 111199 595
rect 186053 9605 186087 9639
rect 136741 3009 136775 3043
rect 154037 3009 154071 3043
rect 154129 3009 154163 3043
rect 136741 2805 136775 2839
rect 142813 2941 142847 2975
rect 142813 2805 142847 2839
rect 154129 2805 154163 2839
rect 154221 2805 154255 2839
rect 157257 3077 157291 3111
rect 157257 2805 157291 2839
rect 157349 3077 157383 3111
rect 157349 2805 157383 2839
rect 166917 3077 166951 3111
rect 166917 2805 166951 2839
rect 134901 561 134935 595
rect 258641 9605 258675 9639
rect 208593 3825 208627 3859
rect 208501 3145 208535 3179
rect 208593 3145 208627 3179
rect 209513 3349 209547 3383
rect 201509 2941 201543 2975
rect 209513 3077 209547 3111
rect 219541 3349 219575 3383
rect 249073 3349 249107 3383
rect 248981 3213 249015 3247
rect 219541 3077 219575 3111
rect 220093 3145 220127 3179
rect 208501 2873 208535 2907
rect 211077 3009 211111 3043
rect 201509 2805 201543 2839
rect 220829 3145 220863 3179
rect 220829 3009 220863 3043
rect 229109 3009 229143 3043
rect 220093 2873 220127 2907
rect 229109 2873 229143 2907
rect 234905 3009 234939 3043
rect 248981 3009 249015 3043
rect 249073 2941 249107 2975
rect 234905 2873 234939 2907
rect 211077 2805 211111 2839
rect 186053 561 186087 595
rect 351745 9605 351779 9639
rect 351745 4641 351779 4675
rect 370421 9605 370455 9639
rect 349077 4029 349111 4063
rect 305009 3961 305043 3995
rect 258733 3349 258767 3383
rect 283573 3349 283607 3383
rect 305009 3349 305043 3383
rect 326353 3961 326387 3995
rect 326353 3349 326387 3383
rect 349077 3349 349111 3383
rect 283573 3077 283607 3111
rect 297373 3281 297407 3315
rect 297373 3077 297407 3111
rect 258733 2941 258767 2975
rect 258641 561 258675 595
rect 370421 561 370455 595
rect 371617 9605 371651 9639
rect 371617 561 371651 595
rect 372813 9605 372847 9639
rect 377597 9605 377631 9639
rect 374653 4913 374687 4947
rect 374653 4641 374687 4675
rect 372813 561 372847 595
rect 377597 561 377631 595
rect 378793 9605 378827 9639
rect 428749 9605 428783 9639
rect 393973 3621 394007 3655
rect 393973 3077 394007 3111
rect 415593 3621 415627 3655
rect 415593 3077 415627 3111
rect 378793 561 378827 595
rect 437029 9605 437063 9639
rect 430129 3621 430163 3655
rect 430129 3077 430163 3111
rect 428749 561 428783 595
rect 494989 4301 495023 4335
rect 490665 3349 490699 3383
rect 490573 3213 490607 3247
rect 490573 2805 490607 2839
rect 490665 2805 490699 2839
rect 498853 3825 498887 3859
rect 500233 3621 500267 3655
rect 500233 3349 500267 3383
rect 502993 3213 503027 3247
rect 503269 3213 503303 3247
rect 498853 3145 498887 3179
rect 494989 2805 495023 2839
rect 496737 3077 496771 3111
rect 496737 2805 496771 2839
rect 499497 2805 499531 2839
rect 499589 2737 499623 2771
rect 437029 561 437063 595
<< metal1 >>
rect 335262 700816 335268 700868
rect 335320 700856 335326 700868
rect 429838 700856 429844 700868
rect 335320 700828 429844 700856
rect 335320 700816 335326 700828
rect 429838 700816 429844 700828
rect 429896 700816 429902 700868
rect 283834 700748 283840 700800
rect 283892 700788 283898 700800
rect 343634 700788 343640 700800
rect 283892 700760 343640 700788
rect 283892 700748 283898 700760
rect 343634 700748 343640 700760
rect 343692 700748 343698 700800
rect 364978 700748 364984 700800
rect 365036 700788 365042 700800
rect 508130 700788 508136 700800
rect 365036 700760 508136 700788
rect 365036 700748 365042 700760
rect 508130 700748 508136 700760
rect 508188 700748 508194 700800
rect 78214 700680 78220 700732
rect 78272 700720 78278 700732
rect 235166 700720 235172 700732
rect 78272 700692 235172 700720
rect 78272 700680 78278 700692
rect 235166 700680 235172 700692
rect 235224 700680 235230 700732
rect 269022 700680 269028 700732
rect 269080 700720 269086 700732
rect 300118 700720 300124 700732
rect 269080 700692 300124 700720
rect 269080 700680 269086 700692
rect 300118 700680 300124 700692
rect 300176 700680 300182 700732
rect 332502 700680 332508 700732
rect 332560 700720 332566 700732
rect 501598 700720 501604 700732
rect 332560 700692 501604 700720
rect 332560 700680 332566 700692
rect 501598 700680 501604 700692
rect 501656 700680 501662 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 386414 700652 386420 700664
rect 137888 700624 386420 700652
rect 137888 700612 137894 700624
rect 386414 700612 386420 700624
rect 386472 700612 386478 700664
rect 397454 700612 397460 700664
rect 397512 700652 397518 700664
rect 502518 700652 502524 700664
rect 397512 700624 502524 700652
rect 397512 700612 397518 700624
rect 502518 700612 502524 700624
rect 502576 700612 502582 700664
rect 81894 700544 81900 700596
rect 81952 700584 81958 700596
rect 170306 700584 170312 700596
rect 81952 700556 170312 700584
rect 81952 700544 81958 700556
rect 170306 700544 170312 700556
rect 170364 700544 170370 700596
rect 202782 700544 202788 700596
rect 202840 700584 202846 700596
rect 501782 700584 501788 700596
rect 202840 700556 501788 700584
rect 202840 700544 202846 700556
rect 501782 700544 501788 700556
rect 501840 700544 501846 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 402974 700516 402980 700528
rect 40552 700488 402980 700516
rect 40552 700476 40558 700488
rect 402974 700476 402980 700488
rect 403032 700476 403038 700528
rect 81434 700408 81440 700460
rect 81492 700448 81498 700460
rect 462314 700448 462320 700460
rect 81492 700420 462320 700448
rect 81492 700408 81498 700420
rect 462314 700408 462320 700420
rect 462372 700408 462378 700460
rect 494790 700408 494796 700460
rect 494848 700448 494854 700460
rect 508406 700448 508412 700460
rect 494848 700420 508412 700448
rect 494848 700408 494854 700420
rect 508406 700408 508412 700420
rect 508464 700408 508470 700460
rect 79962 700340 79968 700392
rect 80020 700380 80026 700392
rect 478506 700380 478512 700392
rect 80020 700352 478512 700380
rect 80020 700340 80026 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 504450 700340 504456 700392
rect 504508 700380 504514 700392
rect 543458 700380 543464 700392
rect 504508 700352 543464 700380
rect 504508 700340 504514 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 19978 700312 19984 700324
rect 8168 700284 19984 700312
rect 8168 700272 8174 700284
rect 19978 700272 19984 700284
rect 20036 700272 20042 700324
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 77938 700312 77944 700324
rect 73028 700284 77944 700312
rect 73028 700272 73034 700284
rect 77938 700272 77944 700284
rect 77996 700272 78002 700324
rect 78582 700272 78588 700324
rect 78640 700312 78646 700324
rect 105446 700312 105452 700324
rect 78640 700284 105452 700312
rect 78640 700272 78646 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 142062 700272 142068 700324
rect 142120 700312 142126 700324
rect 559650 700312 559656 700324
rect 142120 700284 559656 700312
rect 142120 700272 142126 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 508774 685856 508780 685908
rect 508832 685896 508838 685908
rect 580166 685896 580172 685908
rect 508832 685868 580172 685896
rect 508832 685856 508838 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 9306 681748 9312 681760
rect 3568 681720 9312 681748
rect 3568 681708 3574 681720
rect 9306 681708 9312 681720
rect 9364 681708 9370 681760
rect 81526 673480 81532 673532
rect 81584 673520 81590 673532
rect 580166 673520 580172 673532
rect 81584 673492 580172 673520
rect 81584 673480 81590 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 502610 667944 502616 667956
rect 3476 667916 502616 667944
rect 3476 667904 3482 667916
rect 502610 667904 502616 667916
rect 502668 667904 502674 667956
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 15930 652780 15936 652792
rect 3108 652752 15936 652780
rect 3108 652740 3114 652752
rect 15930 652740 15936 652752
rect 15988 652740 15994 652792
rect 190362 650020 190368 650072
rect 190420 650060 190426 650072
rect 580166 650060 580172 650072
rect 190420 650032 580172 650060
rect 190420 650020 190426 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 507118 638936 507124 638988
rect 507176 638976 507182 638988
rect 580166 638976 580172 638988
rect 507176 638948 580172 638976
rect 507176 638936 507182 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 82078 626560 82084 626612
rect 82136 626600 82142 626612
rect 580166 626600 580172 626612
rect 82136 626572 580172 626600
rect 82136 626560 82142 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 14458 623812 14464 623824
rect 3476 623784 14464 623812
rect 3476 623772 3482 623784
rect 14458 623772 14464 623784
rect 14516 623772 14522 623824
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 8846 610008 8852 610020
rect 3476 609980 8852 610008
rect 3476 609968 3482 609980
rect 8846 609968 8852 609980
rect 8904 609968 8910 610020
rect 412818 608580 412824 608592
rect 412779 608552 412824 608580
rect 412818 608540 412824 608552
rect 412876 608540 412882 608592
rect 83550 603100 83556 603152
rect 83608 603140 83614 603152
rect 580166 603140 580172 603152
rect 83608 603112 580172 603140
rect 83608 603100 83614 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 412821 601715 412879 601721
rect 412821 601681 412833 601715
rect 412867 601712 412879 601715
rect 413002 601712 413008 601724
rect 412867 601684 413008 601712
rect 412867 601681 412879 601684
rect 412821 601675 412879 601681
rect 413002 601672 413008 601684
rect 413060 601672 413066 601724
rect 412913 598927 412971 598933
rect 412913 598893 412925 598927
rect 412959 598924 412971 598927
rect 413002 598924 413008 598936
rect 412959 598896 413008 598924
rect 412959 598893 412971 598896
rect 412913 598887 412971 598893
rect 413002 598884 413008 598896
rect 413060 598884 413066 598936
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 31110 594844 31116 594856
rect 3292 594816 31116 594844
rect 3292 594804 3298 594816
rect 31110 594804 31116 594816
rect 31168 594804 31174 594856
rect 89346 593308 89352 593360
rect 89404 593348 89410 593360
rect 89438 593348 89444 593360
rect 89404 593320 89444 593348
rect 89404 593308 89410 593320
rect 89438 593308 89444 593320
rect 89496 593308 89502 593360
rect 507210 592016 507216 592068
rect 507268 592056 507274 592068
rect 580166 592056 580172 592068
rect 507268 592028 580172 592056
rect 507268 592016 507274 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 83550 590724 83556 590776
rect 83608 590764 83614 590776
rect 83734 590764 83740 590776
rect 83608 590736 83740 590764
rect 83608 590724 83614 590736
rect 83734 590724 83740 590736
rect 83792 590724 83798 590776
rect 412910 589336 412916 589348
rect 412871 589308 412916 589336
rect 412910 589296 412916 589308
rect 412968 589296 412974 589348
rect 78490 586508 78496 586560
rect 78548 586548 78554 586560
rect 236914 586548 236920 586560
rect 78548 586520 236920 586548
rect 78548 586508 78554 586520
rect 236914 586508 236920 586520
rect 236972 586508 236978 586560
rect 83550 586440 83556 586492
rect 83608 586440 83614 586492
rect 83568 586412 83596 586440
rect 83642 586412 83648 586424
rect 83568 586384 83648 586412
rect 83642 586372 83648 586384
rect 83700 586372 83706 586424
rect 46198 585080 46204 585132
rect 46256 585120 46262 585132
rect 163130 585120 163136 585132
rect 46256 585092 163136 585120
rect 46256 585080 46262 585092
rect 163130 585080 163136 585092
rect 163188 585080 163194 585132
rect 189258 585080 189264 585132
rect 189316 585120 189322 585132
rect 190362 585120 190368 585132
rect 189316 585092 190368 585120
rect 189316 585080 189322 585092
rect 190362 585080 190368 585092
rect 190420 585080 190426 585132
rect 197078 585080 197084 585132
rect 197136 585120 197142 585132
rect 477586 585120 477592 585132
rect 197136 585092 477592 585120
rect 197136 585080 197142 585092
rect 477586 585080 477592 585092
rect 477644 585080 477650 585132
rect 487154 585080 487160 585132
rect 487212 585120 487218 585132
rect 509878 585120 509884 585132
rect 487212 585092 509884 585120
rect 487212 585080 487218 585092
rect 509878 585080 509884 585092
rect 509936 585080 509942 585132
rect 90910 585012 90916 585064
rect 90968 585052 90974 585064
rect 432322 585052 432328 585064
rect 90968 585024 432328 585052
rect 90968 585012 90974 585024
rect 432322 585012 432328 585024
rect 432380 585012 432386 585064
rect 439498 585012 439504 585064
rect 439556 585052 439562 585064
rect 511350 585052 511356 585064
rect 439556 585024 511356 585052
rect 439556 585012 439562 585024
rect 511350 585012 511356 585024
rect 511408 585012 511414 585064
rect 71038 584944 71044 584996
rect 71096 584984 71102 584996
rect 468018 584984 468024 584996
rect 71096 584956 468024 584984
rect 71096 584944 71102 584956
rect 468018 584944 468024 584956
rect 468076 584944 468082 584996
rect 475194 584944 475200 584996
rect 475252 584984 475258 584996
rect 508038 584984 508044 584996
rect 475252 584956 508044 584984
rect 475252 584944 475258 584956
rect 508038 584944 508044 584956
rect 508096 584944 508102 584996
rect 57238 584876 57244 584928
rect 57296 584916 57302 584928
rect 470410 584916 470416 584928
rect 57296 584888 470416 584916
rect 57296 584876 57302 584888
rect 470410 584876 470416 584888
rect 470468 584876 470474 584928
rect 479978 584876 479984 584928
rect 480036 584916 480042 584928
rect 511258 584916 511264 584928
rect 480036 584888 511264 584916
rect 480036 584876 480042 584888
rect 511258 584876 511264 584888
rect 511316 584876 511322 584928
rect 92106 584808 92112 584860
rect 92164 584848 92170 584860
rect 167914 584848 167920 584860
rect 92164 584820 167920 584848
rect 92164 584808 92170 584820
rect 167914 584808 167920 584820
rect 167972 584808 167978 584860
rect 182266 584808 182272 584860
rect 182324 584848 182330 584860
rect 191742 584848 191748 584860
rect 182324 584820 191748 584848
rect 182324 584808 182330 584820
rect 191742 584808 191748 584820
rect 191800 584808 191806 584860
rect 446674 584808 446680 584860
rect 446732 584848 446738 584860
rect 506474 584848 506480 584860
rect 446732 584820 506480 584848
rect 446732 584808 446738 584820
rect 506474 584808 506480 584820
rect 506532 584808 506538 584860
rect 89717 584783 89775 584789
rect 89717 584749 89729 584783
rect 89763 584780 89775 584783
rect 96433 584783 96491 584789
rect 96433 584780 96445 584783
rect 89763 584752 96445 584780
rect 89763 584749 89775 584752
rect 89717 584743 89775 584749
rect 96433 584749 96445 584752
rect 96479 584749 96491 584783
rect 96433 584743 96491 584749
rect 105354 584740 105360 584792
rect 105412 584780 105418 584792
rect 215570 584780 215576 584792
rect 105412 584752 215576 584780
rect 105412 584740 105418 584752
rect 215570 584740 215576 584752
rect 215628 584740 215634 584792
rect 226334 584740 226340 584792
rect 226392 584780 226398 584792
rect 294138 584780 294144 584792
rect 226392 584752 294144 584780
rect 226392 584740 226398 584752
rect 294138 584740 294144 584752
rect 294196 584740 294202 584792
rect 437106 584740 437112 584792
rect 437164 584780 437170 584792
rect 506566 584780 506572 584792
rect 437164 584752 506572 584780
rect 437164 584740 437170 584752
rect 506566 584740 506572 584752
rect 506624 584740 506630 584792
rect 77018 584672 77024 584724
rect 77076 584712 77082 584724
rect 103514 584712 103520 584724
rect 77076 584684 103520 584712
rect 77076 584672 77082 584684
rect 103514 584672 103520 584684
rect 103572 584672 103578 584724
rect 117866 584672 117872 584724
rect 117924 584712 117930 584724
rect 233234 584712 233240 584724
rect 117924 584684 233240 584712
rect 117924 584672 117930 584684
rect 233234 584672 233240 584684
rect 233292 584672 233298 584724
rect 238754 584672 238760 584724
rect 238812 584712 238818 584724
rect 244090 584712 244096 584724
rect 238812 584684 244096 584712
rect 238812 584672 238818 584684
rect 244090 584672 244096 584684
rect 244148 584672 244154 584724
rect 456058 584672 456064 584724
rect 456116 584712 456122 584724
rect 507946 584712 507952 584724
rect 456116 584684 507952 584712
rect 456116 584672 456122 584684
rect 507946 584672 507952 584684
rect 508004 584672 508010 584724
rect 61378 584604 61384 584656
rect 61436 584644 61442 584656
rect 217962 584644 217968 584656
rect 61436 584616 217968 584644
rect 61436 584604 61442 584616
rect 217962 584604 217968 584616
rect 218020 584604 218026 584656
rect 227806 584604 227812 584656
rect 227864 584644 227870 584656
rect 234522 584644 234528 584656
rect 227864 584616 234528 584644
rect 227864 584604 227870 584616
rect 234522 584604 234528 584616
rect 234580 584604 234586 584656
rect 249702 584604 249708 584656
rect 249760 584644 249766 584656
rect 372706 584644 372712 584656
rect 249760 584616 372712 584644
rect 249760 584604 249766 584616
rect 372706 584604 372712 584616
rect 372764 584604 372770 584656
rect 377490 584604 377496 584656
rect 377548 584644 377554 584656
rect 494698 584644 494704 584656
rect 377548 584616 494704 584644
rect 377548 584604 377554 584616
rect 494698 584604 494704 584616
rect 494756 584604 494762 584656
rect 498105 584647 498163 584653
rect 498105 584613 498117 584647
rect 498151 584644 498163 584647
rect 508314 584644 508320 584656
rect 498151 584616 508320 584644
rect 498151 584613 498163 584616
rect 498105 584607 498163 584613
rect 508314 584604 508320 584616
rect 508372 584604 508378 584656
rect 59998 584536 60004 584588
rect 60056 584576 60062 584588
rect 248874 584576 248880 584588
rect 60056 584548 248880 584576
rect 60056 584536 60062 584548
rect 248874 584536 248880 584548
rect 248932 584536 248938 584588
rect 348970 584536 348976 584588
rect 349028 584576 349034 584588
rect 485774 584576 485780 584588
rect 349028 584548 485780 584576
rect 349028 584536 349034 584548
rect 485774 584536 485780 584548
rect 485832 584536 485838 584588
rect 491938 584536 491944 584588
rect 491996 584576 492002 584588
rect 511166 584576 511172 584588
rect 491996 584548 511172 584576
rect 491996 584536 492002 584548
rect 511166 584536 511172 584548
rect 511224 584536 511230 584588
rect 64138 584468 64144 584520
rect 64196 584508 64202 584520
rect 270402 584508 270408 584520
rect 64196 584480 270408 584508
rect 64196 584468 64202 584480
rect 270402 584468 270408 584480
rect 270460 584468 270466 584520
rect 382274 584468 382280 584520
rect 382332 584508 382338 584520
rect 524414 584508 524420 584520
rect 382332 584480 524420 584508
rect 382332 584468 382338 584480
rect 524414 584468 524420 584480
rect 524472 584468 524478 584520
rect 50338 584400 50344 584452
rect 50396 584440 50402 584452
rect 272794 584440 272800 584452
rect 50396 584412 272800 584440
rect 50396 584400 50402 584412
rect 272794 584400 272800 584412
rect 272852 584400 272858 584452
rect 444282 584400 444288 584452
rect 444340 584440 444346 584452
rect 498105 584443 498163 584449
rect 498105 584440 498117 584443
rect 444340 584412 498117 584440
rect 444340 584400 444346 584412
rect 498105 584409 498117 584412
rect 498151 584409 498163 584443
rect 498105 584403 498163 584409
rect 500221 584443 500279 584449
rect 500221 584409 500233 584443
rect 500267 584440 500279 584443
rect 505278 584440 505284 584452
rect 500267 584412 505284 584440
rect 500267 584409 500279 584412
rect 500221 584403 500279 584409
rect 505278 584400 505284 584412
rect 505336 584400 505342 584452
rect 53098 584332 53104 584384
rect 53156 584372 53162 584384
rect 322658 584372 322664 584384
rect 53156 584344 322664 584372
rect 53156 584332 53162 584344
rect 322658 584332 322664 584344
rect 322716 584332 322722 584384
rect 367922 584332 367928 584384
rect 367980 584372 367986 584384
rect 510798 584372 510804 584384
rect 367980 584344 510804 584372
rect 367980 584332 367986 584344
rect 510798 584332 510804 584344
rect 510856 584332 510862 584384
rect 31018 584264 31024 584316
rect 31076 584304 31082 584316
rect 310882 584304 310888 584316
rect 31076 584276 310888 584304
rect 31076 584264 31082 584276
rect 310882 584264 310888 584276
rect 310940 584264 310946 584316
rect 341794 584264 341800 584316
rect 341852 584304 341858 584316
rect 501506 584304 501512 584316
rect 341852 584276 501512 584304
rect 341852 584264 341858 584276
rect 501506 584264 501512 584276
rect 501564 584264 501570 584316
rect 76926 584196 76932 584248
rect 76984 584236 76990 584248
rect 210786 584236 210792 584248
rect 76984 584208 210792 584236
rect 76984 584196 76990 584208
rect 210786 584196 210792 584208
rect 210844 584196 210850 584248
rect 339402 584196 339408 584248
rect 339460 584236 339466 584248
rect 456794 584236 456800 584248
rect 339460 584208 456800 584236
rect 339460 584196 339466 584208
rect 456794 584196 456800 584208
rect 456852 584196 456858 584248
rect 458450 584196 458456 584248
rect 458508 584236 458514 584248
rect 500221 584239 500279 584245
rect 500221 584236 500233 584239
rect 458508 584208 500233 584236
rect 458508 584196 458514 584208
rect 500221 584205 500233 584208
rect 500267 584205 500279 584239
rect 500221 584199 500279 584205
rect 500313 584239 500371 584245
rect 500313 584205 500325 584239
rect 500359 584236 500371 584239
rect 505370 584236 505376 584248
rect 500359 584208 505376 584236
rect 500359 584205 500371 584208
rect 500313 584199 500371 584205
rect 505370 584196 505376 584208
rect 505428 584196 505434 584248
rect 51718 584128 51724 584180
rect 51776 584168 51782 584180
rect 356146 584168 356152 584180
rect 51776 584140 356152 584168
rect 51776 584128 51782 584140
rect 356146 584128 356152 584140
rect 356204 584128 356210 584180
rect 370314 584128 370320 584180
rect 370372 584168 370378 584180
rect 556154 584168 556160 584180
rect 370372 584140 556160 584168
rect 370372 584128 370378 584140
rect 556154 584128 556160 584140
rect 556212 584128 556218 584180
rect 75178 584060 75184 584112
rect 75236 584100 75242 584112
rect 89717 584103 89775 584109
rect 89717 584100 89729 584103
rect 75236 584072 89729 584100
rect 75236 584060 75242 584072
rect 89717 584069 89729 584072
rect 89763 584069 89775 584103
rect 106461 584103 106519 584109
rect 106461 584100 106473 584103
rect 89717 584063 89775 584069
rect 106200 584072 106473 584100
rect 77202 583992 77208 584044
rect 77260 584032 77266 584044
rect 96338 584032 96344 584044
rect 77260 584004 96344 584032
rect 77260 583992 77266 584004
rect 96338 583992 96344 584004
rect 96396 583992 96402 584044
rect 96433 584035 96491 584041
rect 96433 584001 96445 584035
rect 96479 584032 96491 584035
rect 106200 584032 106228 584072
rect 106461 584069 106473 584072
rect 106507 584069 106519 584103
rect 106461 584063 106519 584069
rect 124125 584103 124183 584109
rect 124125 584069 124137 584103
rect 124171 584100 124183 584103
rect 124171 584072 128400 584100
rect 124171 584069 124183 584072
rect 124125 584063 124183 584069
rect 96479 584004 106228 584032
rect 128372 584032 128400 584072
rect 131942 584060 131948 584112
rect 132000 584100 132006 584112
rect 449066 584100 449072 584112
rect 132000 584072 449072 584100
rect 132000 584060 132006 584072
rect 449066 584060 449072 584072
rect 449124 584060 449130 584112
rect 453850 584060 453856 584112
rect 453908 584100 453914 584112
rect 534074 584100 534080 584112
rect 453908 584072 534080 584100
rect 453908 584060 453914 584072
rect 534074 584060 534080 584072
rect 534132 584060 534138 584112
rect 136818 584032 136824 584044
rect 128372 584004 136824 584032
rect 96479 584001 96491 584004
rect 96433 583995 96491 584001
rect 136818 583992 136824 584004
rect 136876 583992 136882 584044
rect 141602 583992 141608 584044
rect 141660 584032 141666 584044
rect 142062 584032 142068 584044
rect 141660 584004 142068 584032
rect 141660 583992 141666 584004
rect 142062 583992 142068 584004
rect 142120 583992 142126 584044
rect 170306 583992 170312 584044
rect 170364 584032 170370 584044
rect 490374 584032 490380 584044
rect 170364 584004 490380 584032
rect 170364 583992 170370 584004
rect 490374 583992 490380 584004
rect 490432 583992 490438 584044
rect 494330 583992 494336 584044
rect 494388 584032 494394 584044
rect 511534 584032 511540 584044
rect 494388 584004 511540 584032
rect 494388 583992 494394 584004
rect 511534 583992 511540 584004
rect 511592 583992 511598 584044
rect 73798 583924 73804 583976
rect 73856 583964 73862 583976
rect 127434 583964 127440 583976
rect 73856 583936 127440 583964
rect 73856 583924 73862 583936
rect 127434 583924 127440 583936
rect 127492 583924 127498 583976
rect 268010 583924 268016 583976
rect 268068 583964 268074 583976
rect 269022 583964 269028 583976
rect 268068 583936 269028 583964
rect 268068 583924 268074 583936
rect 269022 583924 269028 583936
rect 269080 583924 269086 583976
rect 289354 583924 289360 583976
rect 289412 583964 289418 583976
rect 455322 583964 455328 583976
rect 289412 583936 455328 583964
rect 289412 583924 289418 583936
rect 455322 583924 455328 583936
rect 455380 583924 455386 583976
rect 484762 583924 484768 583976
rect 484820 583964 484826 583976
rect 509786 583964 509792 583976
rect 484820 583936 509792 583964
rect 484820 583924 484826 583936
rect 509786 583924 509792 583936
rect 509844 583924 509850 583976
rect 42058 583856 42064 583908
rect 42116 583896 42122 583908
rect 413186 583896 413192 583908
rect 42116 583868 413192 583896
rect 42116 583856 42122 583868
rect 413186 583856 413192 583868
rect 413244 583856 413250 583908
rect 422754 583856 422760 583908
rect 422812 583896 422818 583908
rect 509418 583896 509424 583908
rect 422812 583868 509424 583896
rect 422812 583856 422818 583868
rect 509418 583856 509424 583868
rect 509476 583856 509482 583908
rect 78306 583788 78312 583840
rect 78364 583828 78370 583840
rect 105906 583828 105912 583840
rect 78364 583800 105912 583828
rect 78364 583788 78370 583800
rect 105906 583788 105912 583800
rect 105964 583788 105970 583840
rect 107654 583788 107660 583840
rect 107712 583828 107718 583840
rect 125042 583828 125048 583840
rect 107712 583800 125048 583828
rect 107712 583788 107718 583800
rect 125042 583788 125048 583800
rect 125100 583788 125106 583840
rect 415578 583788 415584 583840
rect 415636 583828 415642 583840
rect 502334 583828 502340 583840
rect 415636 583800 502340 583828
rect 415636 583788 415642 583800
rect 502334 583788 502340 583800
rect 502392 583788 502398 583840
rect 78398 583720 78404 583772
rect 78456 583760 78462 583772
rect 113082 583760 113088 583772
rect 78456 583732 113088 583760
rect 78456 583720 78462 583732
rect 113082 583720 113088 583732
rect 113140 583720 113146 583772
rect 308490 583720 308496 583772
rect 308548 583760 308554 583772
rect 314654 583760 314660 583772
rect 308548 583732 314660 583760
rect 308548 583720 308554 583732
rect 314654 583720 314660 583732
rect 314712 583720 314718 583772
rect 408586 583720 408592 583772
rect 408644 583760 408650 583772
rect 424962 583760 424968 583772
rect 408644 583732 424968 583760
rect 408644 583720 408650 583732
rect 424962 583720 424968 583732
rect 425020 583720 425026 583772
rect 429930 583720 429936 583772
rect 429988 583760 429994 583772
rect 500313 583763 500371 583769
rect 500313 583760 500325 583763
rect 429988 583732 500325 583760
rect 429988 583720 429994 583732
rect 500313 583729 500325 583732
rect 500359 583729 500371 583763
rect 500313 583723 500371 583729
rect 501322 583720 501328 583772
rect 501380 583760 501386 583772
rect 505830 583760 505836 583772
rect 501380 583732 505836 583760
rect 501380 583720 501386 583732
rect 505830 583720 505836 583732
rect 505888 583720 505894 583772
rect 106461 583695 106519 583701
rect 106461 583661 106473 583695
rect 106507 583692 106519 583695
rect 124125 583695 124183 583701
rect 124125 583692 124137 583695
rect 106507 583664 124137 583692
rect 106507 583661 106519 583664
rect 106461 583655 106519 583661
rect 124125 583661 124137 583664
rect 124171 583661 124183 583695
rect 124125 583655 124183 583661
rect 35802 583448 35808 583500
rect 35860 583488 35866 583500
rect 441890 583488 441896 583500
rect 35860 583460 441896 583488
rect 35860 583448 35866 583460
rect 441890 583448 441896 583460
rect 441948 583448 441954 583500
rect 485774 583448 485780 583500
rect 485832 583488 485838 583500
rect 502978 583488 502984 583500
rect 485832 583460 502984 583488
rect 485832 583448 485838 583460
rect 502978 583448 502984 583460
rect 503036 583448 503042 583500
rect 75822 583380 75828 583432
rect 75880 583420 75886 583432
rect 131942 583420 131948 583432
rect 75880 583392 131948 583420
rect 75880 583380 75886 583392
rect 131942 583380 131948 583392
rect 132000 583380 132006 583432
rect 456794 583380 456800 583432
rect 456852 583420 456858 583432
rect 509510 583420 509516 583432
rect 456852 583392 509516 583420
rect 456852 583380 456858 583392
rect 509510 583380 509516 583392
rect 509568 583380 509574 583432
rect 77110 583312 77116 583364
rect 77168 583352 77174 583364
rect 197078 583352 197084 583364
rect 77168 583324 197084 583352
rect 77168 583312 77174 583324
rect 197078 583312 197084 583324
rect 197136 583312 197142 583364
rect 455322 583312 455328 583364
rect 455380 583352 455386 583364
rect 510982 583352 510988 583364
rect 455380 583324 510988 583352
rect 455380 583312 455386 583324
rect 510982 583312 510988 583324
rect 511040 583312 511046 583364
rect 75270 583244 75276 583296
rect 75328 583284 75334 583296
rect 279786 583284 279792 583296
rect 75328 583256 279792 583284
rect 75328 583244 75334 583256
rect 279786 583244 279792 583256
rect 279844 583244 279850 583296
rect 410794 583244 410800 583296
rect 410852 583284 410858 583296
rect 503346 583284 503352 583296
rect 410852 583256 503352 583284
rect 410852 583244 410858 583256
rect 503346 583244 503352 583256
rect 503404 583244 503410 583296
rect 10410 583176 10416 583228
rect 10468 583216 10474 583228
rect 256050 583216 256056 583228
rect 10468 583188 256056 583216
rect 10468 583176 10474 583188
rect 256050 583176 256056 583188
rect 256108 583176 256114 583228
rect 379882 583176 379888 583228
rect 379940 583216 379946 583228
rect 503070 583216 503076 583228
rect 379940 583188 503076 583216
rect 379940 583176 379946 583188
rect 503070 583176 503076 583188
rect 503128 583176 503134 583228
rect 9490 583108 9496 583160
rect 9548 583148 9554 583160
rect 265618 583148 265624 583160
rect 9548 583120 265624 583148
rect 9548 583108 9554 583120
rect 265618 583108 265624 583120
rect 265676 583108 265682 583160
rect 337010 583108 337016 583160
rect 337068 583148 337074 583160
rect 509694 583148 509700 583160
rect 337068 583120 509700 583148
rect 337068 583108 337074 583120
rect 509694 583108 509700 583120
rect 509752 583108 509758 583160
rect 10594 583040 10600 583092
rect 10652 583080 10658 583092
rect 284570 583080 284576 583092
rect 10652 583052 284576 583080
rect 10652 583040 10658 583052
rect 284570 583040 284576 583052
rect 284628 583040 284634 583092
rect 327442 583040 327448 583092
rect 327500 583080 327506 583092
rect 507670 583080 507676 583092
rect 327500 583052 507676 583080
rect 327500 583040 327506 583052
rect 507670 583040 507676 583052
rect 507728 583040 507734 583092
rect 77754 582972 77760 583024
rect 77812 583012 77818 583024
rect 353754 583012 353760 583024
rect 77812 582984 353760 583012
rect 77812 582972 77818 582984
rect 353754 582972 353760 582984
rect 353812 582972 353818 583024
rect 360930 582972 360936 583024
rect 360988 583012 360994 583024
rect 510062 583012 510068 583024
rect 360988 582984 510068 583012
rect 360988 582972 360994 582984
rect 510062 582972 510068 582984
rect 510120 582972 510126 583024
rect 80698 582904 80704 582956
rect 80756 582944 80762 582956
rect 198826 582944 198832 582956
rect 80756 582916 198832 582944
rect 80756 582904 80762 582916
rect 198826 582904 198832 582916
rect 198884 582904 198890 582956
rect 229738 582904 229744 582956
rect 229796 582944 229802 582956
rect 510890 582944 510896 582956
rect 229796 582916 510896 582944
rect 229796 582904 229802 582916
rect 510890 582904 510896 582916
rect 510948 582904 510954 582956
rect 184474 582836 184480 582888
rect 184532 582876 184538 582888
rect 503254 582876 503260 582888
rect 184532 582848 503260 582876
rect 184532 582836 184538 582848
rect 503254 582836 503260 582848
rect 503312 582836 503318 582888
rect 15838 582768 15844 582820
rect 15896 582808 15902 582820
rect 110690 582808 110696 582820
rect 15896 582780 110696 582808
rect 15896 582768 15902 582780
rect 110690 582768 110696 582780
rect 110748 582768 110754 582820
rect 177482 582768 177488 582820
rect 177540 582808 177546 582820
rect 501966 582808 501972 582820
rect 177540 582780 501972 582808
rect 177540 582768 177546 582780
rect 501966 582768 501972 582780
rect 502024 582768 502030 582820
rect 8938 582700 8944 582752
rect 8996 582740 9002 582752
rect 146386 582740 146392 582752
rect 8996 582712 146392 582740
rect 8996 582700 9002 582712
rect 146386 582700 146392 582712
rect 146444 582700 146450 582752
rect 220354 582700 220360 582752
rect 220412 582740 220418 582752
rect 560938 582740 560944 582752
rect 220412 582712 560944 582740
rect 220412 582700 220418 582712
rect 560938 582700 560944 582712
rect 560996 582700 561002 582752
rect 10686 582632 10692 582684
rect 10744 582672 10750 582684
rect 129826 582672 129832 582684
rect 10744 582644 129832 582672
rect 10744 582632 10750 582644
rect 129826 582632 129832 582644
rect 129884 582632 129890 582684
rect 132218 582632 132224 582684
rect 132276 582672 132282 582684
rect 503162 582672 503168 582684
rect 132276 582644 503168 582672
rect 132276 582632 132282 582644
rect 503162 582632 503168 582644
rect 503220 582632 503226 582684
rect 86310 582564 86316 582616
rect 86368 582604 86374 582616
rect 96522 582604 96528 582616
rect 86368 582576 96528 582604
rect 86368 582564 86374 582576
rect 96522 582564 96528 582576
rect 96580 582564 96586 582616
rect 96614 582564 96620 582616
rect 96672 582604 96678 582616
rect 99929 582607 99987 582613
rect 99929 582604 99941 582607
rect 96672 582576 99941 582604
rect 96672 582564 96678 582576
rect 99929 582573 99941 582576
rect 99975 582573 99987 582607
rect 99929 582567 99987 582573
rect 101306 582564 101312 582616
rect 101364 582604 101370 582616
rect 115842 582604 115848 582616
rect 101364 582576 115848 582604
rect 101364 582564 101370 582576
rect 115842 582564 115848 582576
rect 115900 582564 115906 582616
rect 425146 582564 425152 582616
rect 425204 582604 425210 582616
rect 514018 582604 514024 582616
rect 425204 582576 514024 582604
rect 425204 582564 425210 582576
rect 514018 582564 514024 582576
rect 514076 582564 514082 582616
rect 64782 582496 64788 582548
rect 64840 582536 64846 582548
rect 499114 582536 499120 582548
rect 64840 582508 499120 582536
rect 64840 582496 64846 582508
rect 499114 582496 499120 582508
rect 499172 582496 499178 582548
rect 9582 582428 9588 582480
rect 9640 582468 9646 582480
rect 463234 582468 463240 582480
rect 9640 582440 463240 582468
rect 9640 582428 9646 582440
rect 463234 582428 463240 582440
rect 463292 582428 463298 582480
rect 482370 582428 482376 582480
rect 482428 582468 482434 582480
rect 507486 582468 507492 582480
rect 482428 582440 507492 582468
rect 482428 582428 482434 582440
rect 507486 582428 507492 582440
rect 507544 582428 507550 582480
rect 6178 582360 6184 582412
rect 6236 582400 6242 582412
rect 489546 582400 489552 582412
rect 6236 582372 489552 582400
rect 6236 582360 6242 582372
rect 489546 582360 489552 582372
rect 489604 582360 489610 582412
rect 490190 582360 490196 582412
rect 490248 582400 490254 582412
rect 497550 582400 497556 582412
rect 490248 582372 497556 582400
rect 490248 582360 490254 582372
rect 497550 582360 497556 582372
rect 497608 582360 497614 582412
rect 90450 582292 90456 582344
rect 90508 582332 90514 582344
rect 99834 582332 99840 582344
rect 90508 582304 99840 582332
rect 90508 582292 90514 582304
rect 99834 582292 99840 582304
rect 99892 582292 99898 582344
rect 99929 582335 99987 582341
rect 99929 582301 99941 582335
rect 99975 582332 99987 582335
rect 111058 582332 111064 582344
rect 99975 582304 111064 582332
rect 99975 582301 99987 582304
rect 99929 582295 99987 582301
rect 111058 582292 111064 582304
rect 111116 582292 111122 582344
rect 460842 582292 460848 582344
rect 460900 582332 460906 582344
rect 510706 582332 510712 582344
rect 460900 582304 510712 582332
rect 460900 582292 460906 582304
rect 510706 582292 510712 582304
rect 510764 582292 510770 582344
rect 10502 582224 10508 582276
rect 10560 582264 10566 582276
rect 93946 582264 93952 582276
rect 10560 582236 93952 582264
rect 10560 582224 10566 582236
rect 93946 582224 93952 582236
rect 94004 582224 94010 582276
rect 100018 582224 100024 582276
rect 100076 582264 100082 582276
rect 105354 582264 105360 582276
rect 100076 582236 105360 582264
rect 100076 582224 100082 582236
rect 105354 582224 105360 582236
rect 105412 582224 105418 582276
rect 118694 582224 118700 582276
rect 118752 582264 118758 582276
rect 123754 582264 123760 582276
rect 118752 582236 123760 582264
rect 118752 582224 118758 582236
rect 123754 582224 123760 582236
rect 123812 582224 123818 582276
rect 150986 582224 150992 582276
rect 151044 582264 151050 582276
rect 157150 582264 157156 582276
rect 151044 582236 157156 582264
rect 151044 582224 151050 582236
rect 157150 582224 157156 582236
rect 157208 582224 157214 582276
rect 157242 582224 157248 582276
rect 157300 582264 157306 582276
rect 162486 582264 162492 582276
rect 157300 582236 162492 582264
rect 157300 582224 157306 582236
rect 162486 582224 162492 582236
rect 162544 582224 162550 582276
rect 494698 582224 494704 582276
rect 494756 582264 494762 582276
rect 511074 582264 511080 582276
rect 494756 582236 511080 582264
rect 494756 582224 494762 582236
rect 511074 582224 511080 582236
rect 511132 582224 511138 582276
rect 93210 582156 93216 582208
rect 93268 582196 93274 582208
rect 122650 582196 122656 582208
rect 93268 582168 122656 582196
rect 93268 582156 93274 582168
rect 122650 582156 122656 582168
rect 122708 582156 122714 582208
rect 128354 582156 128360 582208
rect 128412 582196 128418 582208
rect 137922 582196 137928 582208
rect 128412 582168 137928 582196
rect 128412 582156 128418 582168
rect 137922 582156 137928 582168
rect 137980 582156 137986 582208
rect 146938 582156 146944 582208
rect 146996 582196 147002 582208
rect 160462 582196 160468 582208
rect 146996 582168 160468 582196
rect 146996 582156 147002 582168
rect 160462 582156 160468 582168
rect 160520 582156 160526 582208
rect 167086 582156 167092 582208
rect 167144 582196 167150 582208
rect 176562 582196 176568 582208
rect 167144 582168 176568 582196
rect 167144 582156 167150 582168
rect 176562 582156 176568 582168
rect 176620 582156 176626 582208
rect 401410 582156 401416 582208
rect 401468 582196 401474 582208
rect 502058 582196 502064 582208
rect 401468 582168 502064 582196
rect 401468 582156 401474 582168
rect 502058 582156 502064 582168
rect 502116 582156 502122 582208
rect 73062 582088 73068 582140
rect 73120 582128 73126 582140
rect 226334 582128 226340 582140
rect 73120 582100 226340 582128
rect 73120 582088 73126 582100
rect 226334 582088 226340 582100
rect 226392 582088 226398 582140
rect 406194 582088 406200 582140
rect 406252 582128 406258 582140
rect 509326 582128 509332 582140
rect 406252 582100 509332 582128
rect 406252 582088 406258 582100
rect 509326 582088 509332 582100
rect 509384 582088 509390 582140
rect 89714 582020 89720 582072
rect 89772 582060 89778 582072
rect 91922 582060 91928 582072
rect 89772 582032 91928 582060
rect 89772 582020 89778 582032
rect 91922 582020 91928 582032
rect 91980 582020 91986 582072
rect 92658 582020 92664 582072
rect 92716 582060 92722 582072
rect 286686 582060 286692 582072
rect 92716 582032 286692 582060
rect 92716 582020 92722 582032
rect 286686 582020 286692 582032
rect 286744 582020 286750 582072
rect 394602 582020 394608 582072
rect 394660 582060 394666 582072
rect 509602 582060 509608 582072
rect 394660 582032 509608 582060
rect 394660 582020 394666 582032
rect 509602 582020 509608 582032
rect 509660 582020 509666 582072
rect 85206 581952 85212 582004
rect 85264 581992 85270 582004
rect 320174 581992 320180 582004
rect 85264 581964 320180 581992
rect 85264 581952 85270 581964
rect 320174 581952 320180 581964
rect 320232 581952 320238 582004
rect 321554 581952 321560 582004
rect 321612 581992 321618 582004
rect 326430 581992 326436 582004
rect 321612 581964 326436 581992
rect 321612 581952 321618 581964
rect 326430 581952 326436 581964
rect 326488 581952 326494 582004
rect 363690 581952 363696 582004
rect 363748 581992 363754 582004
rect 501874 581992 501880 582004
rect 363748 581964 501880 581992
rect 363748 581952 363754 581964
rect 501874 581952 501880 581964
rect 501932 581952 501938 582004
rect 48222 581884 48228 581936
rect 48280 581924 48286 581936
rect 372614 581924 372620 581936
rect 48280 581896 372620 581924
rect 48280 581884 48286 581896
rect 372614 581884 372620 581896
rect 372672 581884 372678 581936
rect 399386 581884 399392 581936
rect 399444 581924 399450 581936
rect 543734 581924 543740 581936
rect 399444 581896 543740 581924
rect 399444 581884 399450 581896
rect 543734 581884 543740 581896
rect 543792 581884 543798 581936
rect 3418 581816 3424 581868
rect 3476 581856 3482 581868
rect 262950 581856 262956 581868
rect 3476 581828 262956 581856
rect 3476 581816 3482 581828
rect 262950 581816 262956 581828
rect 263008 581816 263014 581868
rect 296714 581816 296720 581868
rect 296772 581856 296778 581868
rect 510614 581856 510620 581868
rect 296772 581828 510620 581856
rect 296772 581816 296778 581828
rect 510614 581816 510620 581828
rect 510672 581816 510678 581868
rect 85482 581748 85488 581800
rect 85540 581788 85546 581800
rect 172514 581788 172520 581800
rect 85540 581760 172520 581788
rect 85540 581748 85546 581760
rect 172514 581748 172520 581760
rect 172572 581748 172578 581800
rect 186314 581748 186320 581800
rect 186372 581788 186378 581800
rect 192202 581788 192208 581800
rect 186372 581760 192208 581788
rect 186372 581748 186378 581760
rect 192202 581748 192208 581760
rect 192260 581748 192266 581800
rect 246850 581748 246856 581800
rect 246908 581788 246914 581800
rect 508222 581788 508228 581800
rect 246908 581760 508228 581788
rect 246908 581748 246914 581760
rect 508222 581748 508228 581760
rect 508280 581748 508286 581800
rect 52362 581680 52368 581732
rect 52420 581720 52426 581732
rect 249702 581720 249708 581732
rect 52420 581692 249708 581720
rect 52420 581680 52426 581692
rect 249702 581680 249708 581692
rect 249760 581680 249766 581732
rect 251634 581680 251640 581732
rect 251692 581720 251698 581732
rect 554866 581720 554872 581732
rect 251692 581692 554872 581720
rect 251692 581680 251698 581692
rect 554866 581680 554872 581692
rect 554924 581680 554930 581732
rect 9122 581612 9128 581664
rect 9180 581652 9186 581664
rect 120074 581652 120080 581664
rect 9180 581624 120080 581652
rect 9180 581612 9186 581624
rect 120074 581612 120080 581624
rect 120132 581612 120138 581664
rect 134334 581652 134340 581664
rect 134295 581624 134340 581652
rect 134334 581612 134340 581624
rect 134392 581612 134398 581664
rect 144362 581652 144368 581664
rect 144323 581624 144368 581652
rect 144362 581612 144368 581624
rect 144420 581612 144426 581664
rect 157058 581612 157064 581664
rect 157116 581652 157122 581664
rect 157518 581652 157524 581664
rect 157116 581624 157524 581652
rect 157116 581612 157122 581624
rect 157518 581612 157524 581624
rect 157576 581612 157582 581664
rect 197998 581612 198004 581664
rect 198056 581652 198062 581664
rect 200850 581652 200856 581664
rect 198056 581624 200856 581652
rect 198056 581612 198062 581624
rect 200850 581612 200856 581624
rect 200908 581612 200914 581664
rect 227714 581612 227720 581664
rect 227772 581652 227778 581664
rect 532694 581652 532700 581664
rect 227772 581624 532700 581652
rect 227772 581612 227778 581624
rect 532694 581612 532700 581624
rect 532752 581612 532758 581664
rect 4798 581544 4804 581596
rect 4856 581584 4862 581596
rect 313182 581584 313188 581596
rect 4856 581556 313188 581584
rect 4856 581544 4862 581556
rect 313182 581544 313188 581556
rect 313240 581544 313246 581596
rect 375282 581544 375288 581596
rect 375340 581584 375346 581596
rect 569954 581584 569960 581596
rect 375340 581556 569960 581584
rect 375340 581544 375346 581556
rect 569954 581544 569960 581556
rect 570012 581544 570018 581596
rect 10318 581476 10324 581528
rect 10376 581516 10382 581528
rect 165246 581516 165252 581528
rect 10376 581488 165252 581516
rect 10376 581476 10382 581488
rect 165246 581476 165252 581488
rect 165304 581476 165310 581528
rect 176562 581476 176568 581528
rect 176620 581516 176626 581528
rect 176746 581516 176752 581528
rect 176620 581488 176752 581516
rect 176620 581476 176626 581488
rect 176746 581476 176752 581488
rect 176804 581476 176810 581528
rect 194410 581476 194416 581528
rect 194468 581516 194474 581528
rect 505094 581516 505100 581528
rect 194468 581488 505100 581516
rect 194468 581476 194474 581488
rect 505094 581476 505100 581488
rect 505152 581476 505158 581528
rect 67542 581408 67548 581460
rect 67600 581448 67606 581460
rect 420086 581448 420092 581460
rect 67600 581420 420092 581448
rect 67600 581408 67606 581420
rect 420086 581408 420092 581420
rect 420144 581408 420150 581460
rect 435082 581408 435088 581460
rect 435140 581448 435146 581460
rect 580534 581448 580540 581460
rect 435140 581420 580540 581448
rect 435140 581408 435146 581420
rect 580534 581408 580540 581420
rect 580592 581408 580598 581460
rect 9214 581340 9220 581392
rect 9272 581380 9278 581392
rect 98454 581380 98460 581392
rect 9272 581352 98460 581380
rect 9272 581340 9278 581352
rect 98454 581340 98460 581352
rect 98512 581340 98518 581392
rect 99466 581340 99472 581392
rect 99524 581380 99530 581392
rect 103422 581380 103428 581392
rect 99524 581352 103428 581380
rect 99524 581340 99530 581352
rect 103422 581340 103428 581352
rect 103480 581340 103486 581392
rect 108666 581340 108672 581392
rect 108724 581380 108730 581392
rect 491846 581380 491852 581392
rect 108724 581352 491852 581380
rect 108724 581340 108730 581352
rect 491846 581340 491852 581352
rect 491904 581340 491910 581392
rect 494606 581340 494612 581392
rect 494664 581380 494670 581392
rect 504358 581380 504364 581392
rect 494664 581352 504364 581380
rect 494664 581340 494670 581352
rect 504358 581340 504364 581352
rect 504416 581340 504422 581392
rect 82630 581272 82636 581324
rect 82688 581312 82694 581324
rect 580350 581312 580356 581324
rect 82688 581284 580356 581312
rect 82688 581272 82694 581284
rect 580350 581272 580356 581284
rect 580408 581272 580414 581324
rect 9030 581204 9036 581256
rect 9088 581244 9094 581256
rect 134337 581247 134395 581253
rect 134337 581244 134349 581247
rect 9088 581216 134349 581244
rect 9088 581204 9094 581216
rect 134337 581213 134349 581216
rect 134383 581213 134395 581247
rect 134337 581207 134395 581213
rect 144365 581247 144423 581253
rect 144365 581213 144377 581247
rect 144411 581244 144423 581247
rect 580442 581244 580448 581256
rect 144411 581216 580448 581244
rect 144411 581213 144423 581216
rect 144365 581207 144423 581213
rect 580442 581204 580448 581216
rect 580500 581204 580506 581256
rect 501690 581068 501696 581120
rect 501748 581108 501754 581120
rect 501874 581108 501880 581120
rect 501748 581080 501880 581108
rect 501748 581068 501754 581080
rect 501874 581068 501880 581080
rect 501932 581068 501938 581120
rect 502058 581040 502064 581052
rect 501892 581012 502064 581040
rect 501892 580984 501920 581012
rect 502058 581000 502064 581012
rect 502116 581000 502122 581052
rect 501874 580932 501880 580984
rect 501932 580932 501938 580984
rect 507302 579640 507308 579692
rect 507360 579680 507366 579692
rect 580166 579680 580172 579692
rect 507360 579652 580172 579680
rect 507360 579640 507366 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 48958 572704 48964 572756
rect 49016 572744 49022 572756
rect 78674 572744 78680 572756
rect 49016 572716 78680 572744
rect 49016 572704 49022 572716
rect 78674 572704 78680 572716
rect 78732 572704 78738 572756
rect 532694 568556 532700 568608
rect 532752 568596 532758 568608
rect 532878 568596 532884 568608
rect 532752 568568 532884 568596
rect 532752 568556 532758 568568
rect 532878 568556 532884 568568
rect 532936 568556 532942 568608
rect 524414 568528 524420 568540
rect 524375 568500 524420 568528
rect 524414 568488 524420 568500
rect 524472 568488 524478 568540
rect 3510 567196 3516 567248
rect 3568 567236 3574 567248
rect 33778 567236 33784 567248
rect 3568 567208 33784 567236
rect 3568 567196 3574 567208
rect 33778 567196 33784 567208
rect 33836 567196 33842 567248
rect 503806 565836 503812 565888
rect 503864 565876 503870 565888
rect 511718 565876 511724 565888
rect 503864 565848 511724 565876
rect 503864 565836 503870 565848
rect 511718 565836 511724 565848
rect 511776 565836 511782 565888
rect 503806 563048 503812 563100
rect 503864 563088 503870 563100
rect 574094 563088 574100 563100
rect 503864 563060 574100 563088
rect 503864 563048 503870 563060
rect 574094 563048 574100 563060
rect 574152 563048 574158 563100
rect 70302 558900 70308 558952
rect 70360 558940 70366 558952
rect 78674 558940 78680 558952
rect 70360 558912 78680 558940
rect 70360 558900 70366 558912
rect 78674 558900 78680 558912
rect 78732 558900 78738 558952
rect 532418 558900 532424 558952
rect 532476 558940 532482 558952
rect 532510 558940 532516 558952
rect 532476 558912 532516 558940
rect 532476 558900 532482 558912
rect 532510 558900 532516 558912
rect 532568 558900 532574 558952
rect 504910 556248 504916 556300
rect 504968 556288 504974 556300
rect 536834 556288 536840 556300
rect 504968 556260 536840 556288
rect 504968 556248 504974 556260
rect 536834 556248 536840 556260
rect 536892 556248 536898 556300
rect 529198 556180 529204 556232
rect 529256 556220 529262 556232
rect 580166 556220 580172 556232
rect 529256 556192 580172 556220
rect 529256 556180 529262 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 532510 553256 532516 553308
rect 532568 553296 532574 553308
rect 532878 553296 532884 553308
rect 532568 553268 532884 553296
rect 532568 553256 532574 553268
rect 532878 553256 532884 553268
rect 532936 553256 532942 553308
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 42150 552072 42156 552084
rect 3200 552044 42156 552072
rect 3200 552032 3206 552044
rect 42150 552032 42156 552044
rect 42208 552032 42214 552084
rect 504818 552032 504824 552084
rect 504876 552072 504882 552084
rect 507394 552072 507400 552084
rect 504876 552044 507400 552072
rect 504876 552032 504882 552044
rect 507394 552032 507400 552044
rect 507452 552032 507458 552084
rect 524417 550647 524475 550653
rect 524417 550613 524429 550647
rect 524463 550644 524475 550647
rect 524598 550644 524604 550656
rect 524463 550616 524604 550644
rect 524463 550613 524475 550616
rect 524417 550607 524475 550613
rect 524598 550604 524604 550616
rect 524656 550604 524662 550656
rect 505002 549312 505008 549364
rect 505060 549352 505066 549364
rect 508590 549352 508596 549364
rect 505060 549324 508596 549352
rect 505060 549312 505066 549324
rect 508590 549312 508596 549324
rect 508648 549312 508654 549364
rect 529934 545164 529940 545216
rect 529992 545204 529998 545216
rect 531958 545204 531964 545216
rect 529992 545176 531964 545204
rect 529992 545164 529998 545176
rect 531958 545164 531964 545176
rect 532016 545164 532022 545216
rect 524414 543736 524420 543788
rect 524472 543776 524478 543788
rect 524598 543776 524604 543788
rect 524472 543748 524604 543776
rect 524472 543736 524478 543748
rect 524598 543736 524604 543748
rect 524656 543736 524662 543788
rect 532694 540948 532700 541000
rect 532752 540988 532758 541000
rect 532970 540988 532976 541000
rect 532752 540960 532976 540988
rect 532752 540948 532758 540960
rect 532970 540948 532976 540960
rect 533028 540948 533034 541000
rect 3510 538228 3516 538280
rect 3568 538268 3574 538280
rect 9398 538268 9404 538280
rect 3568 538240 9404 538268
rect 3568 538228 3574 538240
rect 9398 538228 9404 538240
rect 9456 538228 9462 538280
rect 503346 534012 503352 534064
rect 503404 534052 503410 534064
rect 580166 534052 580172 534064
rect 503404 534024 580172 534052
rect 503404 534012 503410 534024
rect 580166 534012 580172 534024
rect 580224 534012 580230 534064
rect 82814 529904 82820 529916
rect 82775 529876 82820 529904
rect 82814 529864 82820 529876
rect 82872 529864 82878 529916
rect 505002 527144 505008 527196
rect 505060 527184 505066 527196
rect 510154 527184 510160 527196
rect 505060 527156 510160 527184
rect 505060 527144 505066 527156
rect 510154 527144 510160 527156
rect 510212 527144 510218 527196
rect 532694 521636 532700 521688
rect 532752 521676 532758 521688
rect 532878 521676 532884 521688
rect 532752 521648 532884 521676
rect 532752 521636 532758 521648
rect 532878 521636 532884 521648
rect 532936 521636 532942 521688
rect 82817 520319 82875 520325
rect 82817 520285 82829 520319
rect 82863 520316 82875 520319
rect 82906 520316 82912 520328
rect 82863 520288 82912 520316
rect 82863 520285 82875 520288
rect 82817 520279 82875 520285
rect 82906 520276 82912 520288
rect 82964 520276 82970 520328
rect 503714 514700 503720 514752
rect 503772 514740 503778 514752
rect 503898 514740 503904 514752
rect 503772 514712 503904 514740
rect 503772 514700 503778 514712
rect 503898 514700 503904 514712
rect 503956 514700 503962 514752
rect 504450 510552 504456 510604
rect 504508 510592 504514 510604
rect 580166 510592 580172 510604
rect 504508 510564 580172 510592
rect 504508 510552 504514 510564
rect 580166 510552 580172 510564
rect 580224 510552 580230 510604
rect 2866 509260 2872 509312
rect 2924 509300 2930 509312
rect 17218 509300 17224 509312
rect 2924 509272 17224 509300
rect 2924 509260 2930 509272
rect 17218 509260 17224 509272
rect 17276 509260 17282 509312
rect 503714 505112 503720 505164
rect 503772 505152 503778 505164
rect 503898 505152 503904 505164
rect 503772 505124 503904 505152
rect 503772 505112 503778 505124
rect 503898 505112 503904 505124
rect 503956 505112 503962 505164
rect 532694 502324 532700 502376
rect 532752 502364 532758 502376
rect 532878 502364 532884 502376
rect 532752 502336 532884 502364
rect 532752 502324 532758 502336
rect 532878 502324 532884 502336
rect 532936 502324 532942 502376
rect 82814 501032 82820 501084
rect 82872 501032 82878 501084
rect 82832 501004 82860 501032
rect 82906 501004 82912 501016
rect 82832 500976 82912 501004
rect 82906 500964 82912 500976
rect 82964 500964 82970 501016
rect 82814 500936 82820 500948
rect 82775 500908 82820 500936
rect 82814 500896 82820 500908
rect 82872 500896 82878 500948
rect 501966 499468 501972 499520
rect 502024 499508 502030 499520
rect 579982 499508 579988 499520
rect 502024 499480 579988 499508
rect 502024 499468 502030 499480
rect 579982 499468 579988 499480
rect 580040 499468 580046 499520
rect 3510 496748 3516 496800
rect 3568 496788 3574 496800
rect 80698 496788 80704 496800
rect 3568 496760 80704 496788
rect 3568 496748 3574 496760
rect 80698 496748 80704 496760
rect 80756 496748 80762 496800
rect 505002 492668 505008 492720
rect 505060 492708 505066 492720
rect 510246 492708 510252 492720
rect 505060 492680 510252 492708
rect 505060 492668 505066 492680
rect 510246 492668 510252 492680
rect 510304 492668 510310 492720
rect 532694 492600 532700 492652
rect 532752 492640 532758 492652
rect 532878 492640 532884 492652
rect 532752 492612 532884 492640
rect 532752 492600 532758 492612
rect 532878 492600 532884 492612
rect 532936 492600 532942 492652
rect 82814 491348 82820 491360
rect 82775 491320 82820 491348
rect 82814 491308 82820 491320
rect 82872 491308 82878 491360
rect 504450 485800 504456 485852
rect 504508 485840 504514 485852
rect 504508 485812 506520 485840
rect 504508 485800 504514 485812
rect 506492 485772 506520 485812
rect 519538 485800 519544 485852
rect 519596 485840 519602 485852
rect 580166 485840 580172 485852
rect 519596 485812 580172 485840
rect 519596 485800 519602 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 511626 485772 511632 485784
rect 506492 485744 511632 485772
rect 511626 485732 511632 485744
rect 511684 485732 511690 485784
rect 3326 481516 3332 481568
rect 3384 481556 3390 481568
rect 8754 481556 8760 481568
rect 3384 481528 8760 481556
rect 3384 481516 3390 481528
rect 8754 481516 8760 481528
rect 8812 481516 8818 481568
rect 505002 478864 505008 478916
rect 505060 478904 505066 478916
rect 513374 478904 513380 478916
rect 505060 478876 513380 478904
rect 505060 478864 505066 478876
rect 513374 478864 513380 478876
rect 513432 478864 513438 478916
rect 8846 478796 8852 478848
rect 8904 478836 8910 478848
rect 77570 478836 77576 478848
rect 8904 478808 77576 478836
rect 8904 478796 8910 478808
rect 77570 478796 77576 478808
rect 77628 478796 77634 478848
rect 503714 475736 503720 475788
rect 503772 475776 503778 475788
rect 504082 475776 504088 475788
rect 503772 475748 504088 475776
rect 503772 475736 503778 475748
rect 504082 475736 504088 475748
rect 504140 475736 504146 475788
rect 82630 474036 82636 474088
rect 82688 474076 82694 474088
rect 82906 474076 82912 474088
rect 82688 474048 82912 474076
rect 82688 474036 82694 474048
rect 82906 474036 82912 474048
rect 82964 474036 82970 474088
rect 524414 471968 524420 471980
rect 524375 471940 524420 471968
rect 524414 471928 524420 471940
rect 524472 471928 524478 471980
rect 503530 470568 503536 470620
rect 503588 470608 503594 470620
rect 531958 470608 531964 470620
rect 503588 470580 531964 470608
rect 503588 470568 503594 470580
rect 531958 470568 531964 470580
rect 532016 470568 532022 470620
rect 524414 462448 524420 462460
rect 524375 462420 524420 462448
rect 524414 462408 524420 462420
rect 524472 462408 524478 462460
rect 505738 462340 505744 462392
rect 505796 462380 505802 462392
rect 580166 462380 580172 462392
rect 505796 462352 580172 462380
rect 505796 462340 505802 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 503714 461388 503720 461440
rect 503772 461428 503778 461440
rect 504082 461428 504088 461440
rect 503772 461400 504088 461428
rect 503772 461388 503778 461400
rect 504082 461388 504088 461400
rect 504140 461388 504146 461440
rect 503714 456424 503720 456476
rect 503772 456464 503778 456476
rect 504082 456464 504088 456476
rect 503772 456436 504088 456464
rect 503772 456424 503778 456436
rect 504082 456424 504088 456436
rect 504140 456424 504146 456476
rect 504542 454044 504548 454096
rect 504600 454084 504606 454096
rect 510338 454084 510344 454096
rect 504600 454056 510344 454084
rect 504600 454044 504606 454056
rect 510338 454044 510344 454056
rect 510396 454044 510402 454096
rect 524414 452588 524420 452600
rect 524375 452560 524420 452588
rect 524414 452548 524420 452560
rect 524472 452548 524478 452600
rect 82630 450168 82636 450220
rect 82688 450208 82694 450220
rect 82906 450208 82912 450220
rect 82688 450180 82912 450208
rect 82688 450168 82694 450180
rect 82906 450168 82912 450180
rect 82964 450168 82970 450220
rect 82817 447831 82875 447837
rect 82817 447797 82829 447831
rect 82863 447828 82875 447831
rect 82998 447828 83004 447840
rect 82863 447800 83004 447828
rect 82863 447797 82875 447800
rect 82817 447791 82875 447797
rect 82998 447788 83004 447800
rect 83056 447788 83062 447840
rect 503714 447108 503720 447160
rect 503772 447148 503778 447160
rect 504082 447148 504088 447160
rect 503772 447120 504088 447148
rect 503772 447108 503778 447120
rect 504082 447108 504088 447120
rect 504140 447108 504146 447160
rect 524414 443000 524420 443012
rect 524375 442972 524420 443000
rect 524414 442960 524420 442972
rect 524472 442960 524478 443012
rect 82725 442935 82783 442941
rect 82725 442901 82737 442935
rect 82771 442932 82783 442935
rect 82814 442932 82820 442944
rect 82771 442904 82820 442932
rect 82771 442901 82783 442904
rect 82725 442895 82783 442901
rect 82814 442892 82820 442904
rect 82872 442892 82878 442944
rect 82814 442144 82820 442196
rect 82872 442184 82878 442196
rect 82998 442184 83004 442196
rect 82872 442156 83004 442184
rect 82872 442144 82878 442156
rect 82998 442144 83004 442156
rect 83056 442144 83062 442196
rect 503254 440172 503260 440224
rect 503312 440212 503318 440224
rect 579982 440212 579988 440224
rect 503312 440184 579988 440212
rect 503312 440172 503318 440184
rect 579982 440172 579988 440184
rect 580040 440172 580046 440224
rect 82817 439535 82875 439541
rect 82817 439501 82829 439535
rect 82863 439532 82875 439535
rect 82906 439532 82912 439544
rect 82863 439504 82912 439532
rect 82863 439501 82875 439504
rect 82817 439495 82875 439501
rect 82906 439492 82912 439504
rect 82964 439492 82970 439544
rect 82725 438175 82783 438181
rect 82725 438141 82737 438175
rect 82771 438172 82783 438175
rect 82814 438172 82820 438184
rect 82771 438144 82820 438172
rect 82771 438141 82783 438144
rect 82725 438135 82783 438141
rect 82814 438132 82820 438144
rect 82872 438132 82878 438184
rect 503714 437384 503720 437436
rect 503772 437424 503778 437436
rect 504266 437424 504272 437436
rect 503772 437396 504272 437424
rect 503772 437384 503778 437396
rect 504266 437384 504272 437396
rect 504324 437384 504330 437436
rect 12342 436092 12348 436144
rect 12400 436132 12406 436144
rect 75086 436132 75092 436144
rect 12400 436104 75092 436132
rect 12400 436092 12406 436104
rect 75086 436092 75092 436104
rect 75144 436092 75150 436144
rect 524414 433276 524420 433288
rect 524375 433248 524420 433276
rect 524414 433236 524420 433248
rect 524472 433236 524478 433288
rect 38562 427796 38568 427848
rect 38620 427836 38626 427848
rect 77570 427836 77576 427848
rect 38620 427808 77576 427836
rect 38620 427796 38626 427808
rect 77570 427796 77576 427808
rect 77628 427796 77634 427848
rect 503714 427796 503720 427848
rect 503772 427836 503778 427848
rect 504266 427836 504272 427848
rect 503772 427808 504272 427836
rect 503772 427796 503778 427808
rect 504266 427796 504272 427808
rect 504324 427796 504330 427848
rect 2958 424192 2964 424244
rect 3016 424232 3022 424244
rect 9582 424232 9588 424244
rect 3016 424204 9588 424232
rect 3016 424192 3022 424204
rect 9582 424192 9588 424204
rect 9640 424192 9646 424244
rect 524414 423688 524420 423700
rect 524375 423660 524420 423688
rect 524414 423648 524420 423660
rect 524472 423648 524478 423700
rect 82814 423620 82820 423632
rect 82775 423592 82820 423620
rect 82814 423580 82820 423592
rect 82872 423580 82878 423632
rect 82906 423008 82912 423020
rect 82867 422980 82912 423008
rect 82906 422968 82912 422980
rect 82964 422968 82970 423020
rect 82906 418996 82912 419008
rect 82867 418968 82912 418996
rect 82906 418956 82912 418968
rect 82964 418956 82970 419008
rect 503254 418208 503260 418260
rect 503312 418248 503318 418260
rect 505462 418248 505468 418260
rect 503312 418220 505468 418248
rect 503312 418208 503318 418220
rect 505462 418208 505468 418220
rect 505520 418208 505526 418260
rect 503714 418072 503720 418124
rect 503772 418112 503778 418124
rect 504266 418112 504272 418124
rect 503772 418084 504272 418112
rect 503772 418072 503778 418084
rect 504266 418072 504272 418084
rect 504324 418072 504330 418124
rect 514018 416712 514024 416764
rect 514076 416752 514082 416764
rect 580166 416752 580172 416764
rect 514076 416724 580172 416752
rect 514076 416712 514082 416724
rect 580166 416712 580172 416724
rect 580224 416712 580230 416764
rect 82814 414032 82820 414044
rect 82775 414004 82820 414032
rect 82814 413992 82820 414004
rect 82872 413992 82878 414044
rect 524414 413964 524420 413976
rect 524375 413936 524420 413964
rect 524414 413924 524420 413936
rect 524472 413924 524478 413976
rect 503714 408484 503720 408536
rect 503772 408524 503778 408536
rect 504266 408524 504272 408536
rect 503772 408496 504272 408524
rect 503772 408484 503778 408496
rect 504266 408484 504272 408496
rect 504324 408484 504330 408536
rect 4890 407124 4896 407176
rect 4948 407164 4954 407176
rect 77662 407164 77668 407176
rect 4948 407136 77668 407164
rect 4948 407124 4954 407136
rect 77662 407124 77668 407136
rect 77720 407124 77726 407176
rect 82906 406280 82912 406292
rect 82867 406252 82912 406280
rect 82906 406240 82912 406252
rect 82964 406240 82970 406292
rect 524414 404376 524420 404388
rect 524375 404348 524420 404376
rect 524414 404336 524420 404348
rect 524472 404336 524478 404388
rect 505002 402772 505008 402824
rect 505060 402812 505066 402824
rect 505922 402812 505928 402824
rect 505060 402784 505928 402812
rect 505060 402772 505066 402784
rect 505922 402772 505928 402784
rect 505980 402772 505986 402824
rect 82725 400707 82783 400713
rect 82725 400673 82737 400707
rect 82771 400704 82783 400707
rect 82998 400704 83004 400716
rect 82771 400676 83004 400704
rect 82771 400673 82783 400676
rect 82725 400667 82783 400673
rect 82998 400664 83004 400676
rect 83056 400664 83062 400716
rect 82817 400367 82875 400373
rect 82817 400333 82829 400367
rect 82863 400364 82875 400367
rect 82998 400364 83004 400376
rect 82863 400336 83004 400364
rect 82863 400333 82875 400336
rect 82817 400327 82875 400333
rect 82998 400324 83004 400336
rect 83056 400324 83062 400376
rect 77846 400188 77852 400240
rect 77904 400228 77910 400240
rect 78766 400228 78772 400240
rect 77904 400200 78772 400228
rect 77904 400188 77910 400200
rect 78766 400188 78772 400200
rect 78824 400188 78830 400240
rect 82725 400231 82783 400237
rect 82725 400197 82737 400231
rect 82771 400228 82783 400231
rect 82998 400228 83004 400240
rect 82771 400200 83004 400228
rect 82771 400197 82783 400200
rect 82725 400191 82783 400197
rect 82998 400188 83004 400200
rect 83056 400188 83062 400240
rect 82817 399551 82875 399557
rect 82817 399517 82829 399551
rect 82863 399548 82875 399551
rect 82998 399548 83004 399560
rect 82863 399520 83004 399548
rect 82863 399517 82875 399520
rect 82817 399511 82875 399517
rect 82998 399508 83004 399520
rect 83056 399508 83062 399560
rect 3326 394680 3332 394732
rect 3384 394720 3390 394732
rect 9582 394720 9588 394732
rect 3384 394692 9588 394720
rect 3384 394680 3390 394692
rect 9582 394680 9588 394692
rect 9640 394680 9646 394732
rect 524414 394652 524420 394664
rect 524375 394624 524420 394652
rect 524414 394612 524420 394624
rect 524472 394612 524478 394664
rect 69658 393320 69664 393372
rect 69716 393360 69722 393372
rect 78766 393360 78772 393372
rect 69716 393332 78772 393360
rect 69716 393320 69722 393332
rect 78766 393320 78772 393332
rect 78824 393320 78830 393372
rect 503162 393252 503168 393304
rect 503220 393292 503226 393304
rect 579706 393292 579712 393304
rect 503220 393264 579712 393292
rect 503220 393252 503226 393264
rect 579706 393252 579712 393264
rect 579764 393252 579770 393304
rect 504542 390532 504548 390584
rect 504600 390572 504606 390584
rect 508682 390572 508688 390584
rect 504600 390544 508688 390572
rect 504600 390532 504606 390544
rect 508682 390532 508688 390544
rect 508740 390532 508746 390584
rect 82078 387948 82084 388000
rect 82136 387988 82142 388000
rect 82262 387988 82268 388000
rect 82136 387960 82268 387988
rect 82136 387948 82142 387960
rect 82262 387948 82268 387960
rect 82320 387948 82326 388000
rect 82909 387991 82967 387997
rect 82909 387957 82921 387991
rect 82955 387957 82967 387991
rect 82909 387951 82967 387957
rect 82924 387920 82952 387951
rect 82998 387920 83004 387932
rect 82924 387892 83004 387920
rect 82998 387880 83004 387892
rect 83056 387880 83062 387932
rect 524414 385064 524420 385076
rect 524375 385036 524420 385064
rect 524414 385024 524420 385036
rect 524472 385024 524478 385076
rect 82814 384996 82820 385008
rect 82775 384968 82820 384996
rect 82814 384956 82820 384968
rect 82872 384956 82878 385008
rect 3050 379516 3056 379568
rect 3108 379556 3114 379568
rect 21358 379556 21364 379568
rect 3108 379528 21364 379556
rect 3108 379516 3114 379528
rect 21358 379516 21364 379528
rect 21416 379516 21422 379568
rect 49602 379516 49608 379568
rect 49660 379556 49666 379568
rect 77570 379556 77576 379568
rect 49660 379528 77576 379556
rect 49660 379516 49666 379528
rect 77570 379516 77576 379528
rect 77628 379516 77634 379568
rect 504174 376728 504180 376780
rect 504232 376768 504238 376780
rect 507762 376768 507768 376780
rect 504232 376740 507768 376768
rect 504232 376728 504238 376740
rect 507762 376728 507768 376740
rect 507820 376728 507826 376780
rect 82814 375476 82820 375488
rect 82775 375448 82820 375476
rect 82814 375436 82820 375448
rect 82872 375436 82878 375488
rect 82262 375300 82268 375352
rect 82320 375340 82326 375352
rect 82814 375340 82820 375352
rect 82320 375312 82820 375340
rect 82320 375300 82326 375312
rect 82814 375300 82820 375312
rect 82872 375300 82878 375352
rect 524414 375340 524420 375352
rect 524375 375312 524420 375340
rect 524414 375300 524420 375312
rect 524472 375300 524478 375352
rect 82998 372756 83004 372768
rect 82832 372728 83004 372756
rect 10962 372580 10968 372632
rect 11020 372620 11026 372632
rect 77570 372620 77576 372632
rect 11020 372592 77576 372620
rect 11020 372580 11026 372592
rect 77570 372580 77576 372592
rect 77628 372580 77634 372632
rect 82832 372484 82860 372728
rect 82998 372716 83004 372728
rect 83056 372716 83062 372768
rect 82909 372623 82967 372629
rect 82909 372589 82921 372623
rect 82955 372620 82967 372623
rect 82998 372620 83004 372632
rect 82955 372592 83004 372620
rect 82955 372589 82967 372592
rect 82909 372583 82967 372589
rect 82998 372580 83004 372592
rect 83056 372580 83062 372632
rect 504174 372580 504180 372632
rect 504232 372620 504238 372632
rect 540238 372620 540244 372632
rect 504232 372592 540244 372620
rect 504232 372580 504238 372592
rect 540238 372580 540244 372592
rect 540296 372580 540302 372632
rect 82998 372484 83004 372496
rect 82832 372456 83004 372484
rect 82998 372444 83004 372456
rect 83056 372444 83062 372496
rect 82262 370852 82268 370864
rect 82223 370824 82268 370852
rect 82262 370812 82268 370824
rect 82320 370812 82326 370864
rect 504542 369860 504548 369912
rect 504600 369900 504606 369912
rect 511810 369900 511816 369912
rect 504600 369872 511816 369900
rect 504600 369860 504606 369872
rect 511810 369860 511816 369872
rect 511868 369860 511874 369912
rect 82909 369359 82967 369365
rect 82909 369325 82921 369359
rect 82955 369356 82967 369359
rect 82998 369356 83004 369368
rect 82955 369328 83004 369356
rect 82955 369325 82967 369328
rect 82909 369319 82967 369325
rect 82998 369316 83004 369328
rect 83056 369316 83062 369368
rect 507578 368500 507584 368552
rect 507636 368540 507642 368552
rect 580166 368540 580172 368552
rect 507636 368512 580172 368540
rect 507636 368500 507642 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 82538 366800 82544 366852
rect 82596 366840 82602 366852
rect 82906 366840 82912 366852
rect 82596 366812 82912 366840
rect 82596 366800 82602 366812
rect 82906 366800 82912 366812
rect 82964 366800 82970 366852
rect 3602 365712 3608 365764
rect 3660 365752 3666 365764
rect 42242 365752 42248 365764
rect 3660 365724 42248 365752
rect 3660 365712 3666 365724
rect 42242 365712 42248 365724
rect 42300 365712 42306 365764
rect 524414 365752 524420 365764
rect 524375 365724 524420 365752
rect 524414 365712 524420 365724
rect 524472 365712 524478 365764
rect 82265 365279 82323 365285
rect 82265 365245 82277 365279
rect 82311 365276 82323 365279
rect 82538 365276 82544 365288
rect 82311 365248 82544 365276
rect 82311 365245 82323 365248
rect 82265 365239 82323 365245
rect 82538 365236 82544 365248
rect 82596 365236 82602 365288
rect 21358 362856 21364 362908
rect 21416 362896 21422 362908
rect 77570 362896 77576 362908
rect 21416 362868 77576 362896
rect 21416 362856 21422 362868
rect 77570 362856 77576 362868
rect 77628 362856 77634 362908
rect 504542 362788 504548 362840
rect 504600 362828 504606 362840
rect 508774 362828 508780 362840
rect 504600 362800 508780 362828
rect 504600 362788 504606 362800
rect 508774 362788 508780 362800
rect 508832 362788 508838 362840
rect 505922 358028 505928 358080
rect 505980 358068 505986 358080
rect 506106 358068 506112 358080
rect 505980 358040 506112 358068
rect 505980 358028 505986 358040
rect 506106 358028 506112 358040
rect 506164 358028 506170 358080
rect 33870 357416 33876 357468
rect 33928 357456 33934 357468
rect 74166 357456 74172 357468
rect 33928 357428 74172 357456
rect 33928 357416 33934 357428
rect 74166 357416 74172 357428
rect 74224 357416 74230 357468
rect 524414 356028 524420 356040
rect 524375 356000 524420 356028
rect 524414 355988 524420 356000
rect 524472 355988 524478 356040
rect 504174 351908 504180 351960
rect 504232 351948 504238 351960
rect 508774 351948 508780 351960
rect 504232 351920 508780 351948
rect 504232 351908 504238 351920
rect 508774 351908 508780 351920
rect 508832 351908 508838 351960
rect 524414 346440 524420 346452
rect 524375 346412 524420 346440
rect 524414 346400 524420 346412
rect 524472 346400 524478 346452
rect 507670 346332 507676 346384
rect 507728 346372 507734 346384
rect 580166 346372 580172 346384
rect 507728 346344 580172 346372
rect 507728 346332 507734 346344
rect 580166 346332 580172 346344
rect 580224 346332 580230 346384
rect 82814 344972 82820 345024
rect 82872 345012 82878 345024
rect 82906 345012 82912 345024
rect 82872 344984 82912 345012
rect 82872 344972 82878 344984
rect 82906 344972 82912 344984
rect 82964 344972 82970 345024
rect 63402 343612 63408 343664
rect 63460 343652 63466 343664
rect 77570 343652 77576 343664
rect 63460 343624 77576 343652
rect 63460 343612 63466 343624
rect 77570 343612 77576 343624
rect 77628 343612 77634 343664
rect 15930 342184 15936 342236
rect 15988 342224 15994 342236
rect 73614 342224 73620 342236
rect 15988 342196 73620 342224
rect 15988 342184 15994 342196
rect 73614 342184 73620 342196
rect 73672 342184 73678 342236
rect 503438 340892 503444 340944
rect 503496 340932 503502 340944
rect 511902 340932 511908 340944
rect 503496 340904 511908 340932
rect 503496 340892 503502 340904
rect 511902 340892 511908 340904
rect 511960 340892 511966 340944
rect 505922 339668 505928 339720
rect 505980 339708 505986 339720
rect 506198 339708 506204 339720
rect 505980 339680 506204 339708
rect 505980 339668 505986 339680
rect 506198 339668 506204 339680
rect 506256 339668 506262 339720
rect 2958 336744 2964 336796
rect 3016 336784 3022 336796
rect 8846 336784 8852 336796
rect 3016 336756 8852 336784
rect 3016 336744 3022 336756
rect 8846 336744 8852 336756
rect 8904 336744 8910 336796
rect 524414 336716 524420 336728
rect 524375 336688 524420 336716
rect 524414 336676 524420 336688
rect 524472 336676 524478 336728
rect 17218 333888 17224 333940
rect 17276 333928 17282 333940
rect 76466 333928 76472 333940
rect 17276 333900 76472 333928
rect 17276 333888 17282 333900
rect 76466 333888 76472 333900
rect 76524 333888 76530 333940
rect 17218 329808 17224 329860
rect 17276 329848 17282 329860
rect 77570 329848 77576 329860
rect 17276 329820 77576 329848
rect 17276 329808 17282 329820
rect 77570 329808 77576 329820
rect 77628 329808 77634 329860
rect 504450 329808 504456 329860
rect 504508 329848 504514 329860
rect 538858 329848 538864 329860
rect 504508 329820 538864 329848
rect 504508 329808 504514 329820
rect 538858 329808 538864 329820
rect 538916 329808 538922 329860
rect 82906 328556 82912 328568
rect 82832 328528 82912 328556
rect 82832 328500 82860 328528
rect 82906 328516 82912 328528
rect 82964 328516 82970 328568
rect 82814 328448 82820 328500
rect 82872 328448 82878 328500
rect 79594 327972 79600 328024
rect 79652 328012 79658 328024
rect 79962 328012 79968 328024
rect 79652 327984 79968 328012
rect 79652 327972 79658 327984
rect 79962 327972 79968 327984
rect 80020 327972 80026 328024
rect 524414 327128 524420 327140
rect 524375 327100 524420 327128
rect 524414 327088 524420 327100
rect 524472 327088 524478 327140
rect 82909 326995 82967 327001
rect 82909 326961 82921 326995
rect 82955 326992 82967 326995
rect 82998 326992 83004 327004
rect 82955 326964 83004 326992
rect 82955 326961 82967 326964
rect 82909 326955 82967 326961
rect 82998 326952 83004 326964
rect 83056 326952 83062 327004
rect 3326 324232 3332 324284
rect 3384 324272 3390 324284
rect 75270 324272 75276 324284
rect 3384 324244 75276 324272
rect 3384 324232 3390 324244
rect 75270 324232 75276 324244
rect 75328 324232 75334 324284
rect 504450 324232 504456 324284
rect 504508 324272 504514 324284
rect 529198 324272 529204 324284
rect 504508 324244 529204 324272
rect 504508 324232 504514 324244
rect 529198 324232 529204 324244
rect 529256 324232 529262 324284
rect 505830 322872 505836 322924
rect 505888 322912 505894 322924
rect 580166 322912 580172 322924
rect 505888 322884 580172 322912
rect 505888 322872 505894 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 79594 319104 79600 319116
rect 79555 319076 79600 319104
rect 79594 319064 79600 319076
rect 79652 319064 79658 319116
rect 506014 318792 506020 318844
rect 506072 318832 506078 318844
rect 506290 318832 506296 318844
rect 506072 318804 506296 318832
rect 506072 318792 506078 318804
rect 506290 318792 506296 318804
rect 506348 318792 506354 318844
rect 82909 317475 82967 317481
rect 82909 317441 82921 317475
rect 82955 317472 82967 317475
rect 82998 317472 83004 317484
rect 82955 317444 83004 317472
rect 82955 317441 82967 317444
rect 82909 317435 82967 317441
rect 82998 317432 83004 317444
rect 83056 317432 83062 317484
rect 524414 317404 524420 317416
rect 524375 317376 524420 317404
rect 524414 317364 524420 317376
rect 524472 317364 524478 317416
rect 82722 316072 82728 316124
rect 82780 316112 82786 316124
rect 82906 316112 82912 316124
rect 82780 316084 82912 316112
rect 82780 316072 82786 316084
rect 82906 316072 82912 316084
rect 82964 316072 82970 316124
rect 82630 315936 82636 315988
rect 82688 315976 82694 315988
rect 82906 315976 82912 315988
rect 82688 315948 82912 315976
rect 82688 315936 82694 315948
rect 82906 315936 82912 315948
rect 82964 315936 82970 315988
rect 82725 313327 82783 313333
rect 82725 313293 82737 313327
rect 82771 313324 82783 313327
rect 82814 313324 82820 313336
rect 82771 313296 82820 313324
rect 82771 313293 82783 313296
rect 82725 313287 82783 313293
rect 82814 313284 82820 313296
rect 82872 313284 82878 313336
rect 82817 311355 82875 311361
rect 82817 311321 82829 311355
rect 82863 311352 82875 311355
rect 82906 311352 82912 311364
rect 82863 311324 82912 311352
rect 82863 311321 82875 311324
rect 82817 311315 82875 311321
rect 82906 311312 82912 311324
rect 82964 311312 82970 311364
rect 82909 310879 82967 310885
rect 82909 310845 82921 310879
rect 82955 310876 82967 310879
rect 82998 310876 83004 310888
rect 82955 310848 83004 310876
rect 82955 310845 82967 310848
rect 82909 310839 82967 310845
rect 82998 310836 83004 310848
rect 83056 310836 83062 310888
rect 82630 310700 82636 310752
rect 82688 310740 82694 310752
rect 82998 310740 83004 310752
rect 82688 310712 83004 310740
rect 82688 310700 82694 310712
rect 82998 310700 83004 310712
rect 83056 310700 83062 310752
rect 82909 310607 82967 310613
rect 82909 310573 82921 310607
rect 82955 310604 82967 310607
rect 82998 310604 83004 310616
rect 82955 310576 83004 310604
rect 82955 310573 82967 310576
rect 82909 310567 82967 310573
rect 82998 310564 83004 310576
rect 83056 310564 83062 310616
rect 70210 309136 70216 309188
rect 70268 309176 70274 309188
rect 77570 309176 77576 309188
rect 70268 309148 77576 309176
rect 70268 309136 70274 309148
rect 77570 309136 77576 309148
rect 77628 309136 77634 309188
rect 504450 309136 504456 309188
rect 504508 309176 504514 309188
rect 506750 309176 506756 309188
rect 504508 309148 506756 309176
rect 504508 309136 504514 309148
rect 506750 309136 506756 309148
rect 506808 309136 506814 309188
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 17218 309108 17224 309120
rect 3384 309080 17224 309108
rect 3384 309068 3390 309080
rect 17218 309068 17224 309080
rect 17276 309068 17282 309120
rect 82725 309111 82783 309117
rect 82725 309077 82737 309111
rect 82771 309108 82783 309111
rect 82814 309108 82820 309120
rect 82771 309080 82820 309108
rect 82771 309077 82783 309080
rect 82725 309071 82783 309077
rect 82814 309068 82820 309080
rect 82872 309068 82878 309120
rect 524414 307816 524420 307828
rect 524375 307788 524420 307816
rect 524414 307776 524420 307788
rect 524472 307776 524478 307828
rect 507026 307096 507032 307148
rect 507084 307136 507090 307148
rect 507670 307136 507676 307148
rect 507084 307108 507676 307136
rect 507084 307096 507090 307108
rect 507670 307096 507676 307108
rect 507728 307096 507734 307148
rect 504450 306348 504456 306400
rect 504508 306388 504514 306400
rect 564434 306388 564440 306400
rect 504508 306360 564440 306388
rect 504508 306348 504514 306360
rect 564434 306348 564440 306360
rect 564492 306348 564498 306400
rect 82725 303331 82783 303337
rect 82725 303297 82737 303331
rect 82771 303328 82783 303331
rect 82814 303328 82820 303340
rect 82771 303300 82820 303328
rect 82771 303297 82783 303300
rect 82725 303291 82783 303297
rect 82814 303288 82820 303300
rect 82872 303288 82878 303340
rect 82906 303288 82912 303340
rect 82964 303328 82970 303340
rect 82964 303300 83044 303328
rect 82964 303288 82970 303300
rect 82906 303056 82912 303068
rect 82867 303028 82912 303056
rect 82906 303016 82912 303028
rect 82964 303016 82970 303068
rect 82725 302923 82783 302929
rect 82725 302889 82737 302923
rect 82771 302920 82783 302923
rect 82814 302920 82820 302932
rect 82771 302892 82820 302920
rect 82771 302889 82783 302892
rect 82725 302883 82783 302889
rect 82814 302880 82820 302892
rect 82872 302880 82878 302932
rect 82906 302880 82912 302932
rect 82964 302920 82970 302932
rect 83016 302920 83044 303300
rect 82964 302892 83044 302920
rect 82964 302880 82970 302892
rect 82630 300500 82636 300552
rect 82688 300540 82694 300552
rect 82906 300540 82912 300552
rect 82688 300512 82912 300540
rect 82688 300500 82694 300512
rect 82906 300500 82912 300512
rect 82964 300500 82970 300552
rect 511718 299412 511724 299464
rect 511776 299452 511782 299464
rect 580166 299452 580172 299464
rect 511776 299424 580172 299452
rect 511776 299412 511782 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 82722 298256 82728 298308
rect 82780 298296 82786 298308
rect 82817 298299 82875 298305
rect 82817 298296 82829 298299
rect 82780 298268 82829 298296
rect 82780 298256 82786 298268
rect 82817 298265 82829 298268
rect 82863 298265 82875 298299
rect 82817 298259 82875 298265
rect 82725 298095 82783 298101
rect 82725 298061 82737 298095
rect 82771 298092 82783 298095
rect 82814 298092 82820 298104
rect 82771 298064 82820 298092
rect 82771 298061 82783 298064
rect 82725 298055 82783 298061
rect 82814 298052 82820 298064
rect 82872 298052 82878 298104
rect 524414 298092 524420 298104
rect 524375 298064 524420 298092
rect 524414 298052 524420 298064
rect 524472 298052 524478 298104
rect 504450 296624 504456 296676
rect 504508 296664 504514 296676
rect 519538 296664 519544 296676
rect 504508 296636 519544 296664
rect 504508 296624 504514 296636
rect 519538 296624 519544 296636
rect 519596 296624 519602 296676
rect 79318 296080 79324 296132
rect 79376 296120 79382 296132
rect 79505 296123 79563 296129
rect 79505 296120 79517 296123
rect 79376 296092 79517 296120
rect 79376 296080 79382 296092
rect 79505 296089 79517 296092
rect 79551 296089 79563 296123
rect 79505 296083 79563 296089
rect 3234 294720 3240 294772
rect 3292 294760 3298 294772
rect 9490 294760 9496 294772
rect 3292 294732 9496 294760
rect 3292 294720 3298 294732
rect 9490 294720 9496 294732
rect 9548 294720 9554 294772
rect 82817 293403 82875 293409
rect 82817 293369 82829 293403
rect 82863 293400 82875 293403
rect 82906 293400 82912 293412
rect 82863 293372 82912 293400
rect 82863 293369 82875 293372
rect 82817 293363 82875 293369
rect 82906 293360 82912 293372
rect 82964 293360 82970 293412
rect 82814 291864 82820 291916
rect 82872 291904 82878 291916
rect 82909 291907 82967 291913
rect 82909 291904 82921 291907
rect 82872 291876 82921 291904
rect 82872 291864 82878 291876
rect 82909 291873 82921 291876
rect 82955 291873 82967 291907
rect 82909 291867 82967 291873
rect 82906 291768 82912 291780
rect 82867 291740 82912 291768
rect 82906 291728 82912 291740
rect 82964 291728 82970 291780
rect 501966 290272 501972 290284
rect 501927 290244 501972 290272
rect 501966 290232 501972 290244
rect 502024 290232 502030 290284
rect 82817 288847 82875 288853
rect 82817 288813 82829 288847
rect 82863 288844 82875 288847
rect 82906 288844 82912 288856
rect 82863 288816 82912 288844
rect 82863 288813 82875 288816
rect 82817 288807 82875 288813
rect 82906 288804 82912 288816
rect 82964 288804 82970 288856
rect 524414 288436 524420 288448
rect 524375 288408 524420 288436
rect 524414 288396 524420 288408
rect 524472 288396 524478 288448
rect 82906 287756 82912 287768
rect 82867 287728 82912 287756
rect 82906 287716 82912 287728
rect 82964 287716 82970 287768
rect 79318 287348 79324 287360
rect 79279 287320 79324 287348
rect 79318 287308 79324 287320
rect 79376 287308 79382 287360
rect 79778 287348 79784 287360
rect 79739 287320 79784 287348
rect 79778 287308 79784 287320
rect 79836 287308 79842 287360
rect 82725 286399 82783 286405
rect 82725 286365 82737 286399
rect 82771 286396 82783 286399
rect 82814 286396 82820 286408
rect 82771 286368 82820 286396
rect 82771 286365 82783 286368
rect 82725 286359 82783 286365
rect 82814 286356 82820 286368
rect 82872 286356 82878 286408
rect 82722 286220 82728 286272
rect 82780 286260 82786 286272
rect 82906 286260 82912 286272
rect 82780 286232 82912 286260
rect 82780 286220 82786 286232
rect 82906 286220 82912 286232
rect 82964 286220 82970 286272
rect 77570 284588 77576 284640
rect 77628 284628 77634 284640
rect 82630 284628 82636 284640
rect 77628 284600 82636 284628
rect 77628 284588 77634 284600
rect 82630 284588 82636 284600
rect 82688 284588 82694 284640
rect 82906 282248 82912 282260
rect 82867 282220 82912 282248
rect 82906 282208 82912 282220
rect 82964 282208 82970 282260
rect 501877 282251 501935 282257
rect 501877 282217 501889 282251
rect 501923 282248 501935 282251
rect 501966 282248 501972 282260
rect 501923 282220 501972 282248
rect 501923 282217 501935 282220
rect 501877 282211 501935 282217
rect 501966 282208 501972 282220
rect 502024 282208 502030 282260
rect 79321 280823 79379 280829
rect 79321 280789 79333 280823
rect 79367 280820 79379 280823
rect 79594 280820 79600 280832
rect 79367 280792 79600 280820
rect 79367 280789 79379 280792
rect 79321 280783 79379 280789
rect 79594 280780 79600 280792
rect 79652 280780 79658 280832
rect 79778 280820 79784 280832
rect 79739 280792 79784 280820
rect 79778 280780 79784 280792
rect 79836 280780 79842 280832
rect 57882 280168 57888 280220
rect 57940 280208 57946 280220
rect 75638 280208 75644 280220
rect 57940 280180 75644 280208
rect 57940 280168 57946 280180
rect 75638 280168 75644 280180
rect 75696 280168 75702 280220
rect 14458 278672 14464 278724
rect 14516 278712 14522 278724
rect 75454 278712 75460 278724
rect 14516 278684 75460 278712
rect 14516 278672 14522 278684
rect 75454 278672 75460 278684
rect 75512 278672 75518 278724
rect 501785 278443 501843 278449
rect 501785 278409 501797 278443
rect 501831 278440 501843 278443
rect 501966 278440 501972 278452
rect 501831 278412 501972 278440
rect 501831 278409 501843 278412
rect 501785 278403 501843 278409
rect 501966 278400 501972 278412
rect 502024 278400 502030 278452
rect 501966 278264 501972 278316
rect 502024 278304 502030 278316
rect 502242 278304 502248 278316
rect 502024 278276 502248 278304
rect 502024 278264 502030 278276
rect 502242 278264 502248 278276
rect 502300 278264 502306 278316
rect 506106 277856 506112 277908
rect 506164 277896 506170 277908
rect 506201 277899 506259 277905
rect 506201 277896 506213 277899
rect 506164 277868 506213 277896
rect 506164 277856 506170 277868
rect 506201 277865 506213 277868
rect 506247 277865 506259 277899
rect 506201 277859 506259 277865
rect 502242 277788 502248 277840
rect 502300 277828 502306 277840
rect 509050 277828 509056 277840
rect 502300 277800 509056 277828
rect 502300 277788 502306 277800
rect 509050 277788 509056 277800
rect 509108 277788 509114 277840
rect 502242 277584 502248 277636
rect 502300 277624 502306 277636
rect 504174 277624 504180 277636
rect 502300 277596 504180 277624
rect 502300 277584 502306 277596
rect 504174 277584 504180 277596
rect 504232 277584 504238 277636
rect 82906 277420 82912 277432
rect 82867 277392 82912 277420
rect 82906 277380 82912 277392
rect 82964 277380 82970 277432
rect 560938 275952 560944 276004
rect 560996 275992 561002 276004
rect 580166 275992 580172 276004
rect 560996 275964 580172 275992
rect 560996 275952 561002 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 504174 274660 504180 274712
rect 504232 274700 504238 274712
rect 545114 274700 545120 274712
rect 504232 274672 545120 274700
rect 504232 274660 504238 274672
rect 545114 274660 545120 274672
rect 545172 274660 545178 274712
rect 504174 274524 504180 274576
rect 504232 274564 504238 274576
rect 504726 274564 504732 274576
rect 504232 274536 504732 274564
rect 504232 274524 504238 274536
rect 504726 274524 504732 274536
rect 504784 274524 504790 274576
rect 82906 273816 82912 273828
rect 82867 273788 82912 273816
rect 82906 273776 82912 273788
rect 82964 273776 82970 273828
rect 501966 272756 501972 272808
rect 502024 272796 502030 272808
rect 502061 272799 502119 272805
rect 502061 272796 502073 272799
rect 502024 272768 502073 272796
rect 502024 272756 502030 272768
rect 502061 272765 502073 272768
rect 502107 272765 502119 272799
rect 502061 272759 502119 272765
rect 501877 272663 501935 272669
rect 501877 272629 501889 272663
rect 501923 272660 501935 272663
rect 501966 272660 501972 272672
rect 501923 272632 501972 272660
rect 501923 272629 501935 272632
rect 501877 272623 501935 272629
rect 501966 272620 501972 272632
rect 502024 272620 502030 272672
rect 501966 272524 501972 272536
rect 501927 272496 501972 272524
rect 501966 272484 501972 272496
rect 502024 272484 502030 272536
rect 501785 272391 501843 272397
rect 501785 272357 501797 272391
rect 501831 272388 501843 272391
rect 501966 272388 501972 272400
rect 501831 272360 501972 272388
rect 501831 272357 501843 272360
rect 501785 272351 501843 272357
rect 501966 272348 501972 272360
rect 502024 272348 502030 272400
rect 79594 272144 79600 272196
rect 79652 272184 79658 272196
rect 79962 272184 79968 272196
rect 79652 272156 79968 272184
rect 79652 272144 79658 272156
rect 79962 272144 79968 272156
rect 80020 272144 80026 272196
rect 501966 270852 501972 270904
rect 502024 270892 502030 270904
rect 502061 270895 502119 270901
rect 502061 270892 502073 270895
rect 502024 270864 502073 270892
rect 502024 270852 502030 270864
rect 502061 270861 502073 270864
rect 502107 270861 502119 270895
rect 502061 270855 502119 270861
rect 501509 270419 501567 270425
rect 501509 270385 501521 270419
rect 501555 270416 501567 270419
rect 501966 270416 501972 270428
rect 501555 270388 501972 270416
rect 501555 270385 501567 270388
rect 501509 270379 501567 270385
rect 501966 270376 501972 270388
rect 502024 270376 502030 270428
rect 82817 269807 82875 269813
rect 82817 269773 82829 269807
rect 82863 269804 82875 269807
rect 82906 269804 82912 269816
rect 82863 269776 82912 269804
rect 82863 269773 82875 269776
rect 82817 269767 82875 269773
rect 82906 269764 82912 269776
rect 82964 269764 82970 269816
rect 82633 269603 82691 269609
rect 82633 269569 82645 269603
rect 82679 269600 82691 269603
rect 82906 269600 82912 269612
rect 82679 269572 82912 269600
rect 82679 269569 82691 269572
rect 82633 269563 82691 269569
rect 82906 269560 82912 269572
rect 82964 269560 82970 269612
rect 82725 269467 82783 269473
rect 82725 269433 82737 269467
rect 82771 269464 82783 269467
rect 82906 269464 82912 269476
rect 82771 269436 82912 269464
rect 82771 269433 82783 269436
rect 82725 269427 82783 269433
rect 82906 269424 82912 269436
rect 82964 269424 82970 269476
rect 524414 269084 524420 269136
rect 524472 269124 524478 269136
rect 524598 269124 524604 269136
rect 524472 269096 524604 269124
rect 524472 269084 524478 269096
rect 524598 269084 524604 269096
rect 524656 269084 524662 269136
rect 501966 267112 501972 267164
rect 502024 267152 502030 267164
rect 503622 267152 503628 267164
rect 502024 267124 503628 267152
rect 502024 267112 502030 267124
rect 503622 267112 503628 267124
rect 503680 267112 503686 267164
rect 501601 267019 501659 267025
rect 501601 266985 501613 267019
rect 501647 267016 501659 267019
rect 501966 267016 501972 267028
rect 501647 266988 501972 267016
rect 501647 266985 501659 266988
rect 501601 266979 501659 266985
rect 501966 266976 501972 266988
rect 502024 266976 502030 267028
rect 82630 265888 82636 265940
rect 82688 265928 82694 265940
rect 82998 265928 83004 265940
rect 82688 265900 83004 265928
rect 82688 265888 82694 265900
rect 82998 265888 83004 265900
rect 83056 265888 83062 265940
rect 82725 265863 82783 265869
rect 82725 265829 82737 265863
rect 82771 265860 82783 265863
rect 82906 265860 82912 265872
rect 82771 265832 82912 265860
rect 82771 265829 82783 265832
rect 82725 265823 82783 265829
rect 82906 265820 82912 265832
rect 82964 265820 82970 265872
rect 82633 265455 82691 265461
rect 82633 265421 82645 265455
rect 82679 265452 82691 265455
rect 82906 265452 82912 265464
rect 82679 265424 82912 265452
rect 82679 265421 82691 265424
rect 82633 265415 82691 265421
rect 82906 265412 82912 265424
rect 82964 265412 82970 265464
rect 2958 264936 2964 264988
rect 3016 264976 3022 264988
rect 77294 264976 77300 264988
rect 3016 264948 77300 264976
rect 3016 264936 3022 264948
rect 77294 264936 77300 264948
rect 77352 264936 77358 264988
rect 506201 264843 506259 264849
rect 506201 264809 506213 264843
rect 506247 264840 506259 264843
rect 506290 264840 506296 264852
rect 506247 264812 506296 264840
rect 506247 264809 506259 264812
rect 506201 264803 506259 264809
rect 506290 264800 506296 264812
rect 506348 264800 506354 264852
rect 79410 264596 79416 264648
rect 79468 264636 79474 264648
rect 80054 264636 80060 264648
rect 79468 264608 80060 264636
rect 79468 264596 79474 264608
rect 80054 264596 80060 264608
rect 80112 264596 80118 264648
rect 82817 263551 82875 263557
rect 82817 263517 82829 263551
rect 82863 263548 82875 263551
rect 82906 263548 82912 263560
rect 82863 263520 82912 263548
rect 82863 263517 82875 263520
rect 82817 263511 82875 263517
rect 82906 263508 82912 263520
rect 82964 263508 82970 263560
rect 82906 263140 82912 263152
rect 82867 263112 82912 263140
rect 82906 263100 82912 263112
rect 82964 263100 82970 263152
rect 79594 260448 79600 260500
rect 79652 260488 79658 260500
rect 79962 260488 79968 260500
rect 79652 260460 79968 260488
rect 79652 260448 79658 260460
rect 79962 260448 79968 260460
rect 80020 260448 80026 260500
rect 505830 254844 505836 254856
rect 505791 254816 505836 254844
rect 505830 254804 505836 254816
rect 505888 254804 505894 254856
rect 501601 254643 501659 254649
rect 501601 254609 501613 254643
rect 501647 254640 501659 254643
rect 503346 254640 503352 254652
rect 501647 254612 503352 254640
rect 501647 254609 501659 254612
rect 501601 254603 501659 254609
rect 503346 254600 503352 254612
rect 503404 254600 503410 254652
rect 501509 253215 501567 253221
rect 501509 253181 501521 253215
rect 501555 253212 501567 253215
rect 503438 253212 503444 253224
rect 501555 253184 503444 253212
rect 501555 253181 501567 253184
rect 501509 253175 501567 253181
rect 503438 253172 503444 253184
rect 503496 253172 503502 253224
rect 503438 252968 503444 253020
rect 503496 253008 503502 253020
rect 504637 253011 504695 253017
rect 504637 253008 504649 253011
rect 503496 252980 504649 253008
rect 503496 252968 503502 252980
rect 504637 252977 504649 252980
rect 504683 252977 504695 253011
rect 504637 252971 504695 252977
rect 79594 252560 79600 252612
rect 79652 252600 79658 252612
rect 79962 252600 79968 252612
rect 79652 252572 79968 252600
rect 79652 252560 79658 252572
rect 79962 252560 79968 252572
rect 80020 252560 80026 252612
rect 505833 251311 505891 251317
rect 505833 251277 505845 251311
rect 505879 251308 505891 251311
rect 506198 251308 506204 251320
rect 505879 251280 506204 251308
rect 505879 251277 505891 251280
rect 505833 251271 505891 251277
rect 506198 251268 506204 251280
rect 506256 251268 506262 251320
rect 3326 251200 3332 251252
rect 3384 251240 3390 251252
rect 14458 251240 14464 251252
rect 3384 251212 14464 251240
rect 3384 251200 3390 251212
rect 14458 251200 14464 251212
rect 14516 251200 14522 251252
rect 506106 251200 506112 251252
rect 506164 251240 506170 251252
rect 580166 251240 580172 251252
rect 506164 251212 580172 251240
rect 506164 251200 506170 251212
rect 580166 251200 580172 251212
rect 580224 251200 580230 251252
rect 505922 249772 505928 249824
rect 505980 249812 505986 249824
rect 506290 249812 506296 249824
rect 505980 249784 506296 249812
rect 505980 249772 505986 249784
rect 506290 249772 506296 249784
rect 506348 249772 506354 249824
rect 524414 249772 524420 249824
rect 524472 249812 524478 249824
rect 524598 249812 524604 249824
rect 524472 249784 524604 249812
rect 524472 249772 524478 249784
rect 524598 249772 524604 249784
rect 524656 249772 524662 249824
rect 41322 248412 41328 248464
rect 41380 248452 41386 248464
rect 76006 248452 76012 248464
rect 41380 248424 76012 248452
rect 41380 248412 41386 248424
rect 76006 248412 76012 248424
rect 76064 248412 76070 248464
rect 82906 248452 82912 248464
rect 82867 248424 82912 248452
rect 82906 248412 82912 248424
rect 82964 248412 82970 248464
rect 504634 246412 504640 246424
rect 504595 246384 504640 246412
rect 504634 246372 504640 246384
rect 504692 246372 504698 246424
rect 82817 246347 82875 246353
rect 82817 246313 82829 246347
rect 82863 246344 82875 246347
rect 82906 246344 82912 246356
rect 82863 246316 82912 246344
rect 82863 246313 82875 246316
rect 82817 246307 82875 246313
rect 82906 246304 82912 246316
rect 82964 246304 82970 246356
rect 82725 246211 82783 246217
rect 82725 246177 82737 246211
rect 82771 246208 82783 246211
rect 82814 246208 82820 246220
rect 82771 246180 82820 246208
rect 82771 246177 82783 246180
rect 82725 246171 82783 246177
rect 82814 246168 82820 246180
rect 82872 246168 82878 246220
rect 82633 245939 82691 245945
rect 82633 245905 82645 245939
rect 82679 245936 82691 245939
rect 82906 245936 82912 245948
rect 82679 245908 82912 245936
rect 82679 245905 82691 245908
rect 82633 245899 82691 245905
rect 82906 245896 82912 245908
rect 82964 245896 82970 245948
rect 503438 245284 503444 245336
rect 503496 245284 503502 245336
rect 503456 245200 503484 245284
rect 503438 245148 503444 245200
rect 503496 245148 503502 245200
rect 82906 245052 82912 245064
rect 82867 245024 82912 245052
rect 82906 245012 82912 245024
rect 82964 245012 82970 245064
rect 82725 244987 82783 244993
rect 82725 244953 82737 244987
rect 82771 244984 82783 244987
rect 82814 244984 82820 244996
rect 82771 244956 82820 244984
rect 82771 244953 82783 244956
rect 82725 244947 82783 244953
rect 82814 244944 82820 244956
rect 82872 244944 82878 244996
rect 82722 243788 82728 243840
rect 82780 243828 82786 243840
rect 82906 243828 82912 243840
rect 82780 243800 82912 243828
rect 82780 243788 82786 243800
rect 82906 243788 82912 243800
rect 82964 243788 82970 243840
rect 82633 243695 82691 243701
rect 82633 243661 82645 243695
rect 82679 243692 82691 243695
rect 82906 243692 82912 243704
rect 82679 243664 82912 243692
rect 82679 243661 82691 243664
rect 82633 243655 82691 243661
rect 82906 243652 82912 243664
rect 82964 243652 82970 243704
rect 82817 243559 82875 243565
rect 82817 243525 82829 243559
rect 82863 243556 82875 243559
rect 82906 243556 82912 243568
rect 82863 243528 82912 243556
rect 82863 243525 82875 243528
rect 82817 243519 82875 243525
rect 82906 243516 82912 243528
rect 82964 243516 82970 243568
rect 503346 242088 503352 242140
rect 503404 242088 503410 242140
rect 503364 241924 503392 242088
rect 503438 241924 503444 241936
rect 503364 241896 503444 241924
rect 503438 241884 503444 241896
rect 503496 241884 503502 241936
rect 503622 241584 503628 241596
rect 503583 241556 503628 241584
rect 503622 241544 503628 241556
rect 503680 241544 503686 241596
rect 514588 238972 524460 239000
rect 503438 238824 503444 238876
rect 503496 238864 503502 238876
rect 514588 238864 514616 238972
rect 503496 238836 514616 238864
rect 524432 238864 524460 238972
rect 539502 238960 539508 239012
rect 539560 239000 539566 239012
rect 549254 239000 549260 239012
rect 539560 238972 549260 239000
rect 539560 238960 539566 238972
rect 549254 238960 549260 238972
rect 549312 238960 549318 239012
rect 529860 238904 529980 238932
rect 529860 238864 529888 238904
rect 529952 238876 529980 238904
rect 524432 238836 529888 238864
rect 503496 238824 503502 238836
rect 529934 238824 529940 238876
rect 529992 238824 529998 238876
rect 82814 238796 82820 238808
rect 82740 238768 82820 238796
rect 82740 238660 82768 238768
rect 82814 238756 82820 238768
rect 82872 238756 82878 238808
rect 82906 238728 82912 238740
rect 82867 238700 82912 238728
rect 82906 238688 82912 238700
rect 82964 238688 82970 238740
rect 82814 238660 82820 238672
rect 82740 238632 82820 238660
rect 82814 238620 82820 238632
rect 82872 238620 82878 238672
rect 81529 238119 81587 238125
rect 81529 238085 81541 238119
rect 81575 238116 81587 238119
rect 82446 238116 82452 238128
rect 81575 238088 82452 238116
rect 81575 238085 81587 238088
rect 81529 238079 81587 238085
rect 82446 238076 82452 238088
rect 82504 238076 82510 238128
rect 79410 237464 79416 237516
rect 79468 237504 79474 237516
rect 79962 237504 79968 237516
rect 79468 237476 79968 237504
rect 79468 237464 79474 237476
rect 79962 237464 79968 237476
rect 80020 237464 80026 237516
rect 3234 237328 3240 237380
rect 3292 237368 3298 237380
rect 77754 237368 77760 237380
rect 3292 237340 77760 237368
rect 3292 237328 3298 237340
rect 77754 237328 77760 237340
rect 77812 237328 77818 237380
rect 504634 235968 504640 236020
rect 504692 236008 504698 236020
rect 508866 236008 508872 236020
rect 504692 235980 508872 236008
rect 504692 235968 504698 235980
rect 508866 235968 508872 235980
rect 508924 235968 508930 236020
rect 503622 235220 503628 235272
rect 503680 235260 503686 235272
rect 504634 235260 504640 235272
rect 503680 235232 504640 235260
rect 503680 235220 503686 235232
rect 504634 235220 504640 235232
rect 504692 235220 504698 235272
rect 82446 235016 82452 235068
rect 82504 235056 82510 235068
rect 82722 235056 82728 235068
rect 82504 235028 82728 235056
rect 82504 235016 82510 235028
rect 82722 235016 82728 235028
rect 82780 235016 82786 235068
rect 81434 233696 81440 233708
rect 81395 233668 81440 233696
rect 81434 233656 81440 233668
rect 81492 233656 81498 233708
rect 501601 233631 501659 233637
rect 501601 233597 501613 233631
rect 501647 233628 501659 233631
rect 503530 233628 503536 233640
rect 501647 233600 503536 233628
rect 501647 233597 501659 233600
rect 501601 233591 501659 233597
rect 503530 233588 503536 233600
rect 503588 233588 503594 233640
rect 82817 233087 82875 233093
rect 82817 233053 82829 233087
rect 82863 233084 82875 233087
rect 83182 233084 83188 233096
rect 82863 233056 83188 233084
rect 82863 233053 82875 233056
rect 82817 233047 82875 233053
rect 83182 233044 83188 233056
rect 83240 233044 83246 233096
rect 82725 233019 82783 233025
rect 82725 232985 82737 233019
rect 82771 233016 82783 233019
rect 82906 233016 82912 233028
rect 82771 232988 82912 233016
rect 82771 232985 82783 232988
rect 82725 232979 82783 232985
rect 82906 232976 82912 232988
rect 82964 232976 82970 233028
rect 82722 232840 82728 232892
rect 82780 232880 82786 232892
rect 82906 232880 82912 232892
rect 82780 232852 82912 232880
rect 82780 232840 82786 232852
rect 82906 232840 82912 232852
rect 82964 232840 82970 232892
rect 82630 232608 82636 232620
rect 82591 232580 82636 232608
rect 82630 232568 82636 232580
rect 82688 232568 82694 232620
rect 81434 230596 81440 230648
rect 81492 230636 81498 230648
rect 81492 230608 81537 230636
rect 81492 230596 81498 230608
rect 524414 230460 524420 230512
rect 524472 230500 524478 230512
rect 524598 230500 524604 230512
rect 524472 230472 524604 230500
rect 524472 230460 524478 230472
rect 524598 230460 524604 230472
rect 524656 230460 524662 230512
rect 81434 229236 81440 229288
rect 81492 229276 81498 229288
rect 81529 229279 81587 229285
rect 81529 229276 81541 229279
rect 81492 229248 81541 229276
rect 81492 229236 81498 229248
rect 81529 229245 81541 229248
rect 81575 229245 81587 229279
rect 81529 229239 81587 229245
rect 507486 229032 507492 229084
rect 507544 229072 507550 229084
rect 580166 229072 580172 229084
rect 507544 229044 580172 229072
rect 507544 229032 507550 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 82722 228964 82728 229016
rect 82780 229004 82786 229016
rect 82906 229004 82912 229016
rect 82780 228976 82912 229004
rect 82780 228964 82786 228976
rect 82906 228964 82912 228976
rect 82964 228964 82970 229016
rect 82725 228871 82783 228877
rect 82725 228837 82737 228871
rect 82771 228868 82783 228871
rect 82906 228868 82912 228880
rect 82771 228840 82912 228868
rect 82771 228837 82783 228840
rect 82725 228831 82783 228837
rect 82906 228828 82912 228840
rect 82964 228828 82970 228880
rect 81434 227876 81440 227928
rect 81492 227916 81498 227928
rect 82633 227919 82691 227925
rect 82633 227916 82645 227919
rect 81492 227888 82645 227916
rect 81492 227876 81498 227888
rect 82633 227885 82645 227888
rect 82679 227885 82691 227919
rect 82633 227879 82691 227885
rect 503622 227440 503628 227452
rect 503583 227412 503628 227440
rect 503622 227400 503628 227412
rect 503680 227400 503686 227452
rect 82906 226556 82912 226568
rect 82867 226528 82912 226556
rect 82906 226516 82912 226528
rect 82964 226516 82970 226568
rect 79410 225632 79416 225684
rect 79468 225672 79474 225684
rect 79594 225672 79600 225684
rect 79468 225644 79600 225672
rect 79468 225632 79474 225644
rect 79594 225632 79600 225644
rect 79652 225632 79658 225684
rect 82817 225675 82875 225681
rect 82817 225641 82829 225675
rect 82863 225672 82875 225675
rect 82906 225672 82912 225684
rect 82863 225644 82912 225672
rect 82863 225641 82875 225644
rect 82817 225635 82875 225641
rect 82906 225632 82912 225644
rect 82964 225632 82970 225684
rect 503438 225496 503444 225548
rect 503496 225536 503502 225548
rect 503533 225539 503591 225545
rect 503533 225536 503545 225539
rect 503496 225508 503545 225536
rect 503496 225496 503502 225508
rect 503533 225505 503545 225508
rect 503579 225505 503591 225539
rect 503533 225499 503591 225505
rect 503438 224952 503444 225004
rect 503496 224992 503502 225004
rect 519538 224992 519544 225004
rect 503496 224964 519544 224992
rect 503496 224952 503502 224964
rect 519538 224952 519544 224964
rect 519596 224952 519602 225004
rect 505830 224612 505836 224664
rect 505888 224652 505894 224664
rect 506290 224652 506296 224664
rect 505888 224624 506296 224652
rect 505888 224612 505894 224624
rect 506290 224612 506296 224624
rect 506348 224612 506354 224664
rect 505922 224068 505928 224120
rect 505980 224108 505986 224120
rect 506382 224108 506388 224120
rect 505980 224080 506388 224108
rect 505980 224068 505986 224080
rect 506382 224068 506388 224080
rect 506440 224068 506446 224120
rect 3326 223524 3332 223576
rect 3384 223564 3390 223576
rect 10686 223564 10692 223576
rect 3384 223536 10692 223564
rect 3384 223524 3390 223536
rect 10686 223524 10692 223536
rect 10744 223524 10750 223576
rect 503438 221824 503444 221876
rect 503496 221864 503502 221876
rect 508958 221864 508964 221876
rect 503496 221836 508964 221864
rect 503496 221824 503502 221836
rect 508958 221824 508964 221836
rect 509016 221824 509022 221876
rect 503622 221524 503628 221536
rect 503583 221496 503628 221524
rect 503622 221484 503628 221496
rect 503680 221484 503686 221536
rect 503622 221252 503628 221264
rect 503583 221224 503628 221252
rect 503622 221212 503628 221224
rect 503680 221212 503686 221264
rect 82906 220844 82912 220856
rect 82867 220816 82912 220844
rect 82906 220804 82912 220816
rect 82964 220804 82970 220856
rect 501509 220235 501567 220241
rect 501509 220201 501521 220235
rect 501555 220232 501567 220235
rect 503622 220232 503628 220244
rect 501555 220204 503628 220232
rect 501555 220201 501567 220204
rect 501509 220195 501567 220201
rect 503622 220192 503628 220204
rect 503680 220192 503686 220244
rect 501601 220031 501659 220037
rect 501601 219997 501613 220031
rect 501647 220028 501659 220031
rect 503530 220028 503536 220040
rect 501647 220000 503536 220028
rect 501647 219997 501659 220000
rect 501601 219991 501659 219997
rect 503530 219988 503536 220000
rect 503588 219988 503594 220040
rect 503530 219688 503536 219700
rect 503491 219660 503536 219688
rect 503530 219648 503536 219660
rect 503588 219648 503594 219700
rect 82906 219484 82912 219496
rect 82867 219456 82912 219484
rect 82906 219444 82912 219456
rect 82964 219444 82970 219496
rect 506198 217988 506204 218000
rect 506159 217960 506204 217988
rect 506198 217948 506204 217960
rect 506256 217948 506262 218000
rect 509050 217948 509056 218000
rect 509108 217988 509114 218000
rect 580166 217988 580172 218000
rect 509108 217960 580172 217988
rect 509108 217948 509114 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 77754 216656 77760 216708
rect 77812 216696 77818 216708
rect 80330 216696 80336 216708
rect 77812 216668 80336 216696
rect 77812 216656 77818 216668
rect 80330 216656 80336 216668
rect 80388 216656 80394 216708
rect 79594 215228 79600 215280
rect 79652 215268 79658 215280
rect 79962 215268 79968 215280
rect 79652 215240 79968 215268
rect 79652 215228 79658 215240
rect 79962 215228 79968 215240
rect 80020 215228 80026 215280
rect 505922 214344 505928 214396
rect 505980 214384 505986 214396
rect 506382 214384 506388 214396
rect 505980 214356 506388 214384
rect 505980 214344 505986 214356
rect 506382 214344 506388 214356
rect 506440 214344 506446 214396
rect 81526 213392 81532 213444
rect 81584 213432 81590 213444
rect 82722 213432 82728 213444
rect 81584 213404 82728 213432
rect 81584 213392 81590 213404
rect 82722 213392 82728 213404
rect 82780 213392 82786 213444
rect 505830 212304 505836 212356
rect 505888 212344 505894 212356
rect 506290 212344 506296 212356
rect 505888 212316 506296 212344
rect 505888 212304 505894 212316
rect 506290 212304 506296 212316
rect 506348 212304 506354 212356
rect 506201 212211 506259 212217
rect 506201 212177 506213 212211
rect 506247 212208 506259 212211
rect 506290 212208 506296 212220
rect 506247 212180 506296 212208
rect 506247 212177 506259 212180
rect 506201 212171 506259 212177
rect 506290 212168 506296 212180
rect 506348 212168 506354 212220
rect 82906 211148 82912 211200
rect 82964 211188 82970 211200
rect 82998 211188 83004 211200
rect 82964 211160 83004 211188
rect 82964 211148 82970 211160
rect 82998 211148 83004 211160
rect 83056 211148 83062 211200
rect 501509 210783 501567 210789
rect 501509 210749 501521 210783
rect 501555 210780 501567 210783
rect 503622 210780 503628 210792
rect 501555 210752 503628 210780
rect 501555 210749 501567 210752
rect 501509 210743 501567 210749
rect 503622 210740 503628 210752
rect 503680 210740 503686 210792
rect 82630 209488 82636 209500
rect 82591 209460 82636 209488
rect 82630 209448 82636 209460
rect 82688 209448 82694 209500
rect 502150 209352 502156 209364
rect 502111 209324 502156 209352
rect 502150 209312 502156 209324
rect 502208 209312 502214 209364
rect 3142 208292 3148 208344
rect 3200 208332 3206 208344
rect 10594 208332 10600 208344
rect 3200 208304 10600 208332
rect 3200 208292 3206 208304
rect 10594 208292 10600 208304
rect 10652 208292 10658 208344
rect 501601 207859 501659 207865
rect 501601 207825 501613 207859
rect 501647 207856 501659 207859
rect 504818 207856 504824 207868
rect 501647 207828 504824 207856
rect 501647 207825 501659 207828
rect 501601 207819 501659 207825
rect 504818 207816 504824 207828
rect 504876 207816 504882 207868
rect 503622 207000 503628 207052
rect 503680 207040 503686 207052
rect 572714 207040 572720 207052
rect 503680 207012 572720 207040
rect 503680 207000 503686 207012
rect 572714 207000 572720 207012
rect 572772 207000 572778 207052
rect 79594 205640 79600 205692
rect 79652 205680 79658 205692
rect 79962 205680 79968 205692
rect 79652 205652 79968 205680
rect 79652 205640 79658 205652
rect 79962 205640 79968 205652
rect 80020 205640 80026 205692
rect 503530 204864 503536 204876
rect 503491 204836 503536 204864
rect 503530 204824 503536 204836
rect 503588 204824 503594 204876
rect 506198 204280 506204 204332
rect 506256 204320 506262 204332
rect 580166 204320 580172 204332
rect 506256 204292 580172 204320
rect 506256 204280 506262 204292
rect 580166 204280 580172 204292
rect 580224 204280 580230 204332
rect 505830 203940 505836 203992
rect 505888 203980 505894 203992
rect 506382 203980 506388 203992
rect 505888 203952 506388 203980
rect 505888 203940 505894 203952
rect 506382 203940 506388 203952
rect 506440 203940 506446 203992
rect 81526 202484 81532 202496
rect 81487 202456 81532 202484
rect 81526 202444 81532 202456
rect 81584 202444 81590 202496
rect 79134 202104 79140 202156
rect 79192 202144 79198 202156
rect 80330 202144 80336 202156
rect 79192 202116 80336 202144
rect 79192 202104 79198 202116
rect 80330 202104 80336 202116
rect 80388 202104 80394 202156
rect 81526 201764 81532 201816
rect 81584 201804 81590 201816
rect 82265 201807 82323 201813
rect 82265 201804 82277 201807
rect 81584 201776 82277 201804
rect 81584 201764 81590 201776
rect 82265 201773 82277 201776
rect 82311 201773 82323 201807
rect 82265 201767 82323 201773
rect 524414 201424 524420 201476
rect 524472 201464 524478 201476
rect 524598 201464 524604 201476
rect 524472 201436 524604 201464
rect 524472 201424 524478 201436
rect 524598 201424 524604 201436
rect 524656 201424 524662 201476
rect 81526 201220 81532 201272
rect 81584 201260 81590 201272
rect 82633 201263 82691 201269
rect 82633 201260 82645 201263
rect 81584 201232 82645 201260
rect 81584 201220 81590 201232
rect 82633 201229 82645 201232
rect 82679 201229 82691 201263
rect 82633 201223 82691 201229
rect 76466 200744 76472 200796
rect 76524 200784 76530 200796
rect 76926 200784 76932 200796
rect 76524 200756 76932 200784
rect 76524 200744 76530 200756
rect 76926 200744 76932 200756
rect 76984 200744 76990 200796
rect 81526 200268 81532 200320
rect 81584 200308 81590 200320
rect 82541 200311 82599 200317
rect 82541 200308 82553 200311
rect 81584 200280 82553 200308
rect 81584 200268 81590 200280
rect 82541 200277 82553 200280
rect 82587 200277 82599 200311
rect 82541 200271 82599 200277
rect 80330 200200 80336 200252
rect 80388 200240 80394 200252
rect 81434 200240 81440 200252
rect 80388 200212 81440 200240
rect 80388 200200 80394 200212
rect 81434 200200 81440 200212
rect 81492 200200 81498 200252
rect 81526 200172 81532 200184
rect 81487 200144 81532 200172
rect 81526 200132 81532 200144
rect 81584 200132 81590 200184
rect 505922 199628 505928 199640
rect 505883 199600 505928 199628
rect 505922 199588 505928 199600
rect 505980 199588 505986 199640
rect 76926 199520 76932 199572
rect 76984 199560 76990 199572
rect 77110 199560 77116 199572
rect 76984 199532 77116 199560
rect 76984 199520 76990 199532
rect 77110 199520 77116 199532
rect 77168 199520 77174 199572
rect 503622 199492 503628 199504
rect 503583 199464 503628 199492
rect 503622 199452 503628 199464
rect 503680 199452 503686 199504
rect 503533 199359 503591 199365
rect 503533 199325 503545 199359
rect 503579 199356 503591 199359
rect 503622 199356 503628 199368
rect 503579 199328 503628 199356
rect 503579 199325 503591 199328
rect 503533 199319 503591 199325
rect 503622 199316 503628 199328
rect 503680 199316 503686 199368
rect 502150 197724 502156 197736
rect 502111 197696 502156 197724
rect 502150 197684 502156 197696
rect 502208 197684 502214 197736
rect 79594 196800 79600 196852
rect 79652 196840 79658 196852
rect 79962 196840 79968 196852
rect 79652 196812 79968 196840
rect 79652 196800 79658 196812
rect 79962 196800 79968 196812
rect 80020 196800 80026 196852
rect 503530 196188 503536 196240
rect 503588 196228 503594 196240
rect 503625 196231 503683 196237
rect 503625 196228 503637 196231
rect 503588 196200 503637 196228
rect 503588 196188 503594 196200
rect 503625 196197 503637 196200
rect 503671 196197 503683 196231
rect 503625 196191 503683 196197
rect 504818 195984 504824 196036
rect 504876 196024 504882 196036
rect 509142 196024 509148 196036
rect 504876 195996 509148 196024
rect 504876 195984 504882 195996
rect 509142 195984 509148 195996
rect 509200 195984 509206 196036
rect 82817 195347 82875 195353
rect 82817 195313 82829 195347
rect 82863 195344 82875 195347
rect 82906 195344 82912 195356
rect 82863 195316 82912 195344
rect 82863 195313 82875 195316
rect 82817 195307 82875 195313
rect 82906 195304 82912 195316
rect 82964 195304 82970 195356
rect 82722 195276 82728 195288
rect 82683 195248 82728 195276
rect 82722 195236 82728 195248
rect 82780 195236 82786 195288
rect 82906 195208 82912 195220
rect 82867 195180 82912 195208
rect 82906 195168 82912 195180
rect 82964 195168 82970 195220
rect 82722 195100 82728 195152
rect 82780 195140 82786 195152
rect 82817 195143 82875 195149
rect 82817 195140 82829 195143
rect 82780 195112 82829 195140
rect 82780 195100 82786 195112
rect 82817 195109 82829 195112
rect 82863 195109 82875 195143
rect 82817 195103 82875 195109
rect 82173 195075 82231 195081
rect 82173 195041 82185 195075
rect 82219 195072 82231 195075
rect 82630 195072 82636 195084
rect 82219 195044 82636 195072
rect 82219 195041 82231 195044
rect 82173 195035 82231 195041
rect 82630 195032 82636 195044
rect 82688 195032 82694 195084
rect 82449 194939 82507 194945
rect 82449 194905 82461 194939
rect 82495 194936 82507 194939
rect 82630 194936 82636 194948
rect 82495 194908 82636 194936
rect 82495 194905 82507 194908
rect 82449 194899 82507 194905
rect 82630 194896 82636 194908
rect 82688 194896 82694 194948
rect 82817 194939 82875 194945
rect 82817 194905 82829 194939
rect 82863 194936 82875 194939
rect 82906 194936 82912 194948
rect 82863 194908 82912 194936
rect 82863 194905 82875 194908
rect 82817 194899 82875 194905
rect 82906 194896 82912 194908
rect 82964 194896 82970 194948
rect 82081 194803 82139 194809
rect 82081 194769 82093 194803
rect 82127 194800 82139 194803
rect 82630 194800 82636 194812
rect 82127 194772 82636 194800
rect 82127 194769 82139 194772
rect 82081 194763 82139 194769
rect 82630 194760 82636 194772
rect 82688 194760 82694 194812
rect 82906 194800 82912 194812
rect 82867 194772 82912 194800
rect 82906 194760 82912 194772
rect 82964 194760 82970 194812
rect 503073 194395 503131 194401
rect 503073 194361 503085 194395
rect 503119 194392 503131 194395
rect 503530 194392 503536 194404
rect 503119 194364 503536 194392
rect 503119 194361 503131 194364
rect 503073 194355 503131 194361
rect 503530 194352 503536 194364
rect 503588 194352 503594 194404
rect 503070 192584 503076 192636
rect 503128 192624 503134 192636
rect 510522 192624 510528 192636
rect 503128 192596 510528 192624
rect 503128 192584 503134 192596
rect 510522 192584 510528 192596
rect 510580 192584 510586 192636
rect 81526 192420 81532 192432
rect 81487 192392 81532 192420
rect 81526 192380 81532 192392
rect 81584 192380 81590 192432
rect 81526 192176 81532 192228
rect 81584 192216 81590 192228
rect 82906 192216 82912 192228
rect 81584 192188 82912 192216
rect 81584 192176 81590 192188
rect 82906 192176 82912 192188
rect 82964 192176 82970 192228
rect 81526 191768 81532 191820
rect 81584 191808 81590 191820
rect 81621 191811 81679 191817
rect 81621 191808 81633 191811
rect 81584 191780 81633 191808
rect 81584 191768 81590 191780
rect 81621 191777 81633 191780
rect 81667 191777 81679 191811
rect 81621 191771 81679 191777
rect 82357 191267 82415 191273
rect 82357 191233 82369 191267
rect 82403 191264 82415 191267
rect 82630 191264 82636 191276
rect 82403 191236 82636 191264
rect 82403 191233 82415 191236
rect 82357 191227 82415 191233
rect 82630 191224 82636 191236
rect 82688 191224 82694 191276
rect 82541 191199 82599 191205
rect 82541 191196 82553 191199
rect 82004 191168 82553 191196
rect 76926 191088 76932 191140
rect 76984 191128 76990 191140
rect 77110 191128 77116 191140
rect 76984 191100 77116 191128
rect 76984 191088 76990 191100
rect 77110 191088 77116 191100
rect 77168 191088 77174 191140
rect 80238 191088 80244 191140
rect 80296 191128 80302 191140
rect 82004 191128 82032 191168
rect 82541 191165 82553 191168
rect 82587 191165 82599 191199
rect 82541 191159 82599 191165
rect 82630 191128 82636 191140
rect 80296 191100 82032 191128
rect 82591 191100 82636 191128
rect 80296 191088 80302 191100
rect 82630 191088 82636 191100
rect 82688 191088 82694 191140
rect 76466 190952 76472 191004
rect 76524 190992 76530 191004
rect 76926 190992 76932 191004
rect 76524 190964 76932 190992
rect 76524 190952 76530 190964
rect 76926 190952 76932 190964
rect 76984 190952 76990 191004
rect 82449 190995 82507 191001
rect 82449 190961 82461 190995
rect 82495 190992 82507 190995
rect 82630 190992 82636 191004
rect 82495 190964 82636 190992
rect 82495 190961 82507 190964
rect 82449 190955 82507 190961
rect 82630 190952 82636 190964
rect 82688 190952 82694 191004
rect 82538 190856 82544 190868
rect 82499 190828 82544 190856
rect 82538 190816 82544 190828
rect 82596 190816 82602 190868
rect 82173 190791 82231 190797
rect 82173 190757 82185 190791
rect 82219 190788 82231 190791
rect 82630 190788 82636 190800
rect 82219 190760 82636 190788
rect 82219 190757 82231 190760
rect 82173 190751 82231 190757
rect 82630 190748 82636 190760
rect 82688 190748 82694 190800
rect 505922 190788 505928 190800
rect 505883 190760 505928 190788
rect 505922 190748 505928 190760
rect 505980 190748 505986 190800
rect 81526 190680 81532 190732
rect 81584 190720 81590 190732
rect 82538 190720 82544 190732
rect 81584 190692 82544 190720
rect 81584 190680 81590 190692
rect 82538 190680 82544 190692
rect 82596 190680 82602 190732
rect 81529 190519 81587 190525
rect 81529 190485 81541 190519
rect 81575 190516 81587 190519
rect 82538 190516 82544 190528
rect 81575 190488 82544 190516
rect 81575 190485 81587 190488
rect 81529 190479 81587 190485
rect 82538 190476 82544 190488
rect 82596 190476 82602 190528
rect 503070 189700 503076 189712
rect 503031 189672 503076 189700
rect 503070 189660 503076 189672
rect 503128 189660 503134 189712
rect 82541 189091 82599 189097
rect 82541 189057 82553 189091
rect 82587 189057 82599 189091
rect 82541 189051 82599 189057
rect 82556 188961 82584 189051
rect 82541 188955 82599 188961
rect 82541 188921 82553 188955
rect 82587 188921 82599 188955
rect 82541 188915 82599 188921
rect 82081 188615 82139 188621
rect 82081 188581 82093 188615
rect 82127 188612 82139 188615
rect 82630 188612 82636 188624
rect 82127 188584 82636 188612
rect 82127 188581 82139 188584
rect 82081 188575 82139 188581
rect 82630 188572 82636 188584
rect 82688 188572 82694 188624
rect 78766 188368 78772 188420
rect 78824 188408 78830 188420
rect 82265 188411 82323 188417
rect 82265 188408 82277 188411
rect 78824 188380 82277 188408
rect 78824 188368 78830 188380
rect 82265 188377 82277 188380
rect 82311 188377 82323 188411
rect 82265 188371 82323 188377
rect 81621 187255 81679 187261
rect 81621 187221 81633 187255
rect 81667 187252 81679 187255
rect 82630 187252 82636 187264
rect 81667 187224 82636 187252
rect 81667 187221 81679 187224
rect 81621 187215 81679 187221
rect 82630 187212 82636 187224
rect 82688 187212 82694 187264
rect 82817 187119 82875 187125
rect 82817 187116 82829 187119
rect 82740 187088 82829 187116
rect 82357 186983 82415 186989
rect 82357 186949 82369 186983
rect 82403 186980 82415 186983
rect 82630 186980 82636 186992
rect 82403 186952 82636 186980
rect 82403 186949 82415 186952
rect 82357 186943 82415 186949
rect 82630 186940 82636 186952
rect 82688 186940 82694 186992
rect 82740 186844 82768 187088
rect 82817 187085 82829 187088
rect 82863 187085 82875 187119
rect 82817 187079 82875 187085
rect 82906 186980 82912 186992
rect 82867 186952 82912 186980
rect 82906 186940 82912 186952
rect 82964 186940 82970 186992
rect 503622 186980 503628 186992
rect 503583 186952 503628 186980
rect 503622 186940 503628 186952
rect 503680 186940 503686 186992
rect 82909 186847 82967 186853
rect 82909 186844 82921 186847
rect 82740 186816 82921 186844
rect 82909 186813 82921 186816
rect 82955 186813 82967 186847
rect 82909 186807 82967 186813
rect 82722 186668 82728 186720
rect 82780 186708 82786 186720
rect 82906 186708 82912 186720
rect 82780 186680 82912 186708
rect 82780 186668 82786 186680
rect 82906 186668 82912 186680
rect 82964 186668 82970 186720
rect 79594 185648 79600 185700
rect 79652 185688 79658 185700
rect 79962 185688 79968 185700
rect 79652 185660 79968 185688
rect 79652 185648 79658 185660
rect 79962 185648 79968 185660
rect 80020 185648 80026 185700
rect 82722 185688 82728 185700
rect 82683 185660 82728 185688
rect 82722 185648 82728 185660
rect 82780 185648 82786 185700
rect 14458 183472 14464 183524
rect 14516 183512 14522 183524
rect 78766 183512 78772 183524
rect 14516 183484 78772 183512
rect 14516 183472 14522 183484
rect 78766 183472 78772 183484
rect 78824 183472 78830 183524
rect 82630 182424 82636 182436
rect 82591 182396 82636 182424
rect 82630 182384 82636 182396
rect 82688 182384 82694 182436
rect 504818 182180 504824 182232
rect 504876 182220 504882 182232
rect 571978 182220 571984 182232
rect 504876 182192 571984 182220
rect 504876 182180 504882 182192
rect 571978 182180 571984 182192
rect 572036 182180 572042 182232
rect 524414 182112 524420 182164
rect 524472 182152 524478 182164
rect 524598 182152 524604 182164
rect 524472 182124 524604 182152
rect 524472 182112 524478 182124
rect 524598 182112 524604 182124
rect 524656 182112 524662 182164
rect 503070 181772 503076 181824
rect 503128 181812 503134 181824
rect 504818 181812 504824 181824
rect 503128 181784 504824 181812
rect 503128 181772 503134 181784
rect 504818 181772 504824 181784
rect 504876 181772 504882 181824
rect 514662 181092 514668 181144
rect 514720 181132 514726 181144
rect 521562 181132 521568 181144
rect 514720 181104 521568 181132
rect 514720 181092 514726 181104
rect 521562 181092 521568 181104
rect 521620 181092 521626 181144
rect 533982 180956 533988 181008
rect 534040 180996 534046 181008
rect 535454 180996 535460 181008
rect 534040 180968 535460 180996
rect 534040 180956 534046 180968
rect 535454 180956 535460 180968
rect 535512 180956 535518 181008
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 10502 180792 10508 180804
rect 3292 180764 10508 180792
rect 3292 180752 3298 180764
rect 10502 180752 10508 180764
rect 10560 180752 10566 180804
rect 503625 180183 503683 180189
rect 503625 180149 503637 180183
rect 503671 180180 503683 180183
rect 503806 180180 503812 180192
rect 503671 180152 503812 180180
rect 503671 180149 503683 180152
rect 503625 180143 503683 180149
rect 503806 180140 503812 180152
rect 503864 180140 503870 180192
rect 82630 178752 82636 178764
rect 82591 178724 82636 178752
rect 82630 178712 82636 178724
rect 82688 178712 82694 178764
rect 82541 178619 82599 178625
rect 82541 178585 82553 178619
rect 82587 178616 82599 178619
rect 82630 178616 82636 178628
rect 82587 178588 82636 178616
rect 82587 178585 82599 178588
rect 82541 178579 82599 178585
rect 82630 178576 82636 178588
rect 82688 178576 82694 178628
rect 501509 178211 501567 178217
rect 501509 178177 501521 178211
rect 501555 178208 501567 178211
rect 505830 178208 505836 178220
rect 501555 178180 505836 178208
rect 501555 178177 501567 178180
rect 501509 178171 501567 178177
rect 505830 178168 505836 178180
rect 505888 178168 505894 178220
rect 82817 177259 82875 177265
rect 82817 177225 82829 177259
rect 82863 177256 82875 177259
rect 82906 177256 82912 177268
rect 82863 177228 82912 177256
rect 82863 177225 82875 177228
rect 82817 177219 82875 177225
rect 82906 177216 82912 177228
rect 82964 177216 82970 177268
rect 82725 177123 82783 177129
rect 82725 177089 82737 177123
rect 82771 177120 82783 177123
rect 82906 177120 82912 177132
rect 82771 177092 82912 177120
rect 82771 177089 82783 177092
rect 82725 177083 82783 177089
rect 82906 177080 82912 177092
rect 82964 177080 82970 177132
rect 82906 176984 82912 176996
rect 82867 176956 82912 176984
rect 82906 176944 82912 176956
rect 82964 176944 82970 176996
rect 19978 176604 19984 176656
rect 20036 176644 20042 176656
rect 79962 176644 79968 176656
rect 20036 176616 79968 176644
rect 20036 176604 20042 176616
rect 79962 176604 79968 176616
rect 80020 176604 80026 176656
rect 82906 176644 82912 176656
rect 82867 176616 82912 176644
rect 82906 176604 82912 176616
rect 82964 176604 82970 176656
rect 79594 176576 79600 176588
rect 79555 176548 79600 176576
rect 79594 176536 79600 176548
rect 79652 176536 79658 176588
rect 79597 175559 79655 175565
rect 79597 175525 79609 175559
rect 79643 175556 79655 175559
rect 79962 175556 79968 175568
rect 79643 175528 79968 175556
rect 79643 175525 79655 175528
rect 79597 175519 79655 175525
rect 79962 175516 79968 175528
rect 80020 175516 80026 175568
rect 82725 173179 82783 173185
rect 82725 173145 82737 173179
rect 82771 173176 82783 173179
rect 82906 173176 82912 173188
rect 82771 173148 82912 173176
rect 82771 173145 82783 173148
rect 82725 173139 82783 173145
rect 82906 173136 82912 173148
rect 82964 173136 82970 173188
rect 503070 172932 503076 172984
rect 503128 172972 503134 172984
rect 505002 172972 505008 172984
rect 503128 172944 505008 172972
rect 503128 172932 503134 172944
rect 505002 172932 505008 172944
rect 505060 172932 505066 172984
rect 77386 171096 77392 171148
rect 77444 171136 77450 171148
rect 78674 171136 78680 171148
rect 77444 171108 78680 171136
rect 77444 171096 77450 171108
rect 78674 171096 78680 171108
rect 78732 171096 78738 171148
rect 510062 171028 510068 171080
rect 510120 171068 510126 171080
rect 580166 171068 580172 171080
rect 510120 171040 580172 171068
rect 510120 171028 510126 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 82630 170348 82636 170400
rect 82688 170388 82694 170400
rect 82688 170360 82768 170388
rect 82688 170348 82694 170360
rect 82630 170252 82636 170264
rect 82591 170224 82636 170252
rect 82630 170212 82636 170224
rect 82688 170212 82694 170264
rect 82630 170076 82636 170128
rect 82688 170116 82694 170128
rect 82740 170116 82768 170360
rect 82688 170088 82768 170116
rect 82688 170076 82694 170088
rect 505830 170008 505836 170060
rect 505888 170048 505894 170060
rect 506382 170048 506388 170060
rect 505888 170020 506388 170048
rect 505888 170008 505894 170020
rect 506382 170008 506388 170020
rect 506440 170008 506446 170060
rect 503622 169232 503628 169244
rect 503583 169204 503628 169232
rect 503622 169192 503628 169204
rect 503680 169192 503686 169244
rect 6822 168376 6828 168428
rect 6880 168416 6886 168428
rect 78674 168416 78680 168428
rect 6880 168388 78680 168416
rect 6880 168376 6886 168388
rect 78674 168376 78680 168388
rect 78732 168376 78738 168428
rect 82817 168419 82875 168425
rect 82817 168385 82829 168419
rect 82863 168416 82875 168419
rect 82998 168416 83004 168428
rect 82863 168388 83004 168416
rect 82863 168385 82875 168388
rect 82817 168379 82875 168385
rect 82998 168376 83004 168388
rect 83056 168376 83062 168428
rect 82725 167263 82783 167269
rect 82725 167229 82737 167263
rect 82771 167260 82783 167263
rect 82998 167260 83004 167272
rect 82771 167232 83004 167260
rect 82771 167229 82783 167232
rect 82725 167223 82783 167229
rect 82998 167220 83004 167232
rect 83056 167220 83062 167272
rect 82817 167127 82875 167133
rect 82817 167093 82829 167127
rect 82863 167124 82875 167127
rect 82998 167124 83004 167136
rect 82863 167096 83004 167124
rect 82863 167093 82875 167096
rect 82817 167087 82875 167093
rect 82998 167084 83004 167096
rect 83056 167084 83062 167136
rect 79594 167016 79600 167068
rect 79652 167056 79658 167068
rect 79962 167056 79968 167068
rect 79652 167028 79968 167056
rect 79652 167016 79658 167028
rect 79962 167016 79968 167028
rect 80020 167016 80026 167068
rect 82725 166719 82783 166725
rect 82725 166685 82737 166719
rect 82771 166716 82783 166719
rect 82998 166716 83004 166728
rect 82771 166688 83004 166716
rect 82771 166685 82783 166688
rect 82725 166679 82783 166685
rect 82998 166676 83004 166688
rect 83056 166676 83062 166728
rect 502978 166676 502984 166728
rect 503036 166716 503042 166728
rect 506382 166716 506388 166728
rect 503036 166688 506388 166716
rect 503036 166676 503042 166688
rect 506382 166676 506388 166688
rect 506440 166676 506446 166728
rect 501877 166379 501935 166385
rect 501877 166345 501889 166379
rect 501923 166376 501935 166379
rect 502978 166376 502984 166388
rect 501923 166348 502984 166376
rect 501923 166345 501935 166348
rect 501877 166339 501935 166345
rect 502978 166336 502984 166348
rect 503036 166336 503042 166388
rect 82909 166039 82967 166045
rect 82909 166005 82921 166039
rect 82955 166036 82967 166039
rect 82998 166036 83004 166048
rect 82955 166008 83004 166036
rect 82955 166005 82967 166008
rect 82909 165999 82967 166005
rect 82998 165996 83004 166008
rect 83056 165996 83062 166048
rect 501509 165631 501567 165637
rect 501509 165597 501521 165631
rect 501555 165628 501567 165631
rect 502978 165628 502984 165640
rect 501555 165600 502984 165628
rect 501555 165597 501567 165600
rect 501509 165591 501567 165597
rect 502978 165588 502984 165600
rect 503036 165588 503042 165640
rect 3418 165520 3424 165572
rect 3476 165560 3482 165572
rect 10410 165560 10416 165572
rect 3476 165532 10416 165560
rect 3476 165520 3482 165532
rect 10410 165520 10416 165532
rect 10468 165520 10474 165572
rect 503898 165520 503904 165572
rect 503956 165560 503962 165572
rect 527174 165560 527180 165572
rect 503956 165532 527180 165560
rect 503956 165520 503962 165532
rect 527174 165520 527180 165532
rect 527232 165520 527238 165572
rect 502978 164948 502984 164960
rect 502939 164920 502984 164948
rect 502978 164908 502984 164920
rect 503036 164908 503042 164960
rect 13722 164228 13728 164280
rect 13780 164268 13786 164280
rect 78674 164268 78680 164280
rect 13780 164240 78680 164268
rect 13780 164228 13786 164240
rect 78674 164228 78680 164240
rect 78732 164228 78738 164280
rect 501509 163795 501567 163801
rect 501509 163761 501521 163795
rect 501555 163792 501567 163795
rect 502978 163792 502984 163804
rect 501555 163764 502984 163792
rect 501555 163761 501567 163764
rect 501509 163755 501567 163761
rect 502978 163752 502984 163764
rect 503036 163752 503042 163804
rect 505830 162976 505836 162988
rect 505791 162948 505836 162976
rect 505830 162936 505836 162948
rect 505888 162936 505894 162988
rect 78766 162800 78772 162852
rect 78824 162840 78830 162852
rect 82633 162843 82691 162849
rect 82633 162840 82645 162843
rect 78824 162812 82645 162840
rect 78824 162800 78830 162812
rect 82633 162809 82645 162812
rect 82679 162809 82691 162843
rect 82633 162803 82691 162809
rect 502978 162800 502984 162852
rect 503036 162840 503042 162852
rect 503717 162843 503775 162849
rect 503717 162840 503729 162843
rect 503036 162812 503729 162840
rect 503036 162800 503042 162812
rect 503717 162809 503729 162812
rect 503763 162809 503775 162843
rect 524414 162840 524420 162852
rect 524375 162812 524420 162840
rect 503717 162803 503775 162809
rect 524414 162800 524420 162812
rect 524472 162800 524478 162852
rect 532694 162840 532700 162852
rect 532655 162812 532700 162840
rect 532694 162800 532700 162812
rect 532752 162800 532758 162852
rect 502889 162435 502947 162441
rect 502889 162401 502901 162435
rect 502935 162432 502947 162435
rect 502978 162432 502984 162444
rect 502935 162404 502984 162432
rect 502935 162401 502947 162404
rect 502889 162395 502947 162401
rect 502978 162392 502984 162404
rect 503036 162392 503042 162444
rect 81526 162120 81532 162172
rect 81584 162160 81590 162172
rect 81621 162163 81679 162169
rect 81621 162160 81633 162163
rect 81584 162132 81633 162160
rect 81584 162120 81590 162132
rect 81621 162129 81633 162132
rect 81667 162129 81679 162163
rect 81621 162123 81679 162129
rect 501969 162163 502027 162169
rect 501969 162129 501981 162163
rect 502015 162160 502027 162163
rect 502978 162160 502984 162172
rect 502015 162132 502984 162160
rect 502015 162129 502027 162132
rect 501969 162123 502027 162129
rect 502978 162120 502984 162132
rect 503036 162120 503042 162172
rect 503622 160692 503628 160744
rect 503680 160732 503686 160744
rect 503898 160732 503904 160744
rect 503680 160704 503904 160732
rect 503680 160692 503686 160704
rect 503898 160692 503904 160704
rect 503956 160692 503962 160744
rect 501690 159100 501696 159112
rect 501651 159072 501696 159100
rect 501690 159060 501696 159072
rect 501748 159060 501754 159112
rect 501874 158788 501880 158840
rect 501932 158828 501938 158840
rect 503622 158828 503628 158840
rect 501932 158800 503628 158828
rect 501932 158788 501938 158800
rect 503622 158788 503628 158800
rect 503680 158788 503686 158840
rect 501874 158652 501880 158704
rect 501932 158692 501938 158704
rect 502889 158695 502947 158701
rect 502889 158692 502901 158695
rect 501932 158664 502901 158692
rect 501932 158652 501938 158664
rect 502889 158661 502901 158664
rect 502935 158661 502947 158695
rect 502889 158655 502947 158661
rect 507762 158652 507768 158704
rect 507820 158692 507826 158704
rect 580166 158692 580172 158704
rect 507820 158664 580172 158692
rect 507820 158652 507826 158664
rect 580166 158652 580172 158664
rect 580224 158652 580230 158704
rect 82725 157607 82783 157613
rect 82725 157573 82737 157607
rect 82771 157604 82783 157607
rect 82906 157604 82912 157616
rect 82771 157576 82912 157604
rect 82771 157573 82783 157576
rect 82725 157567 82783 157573
rect 82906 157564 82912 157576
rect 82964 157564 82970 157616
rect 501598 157564 501604 157616
rect 501656 157604 501662 157616
rect 507486 157604 507492 157616
rect 501656 157576 507492 157604
rect 501656 157564 501662 157576
rect 507486 157564 507492 157576
rect 507544 157564 507550 157616
rect 82817 157539 82875 157545
rect 82817 157505 82829 157539
rect 82863 157536 82875 157539
rect 82998 157536 83004 157548
rect 82863 157508 83004 157536
rect 82863 157505 82875 157508
rect 82817 157499 82875 157505
rect 82998 157496 83004 157508
rect 83056 157496 83062 157548
rect 81526 157468 81532 157480
rect 81487 157440 81532 157468
rect 81526 157428 81532 157440
rect 81584 157428 81590 157480
rect 501509 157471 501567 157477
rect 501509 157437 501521 157471
rect 501555 157468 501567 157471
rect 501598 157468 501604 157480
rect 501555 157440 501604 157468
rect 501555 157437 501567 157440
rect 501509 157431 501567 157437
rect 501598 157428 501604 157440
rect 501656 157428 501662 157480
rect 78766 157292 78772 157344
rect 78824 157332 78830 157344
rect 79594 157332 79600 157344
rect 78824 157304 79600 157332
rect 78824 157292 78830 157304
rect 79594 157292 79600 157304
rect 79652 157292 79658 157344
rect 81526 157292 81532 157344
rect 81584 157332 81590 157344
rect 81621 157335 81679 157341
rect 81621 157332 81633 157335
rect 81584 157304 81633 157332
rect 81584 157292 81590 157304
rect 81621 157301 81633 157304
rect 81667 157301 81679 157335
rect 81621 157295 81679 157301
rect 81526 157196 81532 157208
rect 81487 157168 81532 157196
rect 81526 157156 81532 157168
rect 81584 157156 81590 157208
rect 82998 157060 83004 157072
rect 82832 157032 83004 157060
rect 82832 156856 82860 157032
rect 82998 157020 83004 157032
rect 83056 157020 83062 157072
rect 82906 156952 82912 157004
rect 82964 156992 82970 157004
rect 82964 156964 83044 156992
rect 82964 156952 82970 156964
rect 82906 156856 82912 156868
rect 82832 156828 82912 156856
rect 82906 156816 82912 156828
rect 82964 156816 82970 156868
rect 83016 156800 83044 156964
rect 82998 156748 83004 156800
rect 83056 156748 83062 156800
rect 82630 156340 82636 156392
rect 82688 156380 82694 156392
rect 82906 156380 82912 156392
rect 82688 156352 82912 156380
rect 82688 156340 82694 156352
rect 82906 156340 82912 156352
rect 82964 156340 82970 156392
rect 82630 156244 82636 156256
rect 82591 156216 82636 156244
rect 82630 156204 82636 156216
rect 82688 156204 82694 156256
rect 501874 155524 501880 155576
rect 501932 155564 501938 155576
rect 505557 155567 505615 155573
rect 505557 155564 505569 155567
rect 501932 155536 505569 155564
rect 501932 155524 501938 155536
rect 505557 155533 505569 155536
rect 505603 155533 505615 155567
rect 505557 155527 505615 155533
rect 501874 155388 501880 155440
rect 501932 155428 501938 155440
rect 502981 155431 503039 155437
rect 502981 155428 502993 155431
rect 501932 155400 502993 155428
rect 501932 155388 501938 155400
rect 502981 155397 502993 155400
rect 503027 155397 503039 155431
rect 502981 155391 503039 155397
rect 506290 155320 506296 155372
rect 506348 155360 506354 155372
rect 506348 155332 506428 155360
rect 506348 155320 506354 155332
rect 502334 155224 502340 155236
rect 501892 155196 502340 155224
rect 501892 155168 501920 155196
rect 502334 155184 502340 155196
rect 502392 155184 502398 155236
rect 506400 155168 506428 155332
rect 501874 155116 501880 155168
rect 501932 155116 501938 155168
rect 506382 155116 506388 155168
rect 506440 155116 506446 155168
rect 501693 155091 501751 155097
rect 501693 155057 501705 155091
rect 501739 155088 501751 155091
rect 502334 155088 502340 155100
rect 501739 155060 502340 155088
rect 501739 155057 501751 155060
rect 501693 155051 501751 155057
rect 502334 155048 502340 155060
rect 502392 155048 502398 155100
rect 501598 154844 501604 154896
rect 501656 154884 501662 154896
rect 501785 154887 501843 154893
rect 501785 154884 501797 154887
rect 501656 154856 501797 154884
rect 501656 154844 501662 154856
rect 501785 154853 501797 154856
rect 501831 154853 501843 154887
rect 501785 154847 501843 154853
rect 501690 154708 501696 154760
rect 501748 154748 501754 154760
rect 501969 154751 502027 154757
rect 501969 154748 501981 154751
rect 501748 154720 501981 154748
rect 501748 154708 501754 154720
rect 501969 154717 501981 154720
rect 502015 154717 502027 154751
rect 501969 154711 502027 154717
rect 501690 154572 501696 154624
rect 501748 154612 501754 154624
rect 503625 154615 503683 154621
rect 503625 154612 503637 154615
rect 501748 154584 503637 154612
rect 501748 154572 501754 154584
rect 503625 154581 503637 154584
rect 503671 154581 503683 154615
rect 503625 154575 503683 154581
rect 524414 153252 524420 153264
rect 524375 153224 524420 153252
rect 524414 153212 524420 153224
rect 524472 153212 524478 153264
rect 532694 153252 532700 153264
rect 532655 153224 532700 153252
rect 532694 153212 532700 153224
rect 532752 153212 532758 153264
rect 504545 152575 504603 152581
rect 504545 152541 504557 152575
rect 504591 152572 504603 152575
rect 505830 152572 505836 152584
rect 504591 152544 505836 152572
rect 504591 152541 504603 152544
rect 504545 152535 504603 152541
rect 505830 152532 505836 152544
rect 505888 152532 505894 152584
rect 82906 152504 82912 152516
rect 82867 152476 82912 152504
rect 82906 152464 82912 152476
rect 82964 152464 82970 152516
rect 82817 152371 82875 152377
rect 82817 152337 82829 152371
rect 82863 152368 82875 152371
rect 82906 152368 82912 152380
rect 82863 152340 82912 152368
rect 82863 152337 82875 152340
rect 82817 152331 82875 152337
rect 82906 152328 82912 152340
rect 82964 152328 82970 152380
rect 82725 152167 82783 152173
rect 82725 152133 82737 152167
rect 82771 152164 82783 152167
rect 82906 152164 82912 152176
rect 82771 152136 82912 152164
rect 82771 152133 82783 152136
rect 82725 152127 82783 152133
rect 82906 152124 82912 152136
rect 82964 152124 82970 152176
rect 505741 152099 505799 152105
rect 505741 152065 505753 152099
rect 505787 152096 505799 152099
rect 505830 152096 505836 152108
rect 505787 152068 505836 152096
rect 505787 152065 505799 152068
rect 505741 152059 505799 152065
rect 505830 152056 505836 152068
rect 505888 152056 505894 152108
rect 501506 151920 501512 151972
rect 501564 151960 501570 151972
rect 501564 151932 501644 151960
rect 501564 151920 501570 151932
rect 501506 151824 501512 151836
rect 501467 151796 501512 151824
rect 501506 151784 501512 151796
rect 501564 151784 501570 151836
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 10318 151756 10324 151768
rect 3200 151728 10324 151756
rect 3200 151716 3206 151728
rect 10318 151716 10324 151728
rect 10376 151716 10382 151768
rect 501506 151648 501512 151700
rect 501564 151688 501570 151700
rect 501616 151688 501644 151932
rect 505557 151895 505615 151901
rect 505557 151861 505569 151895
rect 505603 151892 505615 151895
rect 505830 151892 505836 151904
rect 505603 151864 505836 151892
rect 505603 151861 505615 151864
rect 505557 151855 505615 151861
rect 505830 151852 505836 151864
rect 505888 151852 505894 151904
rect 501564 151660 501644 151688
rect 501564 151648 501570 151660
rect 505830 151280 505836 151292
rect 505791 151252 505836 151280
rect 505830 151240 505836 151252
rect 505888 151240 505894 151292
rect 78766 151008 78772 151020
rect 78727 150980 78772 151008
rect 78766 150968 78772 150980
rect 78824 150968 78830 151020
rect 56502 150424 56508 150476
rect 56560 150464 56566 150476
rect 78766 150464 78772 150476
rect 56560 150436 78772 150464
rect 56560 150424 56566 150436
rect 78766 150424 78772 150436
rect 78824 150424 78830 150476
rect 78766 150328 78772 150340
rect 78727 150300 78772 150328
rect 78766 150288 78772 150300
rect 78824 150288 78830 150340
rect 501693 149039 501751 149045
rect 501693 149005 501705 149039
rect 501739 149036 501751 149039
rect 504542 149036 504548 149048
rect 501739 149008 504548 149036
rect 501739 149005 501751 149008
rect 501693 148999 501751 149005
rect 504542 148996 504548 149008
rect 504600 148996 504606 149048
rect 502334 148928 502340 148980
rect 502392 148928 502398 148980
rect 502352 148900 502380 148928
rect 506385 148903 506443 148909
rect 506385 148900 506397 148903
rect 502352 148872 506397 148900
rect 506385 148869 506397 148872
rect 506431 148869 506443 148903
rect 506385 148863 506443 148869
rect 502245 148835 502303 148841
rect 502245 148801 502257 148835
rect 502291 148832 502303 148835
rect 502334 148832 502340 148844
rect 502291 148804 502340 148832
rect 502291 148801 502303 148804
rect 502245 148795 502303 148801
rect 502334 148792 502340 148804
rect 502392 148792 502398 148844
rect 504358 148724 504364 148776
rect 504416 148764 504422 148776
rect 504542 148764 504548 148776
rect 504416 148736 504548 148764
rect 504416 148724 504422 148736
rect 504542 148724 504548 148736
rect 504600 148724 504606 148776
rect 504082 148588 504088 148640
rect 504140 148628 504146 148640
rect 504358 148628 504364 148640
rect 504140 148600 504364 148628
rect 504140 148588 504146 148600
rect 504358 148588 504364 148600
rect 504416 148588 504422 148640
rect 503714 148016 503720 148028
rect 503675 147988 503720 148016
rect 503714 147976 503720 147988
rect 503772 147976 503778 148028
rect 78766 147636 78772 147688
rect 78824 147676 78830 147688
rect 79594 147676 79600 147688
rect 78824 147648 79600 147676
rect 78824 147636 78830 147648
rect 79594 147636 79600 147648
rect 79652 147636 79658 147688
rect 503714 147636 503720 147688
rect 503772 147676 503778 147688
rect 563054 147676 563060 147688
rect 503772 147648 563060 147676
rect 503772 147636 503778 147648
rect 563054 147636 563060 147648
rect 563112 147636 563118 147688
rect 502334 147472 502340 147484
rect 502295 147444 502340 147472
rect 502334 147432 502340 147444
rect 502392 147432 502398 147484
rect 504542 147364 504548 147416
rect 504600 147404 504606 147416
rect 505741 147407 505799 147413
rect 505741 147404 505753 147407
rect 504600 147376 505753 147404
rect 504600 147364 504606 147376
rect 505741 147373 505753 147376
rect 505787 147373 505799 147407
rect 505741 147367 505799 147373
rect 501509 147271 501567 147277
rect 501509 147237 501521 147271
rect 501555 147268 501567 147271
rect 502334 147268 502340 147280
rect 501555 147240 502340 147268
rect 501555 147237 501567 147240
rect 501509 147231 501567 147237
rect 502334 147228 502340 147240
rect 502392 147228 502398 147280
rect 503714 146996 503720 147008
rect 503675 146968 503720 146996
rect 503714 146956 503720 146968
rect 503772 146956 503778 147008
rect 504082 146140 504088 146192
rect 504140 146180 504146 146192
rect 504545 146183 504603 146189
rect 504545 146180 504557 146183
rect 504140 146152 504557 146180
rect 504140 146140 504146 146152
rect 504545 146149 504557 146152
rect 504591 146149 504603 146183
rect 504545 146143 504603 146149
rect 504082 145976 504088 145988
rect 504043 145948 504088 145976
rect 504082 145936 504088 145948
rect 504140 145936 504146 145988
rect 82817 145911 82875 145917
rect 82817 145877 82829 145911
rect 82863 145908 82875 145911
rect 82906 145908 82912 145920
rect 82863 145880 82912 145908
rect 82863 145877 82875 145880
rect 82817 145871 82875 145877
rect 82906 145868 82912 145880
rect 82964 145868 82970 145920
rect 82906 145772 82912 145784
rect 82867 145744 82912 145772
rect 82906 145732 82912 145744
rect 82964 145732 82970 145784
rect 82817 145503 82875 145509
rect 82817 145469 82829 145503
rect 82863 145500 82875 145503
rect 82906 145500 82912 145512
rect 82863 145472 82912 145500
rect 82863 145469 82875 145472
rect 82817 145463 82875 145469
rect 82906 145460 82912 145472
rect 82964 145460 82970 145512
rect 501509 144483 501567 144489
rect 501509 144449 501521 144483
rect 501555 144480 501567 144483
rect 504082 144480 504088 144492
rect 501555 144452 504088 144480
rect 501555 144449 501567 144452
rect 501509 144443 501567 144449
rect 504082 144440 504088 144452
rect 504140 144440 504146 144492
rect 80238 144032 80244 144084
rect 80296 144072 80302 144084
rect 80425 144075 80483 144081
rect 80425 144072 80437 144075
rect 80296 144044 80437 144072
rect 80296 144032 80302 144044
rect 80425 144041 80437 144044
rect 80471 144041 80483 144075
rect 80425 144035 80483 144041
rect 501877 143667 501935 143673
rect 501877 143633 501889 143667
rect 501923 143664 501935 143667
rect 504542 143664 504548 143676
rect 501923 143636 504548 143664
rect 501923 143633 501935 143636
rect 501877 143627 501935 143633
rect 504542 143624 504548 143636
rect 504600 143624 504606 143676
rect 505830 143664 505836 143676
rect 505791 143636 505836 143664
rect 505830 143624 505836 143636
rect 505888 143624 505894 143676
rect 524414 143528 524420 143540
rect 524375 143500 524420 143528
rect 524414 143488 524420 143500
rect 524472 143488 524478 143540
rect 532694 143528 532700 143540
rect 532655 143500 532700 143528
rect 532694 143488 532700 143500
rect 532752 143488 532758 143540
rect 503625 143395 503683 143401
rect 503625 143361 503637 143395
rect 503671 143392 503683 143395
rect 504542 143392 504548 143404
rect 503671 143364 504548 143392
rect 503671 143361 503683 143364
rect 503625 143355 503683 143361
rect 504542 143352 504548 143364
rect 504600 143352 504606 143404
rect 501877 141831 501935 141837
rect 501877 141797 501889 141831
rect 501923 141828 501935 141831
rect 502150 141828 502156 141840
rect 501923 141800 502156 141828
rect 501923 141797 501935 141800
rect 501877 141791 501935 141797
rect 502150 141788 502156 141800
rect 502208 141788 502214 141840
rect 501874 141652 501880 141704
rect 501932 141692 501938 141704
rect 502150 141692 502156 141704
rect 501932 141664 502156 141692
rect 501932 141652 501938 141664
rect 502150 141652 502156 141664
rect 502208 141652 502214 141704
rect 506290 140632 506296 140684
rect 506348 140672 506354 140684
rect 507762 140672 507768 140684
rect 506348 140644 507768 140672
rect 506348 140632 506354 140644
rect 507762 140632 507768 140644
rect 507820 140632 507826 140684
rect 501874 140496 501880 140548
rect 501932 140536 501938 140548
rect 502521 140539 502579 140545
rect 502521 140536 502533 140539
rect 501932 140508 502533 140536
rect 501932 140496 501938 140508
rect 502521 140505 502533 140508
rect 502567 140505 502579 140539
rect 502521 140499 502579 140505
rect 80146 140400 80152 140412
rect 80107 140372 80152 140400
rect 80146 140360 80152 140372
rect 80204 140360 80210 140412
rect 501874 140360 501880 140412
rect 501932 140400 501938 140412
rect 502153 140403 502211 140409
rect 502153 140400 502165 140403
rect 501932 140372 502165 140400
rect 501932 140360 501938 140372
rect 502153 140369 502165 140372
rect 502199 140369 502211 140403
rect 502153 140363 502211 140369
rect 501874 140224 501880 140276
rect 501932 140264 501938 140276
rect 502429 140267 502487 140273
rect 502429 140264 502441 140267
rect 501932 140236 502441 140264
rect 501932 140224 501938 140236
rect 502429 140233 502441 140236
rect 502475 140233 502487 140267
rect 502429 140227 502487 140233
rect 501785 140131 501843 140137
rect 501785 140097 501797 140131
rect 501831 140128 501843 140131
rect 501874 140128 501880 140140
rect 501831 140100 501880 140128
rect 501831 140097 501843 140100
rect 501785 140091 501843 140097
rect 501874 140088 501880 140100
rect 501932 140088 501938 140140
rect 501874 139952 501880 140004
rect 501932 139992 501938 140004
rect 501969 139995 502027 140001
rect 501969 139992 501981 139995
rect 501932 139964 501981 139992
rect 501932 139952 501938 139964
rect 501969 139961 501981 139964
rect 502015 139961 502027 139995
rect 501969 139955 502027 139961
rect 82906 138700 82912 138712
rect 82867 138672 82912 138700
rect 82906 138660 82912 138672
rect 82964 138660 82970 138712
rect 82817 138499 82875 138505
rect 82817 138465 82829 138499
rect 82863 138496 82875 138499
rect 82906 138496 82912 138508
rect 82863 138468 82912 138496
rect 82863 138465 82875 138468
rect 82817 138459 82875 138465
rect 82906 138456 82912 138468
rect 82964 138456 82970 138508
rect 502334 138252 502340 138304
rect 502392 138292 502398 138304
rect 504085 138295 504143 138301
rect 504085 138292 504097 138295
rect 502392 138264 504097 138292
rect 502392 138252 502398 138264
rect 504085 138261 504097 138264
rect 504131 138261 504143 138295
rect 504085 138255 504143 138261
rect 501601 138091 501659 138097
rect 501601 138057 501613 138091
rect 501647 138088 501659 138091
rect 501874 138088 501880 138100
rect 501647 138060 501880 138088
rect 501647 138057 501659 138060
rect 501601 138051 501659 138057
rect 501874 138048 501880 138060
rect 501932 138048 501938 138100
rect 501874 137776 501880 137828
rect 501932 137816 501938 137828
rect 502061 137819 502119 137825
rect 502061 137816 502073 137819
rect 501932 137788 502073 137816
rect 501932 137776 501938 137788
rect 502061 137785 502073 137788
rect 502107 137785 502119 137819
rect 502061 137779 502119 137785
rect 501969 137479 502027 137485
rect 501969 137445 501981 137479
rect 502015 137476 502027 137479
rect 502334 137476 502340 137488
rect 502015 137448 502340 137476
rect 502015 137445 502027 137448
rect 501969 137439 502027 137445
rect 502334 137436 502340 137448
rect 502392 137436 502398 137488
rect 82725 137343 82783 137349
rect 82725 137309 82737 137343
rect 82771 137340 82783 137343
rect 82906 137340 82912 137352
rect 82771 137312 82912 137340
rect 82771 137309 82783 137312
rect 82725 137303 82783 137309
rect 82906 137300 82912 137312
rect 82964 137300 82970 137352
rect 80422 137204 80428 137216
rect 80383 137176 80428 137204
rect 80422 137164 80428 137176
rect 80480 137164 80486 137216
rect 82633 137207 82691 137213
rect 82633 137173 82645 137207
rect 82679 137204 82691 137207
rect 82906 137204 82912 137216
rect 82679 137176 82912 137204
rect 82679 137173 82691 137176
rect 82633 137167 82691 137173
rect 82906 137164 82912 137176
rect 82964 137164 82970 137216
rect 80149 137071 80207 137077
rect 80149 137037 80161 137071
rect 80195 137068 80207 137071
rect 80422 137068 80428 137080
rect 80195 137040 80428 137068
rect 80195 137037 80207 137040
rect 80149 137031 80207 137037
rect 80422 137028 80428 137040
rect 80480 137028 80486 137080
rect 82906 137068 82912 137080
rect 82867 137040 82912 137068
rect 82906 137028 82912 137040
rect 82964 137028 82970 137080
rect 501874 137028 501880 137080
rect 501932 137068 501938 137080
rect 502153 137071 502211 137077
rect 502153 137068 502165 137071
rect 501932 137040 502165 137068
rect 501932 137028 501938 137040
rect 502153 137037 502165 137040
rect 502199 137037 502211 137071
rect 502153 137031 502211 137037
rect 82725 136935 82783 136941
rect 82725 136901 82737 136935
rect 82771 136932 82783 136935
rect 82906 136932 82912 136944
rect 82771 136904 82912 136932
rect 82771 136901 82783 136904
rect 82725 136895 82783 136901
rect 82906 136892 82912 136904
rect 82964 136892 82970 136944
rect 501874 136892 501880 136944
rect 501932 136932 501938 136944
rect 502429 136935 502487 136941
rect 502429 136932 502441 136935
rect 501932 136904 502441 136932
rect 501932 136892 501938 136904
rect 502429 136901 502441 136904
rect 502475 136901 502487 136935
rect 502429 136895 502487 136901
rect 80974 136864 80980 136876
rect 80935 136836 80980 136864
rect 80974 136824 80980 136836
rect 81032 136824 81038 136876
rect 80974 136620 80980 136672
rect 81032 136660 81038 136672
rect 82906 136660 82912 136672
rect 81032 136632 82912 136660
rect 81032 136620 81038 136632
rect 82906 136620 82912 136632
rect 82964 136620 82970 136672
rect 80974 136524 80980 136536
rect 80935 136496 80980 136524
rect 80974 136484 80980 136496
rect 81032 136484 81038 136536
rect 502337 136323 502395 136329
rect 502337 136289 502349 136323
rect 502383 136320 502395 136323
rect 503714 136320 503720 136332
rect 502383 136292 503720 136320
rect 502383 136289 502395 136292
rect 502337 136283 502395 136289
rect 503714 136280 503720 136292
rect 503772 136280 503778 136332
rect 501601 136187 501659 136193
rect 501601 136153 501613 136187
rect 501647 136184 501659 136187
rect 501690 136184 501696 136196
rect 501647 136156 501696 136184
rect 501647 136153 501659 136156
rect 501601 136147 501659 136153
rect 501690 136144 501696 136156
rect 501748 136144 501754 136196
rect 78766 135668 78772 135720
rect 78824 135708 78830 135720
rect 79594 135708 79600 135720
rect 78824 135680 79600 135708
rect 78824 135668 78830 135680
rect 79594 135668 79600 135680
rect 79652 135668 79658 135720
rect 501874 135504 501880 135516
rect 501835 135476 501880 135504
rect 501874 135464 501880 135476
rect 501932 135464 501938 135516
rect 503714 133940 503720 133952
rect 503675 133912 503720 133940
rect 503714 133900 503720 133912
rect 503772 133900 503778 133952
rect 524414 133940 524420 133952
rect 524375 133912 524420 133940
rect 524414 133900 524420 133912
rect 524472 133900 524478 133952
rect 532694 133940 532700 133952
rect 532655 133912 532700 133940
rect 532694 133900 532700 133912
rect 532752 133900 532758 133952
rect 78766 133288 78772 133340
rect 78824 133328 78830 133340
rect 79597 133331 79655 133337
rect 79597 133328 79609 133331
rect 78824 133300 79609 133328
rect 78824 133288 78830 133300
rect 79597 133297 79609 133300
rect 79643 133297 79655 133331
rect 79597 133291 79655 133297
rect 501601 133331 501659 133337
rect 501601 133297 501613 133331
rect 501647 133328 501659 133331
rect 501690 133328 501696 133340
rect 501647 133300 501696 133328
rect 501647 133297 501659 133300
rect 501601 133291 501659 133297
rect 501690 133288 501696 133300
rect 501748 133288 501754 133340
rect 82909 133195 82967 133201
rect 82909 133161 82921 133195
rect 82955 133192 82967 133195
rect 82998 133192 83004 133204
rect 82955 133164 83004 133192
rect 82955 133161 82967 133164
rect 82909 133155 82967 133161
rect 82998 133152 83004 133164
rect 83056 133152 83062 133204
rect 501690 133192 501696 133204
rect 501651 133164 501696 133192
rect 501690 133152 501696 133164
rect 501748 133152 501754 133204
rect 82817 133059 82875 133065
rect 82817 133025 82829 133059
rect 82863 133056 82875 133059
rect 82906 133056 82912 133068
rect 82863 133028 82912 133056
rect 82863 133025 82875 133028
rect 82817 133019 82875 133025
rect 82906 133016 82912 133028
rect 82964 133016 82970 133068
rect 501693 133059 501751 133065
rect 501693 133025 501705 133059
rect 501739 133056 501751 133059
rect 502245 133059 502303 133065
rect 502245 133056 502257 133059
rect 501739 133028 502257 133056
rect 501739 133025 501751 133028
rect 501693 133019 501751 133025
rect 502245 133025 502257 133028
rect 502291 133025 502303 133059
rect 502245 133019 502303 133025
rect 501969 132515 502027 132521
rect 501969 132481 501981 132515
rect 502015 132512 502027 132515
rect 503622 132512 503628 132524
rect 502015 132484 503628 132512
rect 502015 132481 502027 132484
rect 501969 132475 502027 132481
rect 503622 132472 503628 132484
rect 503680 132472 503686 132524
rect 82633 132311 82691 132317
rect 82633 132277 82645 132311
rect 82679 132308 82691 132311
rect 82906 132308 82912 132320
rect 82679 132280 82912 132308
rect 82679 132277 82691 132280
rect 82633 132271 82691 132277
rect 82906 132268 82912 132280
rect 82964 132268 82970 132320
rect 505830 131832 505836 131844
rect 505791 131804 505836 131832
rect 505830 131792 505836 131804
rect 505888 131792 505894 131844
rect 506382 131832 506388 131844
rect 506343 131804 506388 131832
rect 506382 131792 506388 131804
rect 506440 131792 506446 131844
rect 501509 131087 501567 131093
rect 501509 131053 501521 131087
rect 501555 131084 501567 131087
rect 503441 131087 503499 131093
rect 503441 131084 503453 131087
rect 501555 131056 503453 131084
rect 501555 131053 501567 131056
rect 501509 131047 501567 131053
rect 503441 131053 503453 131056
rect 503487 131053 503499 131087
rect 503714 131084 503720 131096
rect 503675 131056 503720 131084
rect 503441 131047 503499 131053
rect 503714 131044 503720 131056
rect 503772 131044 503778 131096
rect 502337 130611 502395 130617
rect 502337 130577 502349 130611
rect 502383 130608 502395 130611
rect 503714 130608 503720 130620
rect 502383 130580 503720 130608
rect 502383 130577 502395 130580
rect 502337 130571 502395 130577
rect 503714 130568 503720 130580
rect 503772 130568 503778 130620
rect 502521 129999 502579 130005
rect 502521 129965 502533 129999
rect 502567 129996 502579 129999
rect 503714 129996 503720 130008
rect 502567 129968 503720 129996
rect 502567 129965 502579 129968
rect 502521 129959 502579 129965
rect 503714 129956 503720 129968
rect 503772 129956 503778 130008
rect 82630 129072 82636 129124
rect 82688 129072 82694 129124
rect 82648 128908 82676 129072
rect 82722 128908 82728 128920
rect 82648 128880 82728 128908
rect 82722 128868 82728 128880
rect 82780 128868 82786 128920
rect 79870 127848 79876 127900
rect 79928 127888 79934 127900
rect 80422 127888 80428 127900
rect 79928 127860 80428 127888
rect 79928 127848 79934 127860
rect 80422 127848 80428 127860
rect 80480 127848 80486 127900
rect 503533 127823 503591 127829
rect 503533 127789 503545 127823
rect 503579 127820 503591 127823
rect 503622 127820 503628 127832
rect 503579 127792 503628 127820
rect 503579 127789 503591 127792
rect 503533 127783 503591 127789
rect 503622 127780 503628 127792
rect 503680 127780 503686 127832
rect 503622 127684 503628 127696
rect 503583 127656 503628 127684
rect 503622 127644 503628 127656
rect 503680 127644 503686 127696
rect 501598 127344 501604 127356
rect 501559 127316 501604 127344
rect 501598 127304 501604 127316
rect 501656 127304 501662 127356
rect 501874 127344 501880 127356
rect 501835 127316 501880 127344
rect 501874 127304 501880 127316
rect 501932 127304 501938 127356
rect 502150 127344 502156 127356
rect 502111 127316 502156 127344
rect 502150 127304 502156 127316
rect 502208 127304 502214 127356
rect 501785 127211 501843 127217
rect 501785 127177 501797 127211
rect 501831 127208 501843 127211
rect 501874 127208 501880 127220
rect 501831 127180 501880 127208
rect 501831 127177 501843 127180
rect 501785 127171 501843 127177
rect 501874 127168 501880 127180
rect 501932 127168 501938 127220
rect 501509 127143 501567 127149
rect 501509 127109 501521 127143
rect 501555 127140 501567 127143
rect 502150 127140 502156 127152
rect 501555 127112 502156 127140
rect 501555 127109 501567 127112
rect 501509 127103 501567 127109
rect 502150 127100 502156 127112
rect 502208 127100 502214 127152
rect 505830 126420 505836 126472
rect 505888 126460 505894 126472
rect 506290 126460 506296 126472
rect 505888 126432 506296 126460
rect 505888 126420 505894 126432
rect 506290 126420 506296 126432
rect 506348 126420 506354 126472
rect 82354 125536 82360 125588
rect 82412 125576 82418 125588
rect 82412 125548 82492 125576
rect 82412 125536 82418 125548
rect 82464 125384 82492 125548
rect 82446 125332 82452 125384
rect 82504 125332 82510 125384
rect 503533 124831 503591 124837
rect 503533 124797 503545 124831
rect 503579 124828 503591 124831
rect 503622 124828 503628 124840
rect 503579 124800 503628 124828
rect 503579 124797 503591 124800
rect 503533 124791 503591 124797
rect 503622 124788 503628 124800
rect 503680 124788 503686 124840
rect 501506 124760 501512 124772
rect 501467 124732 501512 124760
rect 501506 124720 501512 124732
rect 501564 124720 501570 124772
rect 502610 124760 502616 124772
rect 502571 124732 502616 124760
rect 502610 124720 502616 124732
rect 502668 124720 502674 124772
rect 501506 124584 501512 124636
rect 501564 124624 501570 124636
rect 501782 124624 501788 124636
rect 501564 124596 501788 124624
rect 501564 124584 501570 124596
rect 501782 124584 501788 124596
rect 501840 124584 501846 124636
rect 507394 124108 507400 124160
rect 507452 124148 507458 124160
rect 580166 124148 580172 124160
rect 507452 124120 580172 124148
rect 507452 124108 507458 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 524414 124080 524420 124092
rect 524375 124052 524420 124080
rect 524414 124040 524420 124052
rect 524472 124040 524478 124092
rect 532694 124080 532700 124092
rect 532655 124052 532700 124080
rect 532694 124040 532700 124052
rect 532752 124040 532758 124092
rect 501782 123836 501788 123888
rect 501840 123876 501846 123888
rect 501969 123879 502027 123885
rect 501969 123876 501981 123879
rect 501840 123848 501981 123876
rect 501840 123836 501846 123848
rect 501969 123845 501981 123848
rect 502015 123845 502027 123879
rect 501969 123839 502027 123845
rect 502150 123740 502156 123752
rect 502111 123712 502156 123740
rect 502150 123700 502156 123712
rect 502208 123700 502214 123752
rect 82078 123672 82084 123684
rect 82039 123644 82084 123672
rect 82078 123632 82084 123644
rect 82136 123632 82142 123684
rect 82817 123675 82875 123681
rect 82817 123641 82829 123675
rect 82863 123672 82875 123675
rect 82906 123672 82912 123684
rect 82863 123644 82912 123672
rect 82863 123641 82875 123644
rect 82817 123635 82875 123641
rect 82906 123632 82912 123644
rect 82964 123632 82970 123684
rect 82446 123604 82452 123616
rect 82407 123576 82452 123604
rect 82446 123564 82452 123576
rect 82504 123564 82510 123616
rect 81986 123496 81992 123548
rect 82044 123536 82050 123548
rect 82044 123508 82492 123536
rect 82044 123496 82050 123508
rect 80425 123471 80483 123477
rect 80425 123437 80437 123471
rect 80471 123468 80483 123471
rect 82078 123468 82084 123480
rect 80471 123440 82084 123468
rect 80471 123437 80483 123440
rect 80425 123431 80483 123437
rect 82078 123428 82084 123440
rect 82136 123428 82142 123480
rect 81986 123360 81992 123412
rect 82044 123400 82050 123412
rect 82262 123400 82268 123412
rect 82044 123372 82268 123400
rect 82044 123360 82050 123372
rect 82262 123360 82268 123372
rect 82320 123360 82326 123412
rect 82464 123208 82492 123508
rect 501598 123428 501604 123480
rect 501656 123468 501662 123480
rect 501693 123471 501751 123477
rect 501693 123468 501705 123471
rect 501656 123440 501705 123468
rect 501656 123428 501662 123440
rect 501693 123437 501705 123440
rect 501739 123437 501751 123471
rect 501693 123431 501751 123437
rect 501598 123332 501604 123344
rect 501559 123304 501604 123332
rect 501598 123292 501604 123304
rect 501656 123292 501662 123344
rect 82446 123156 82452 123208
rect 82504 123156 82510 123208
rect 501601 123199 501659 123205
rect 501601 123165 501613 123199
rect 501647 123196 501659 123199
rect 502337 123199 502395 123205
rect 502337 123196 502349 123199
rect 501647 123168 502349 123196
rect 501647 123165 501659 123168
rect 501601 123159 501659 123165
rect 502337 123165 502349 123168
rect 502383 123165 502395 123199
rect 502337 123159 502395 123165
rect 82170 123088 82176 123140
rect 82228 123128 82234 123140
rect 82538 123128 82544 123140
rect 82228 123100 82544 123128
rect 82228 123088 82234 123100
rect 82538 123088 82544 123100
rect 82596 123088 82602 123140
rect 76926 122748 76932 122800
rect 76984 122788 76990 122800
rect 103517 122791 103575 122797
rect 103517 122788 103529 122791
rect 76984 122760 103529 122788
rect 76984 122748 76990 122760
rect 103517 122757 103529 122760
rect 103563 122757 103575 122791
rect 103517 122751 103575 122757
rect 326985 122791 327043 122797
rect 326985 122757 326997 122791
rect 327031 122788 327043 122791
rect 510154 122788 510160 122800
rect 327031 122760 510160 122788
rect 327031 122757 327043 122760
rect 326985 122751 327043 122757
rect 510154 122748 510160 122760
rect 510212 122748 510218 122800
rect 80425 122723 80483 122729
rect 80425 122689 80437 122723
rect 80471 122720 80483 122723
rect 81897 122723 81955 122729
rect 81897 122720 81909 122723
rect 80471 122692 81909 122720
rect 80471 122689 80483 122692
rect 80425 122683 80483 122689
rect 81897 122689 81909 122692
rect 81943 122689 81955 122723
rect 81897 122683 81955 122689
rect 83458 122680 83464 122732
rect 83516 122720 83522 122732
rect 120534 122720 120540 122732
rect 83516 122692 120540 122720
rect 83516 122680 83522 122692
rect 120534 122680 120540 122692
rect 120592 122680 120598 122732
rect 124306 122680 124312 122732
rect 124364 122720 124370 122732
rect 133782 122720 133788 122732
rect 124364 122692 133788 122720
rect 124364 122680 124370 122692
rect 133782 122680 133788 122692
rect 133840 122680 133846 122732
rect 286962 122680 286968 122732
rect 287020 122720 287026 122732
rect 504358 122720 504364 122732
rect 287020 122692 504364 122720
rect 287020 122680 287026 122692
rect 504358 122680 504364 122692
rect 504416 122680 504422 122732
rect 81158 122612 81164 122664
rect 81216 122652 81222 122664
rect 128354 122652 128360 122664
rect 81216 122624 128360 122652
rect 81216 122612 81222 122624
rect 128354 122612 128360 122624
rect 128412 122612 128418 122664
rect 143626 122612 143632 122664
rect 143684 122652 143690 122664
rect 153102 122652 153108 122664
rect 143684 122624 153108 122652
rect 143684 122612 143690 122624
rect 153102 122612 153108 122624
rect 153160 122612 153166 122664
rect 249886 122612 249892 122664
rect 249944 122652 249950 122664
rect 259362 122652 259368 122664
rect 249944 122624 259368 122652
rect 249944 122612 249950 122624
rect 259362 122612 259368 122624
rect 259420 122612 259426 122664
rect 284202 122612 284208 122664
rect 284260 122652 284266 122664
rect 507026 122652 507032 122664
rect 284260 122624 507032 122652
rect 284260 122612 284266 122624
rect 507026 122612 507032 122624
rect 507084 122612 507090 122664
rect 81342 122544 81348 122596
rect 81400 122584 81406 122596
rect 156049 122587 156107 122593
rect 156049 122584 156061 122587
rect 81400 122556 156061 122584
rect 81400 122544 81406 122556
rect 156049 122553 156061 122556
rect 156095 122553 156107 122587
rect 156049 122547 156107 122553
rect 253842 122544 253848 122596
rect 253900 122584 253906 122596
rect 503806 122584 503812 122596
rect 253900 122556 503812 122584
rect 253900 122544 253906 122556
rect 503806 122544 503812 122556
rect 503864 122544 503870 122596
rect 82354 122476 82360 122528
rect 82412 122516 82418 122528
rect 338117 122519 338175 122525
rect 338117 122516 338129 122519
rect 82412 122488 338129 122516
rect 82412 122476 82418 122488
rect 338117 122485 338129 122488
rect 338163 122485 338175 122519
rect 338117 122479 338175 122485
rect 365622 122476 365628 122528
rect 365680 122516 365686 122528
rect 505278 122516 505284 122528
rect 365680 122488 505284 122516
rect 365680 122476 365686 122488
rect 505278 122476 505284 122488
rect 505336 122476 505342 122528
rect 83550 122408 83556 122460
rect 83608 122448 83614 122460
rect 166994 122448 167000 122460
rect 83608 122420 167000 122448
rect 83608 122408 83614 122420
rect 166994 122408 167000 122420
rect 167052 122408 167058 122460
rect 172606 122408 172612 122460
rect 172664 122448 172670 122460
rect 182082 122448 182088 122460
rect 172664 122420 182088 122448
rect 172664 122408 172670 122420
rect 182082 122408 182088 122420
rect 182140 122408 182146 122460
rect 241422 122408 241428 122460
rect 241480 122448 241486 122460
rect 506750 122448 506756 122460
rect 241480 122420 506756 122448
rect 241480 122408 241486 122420
rect 506750 122408 506756 122420
rect 506808 122408 506814 122460
rect 82081 122383 82139 122389
rect 82081 122349 82093 122383
rect 82127 122380 82139 122383
rect 212534 122380 212540 122392
rect 82127 122352 212540 122380
rect 82127 122349 82139 122352
rect 82081 122343 82139 122349
rect 212534 122340 212540 122352
rect 212592 122340 212598 122392
rect 229002 122340 229008 122392
rect 229060 122380 229066 122392
rect 503717 122383 503775 122389
rect 503717 122380 503729 122383
rect 229060 122352 503729 122380
rect 229060 122340 229066 122352
rect 503717 122349 503729 122352
rect 503763 122349 503775 122383
rect 503717 122343 503775 122349
rect 80790 122272 80796 122324
rect 80848 122312 80854 122324
rect 223574 122312 223580 122324
rect 80848 122284 223580 122312
rect 80848 122272 80854 122284
rect 223574 122272 223580 122284
rect 223632 122272 223638 122324
rect 227622 122272 227628 122324
rect 227680 122312 227686 122324
rect 509050 122312 509056 122324
rect 227680 122284 509056 122312
rect 227680 122272 227686 122284
rect 509050 122272 509056 122284
rect 509108 122272 509114 122324
rect 80698 122204 80704 122256
rect 80756 122244 80762 122256
rect 205634 122244 205640 122256
rect 80756 122216 205640 122244
rect 80756 122204 80762 122216
rect 205634 122204 205640 122216
rect 205692 122204 205698 122256
rect 212442 122204 212448 122256
rect 212500 122244 212506 122256
rect 508774 122244 508780 122256
rect 212500 122216 508780 122244
rect 212500 122204 212506 122216
rect 508774 122204 508780 122216
rect 508832 122204 508838 122256
rect 82814 122136 82820 122188
rect 82872 122176 82878 122188
rect 196066 122176 196072 122188
rect 82872 122148 196072 122176
rect 82872 122136 82878 122148
rect 196066 122136 196072 122148
rect 196124 122136 196130 122188
rect 198642 122136 198648 122188
rect 198700 122176 198706 122188
rect 506934 122176 506940 122188
rect 198700 122148 506940 122176
rect 198700 122136 198706 122148
rect 506934 122136 506940 122148
rect 506992 122136 506998 122188
rect 78766 122068 78772 122120
rect 78824 122108 78830 122120
rect 393961 122111 394019 122117
rect 393961 122108 393973 122111
rect 78824 122080 393973 122108
rect 78824 122068 78830 122080
rect 393961 122077 393973 122080
rect 394007 122077 394019 122111
rect 393961 122071 394019 122077
rect 400122 122068 400128 122120
rect 400180 122108 400186 122120
rect 509878 122108 509884 122120
rect 400180 122080 509884 122108
rect 400180 122068 400186 122080
rect 509878 122068 509884 122080
rect 509936 122068 509942 122120
rect 80882 122000 80888 122052
rect 80940 122040 80946 122052
rect 99374 122040 99380 122052
rect 80940 122012 99380 122040
rect 80940 122000 80946 122012
rect 99374 122000 99380 122012
rect 99432 122000 99438 122052
rect 103514 122040 103520 122052
rect 103475 122012 103520 122040
rect 103514 122000 103520 122012
rect 103572 122000 103578 122052
rect 124306 122000 124312 122052
rect 124364 122040 124370 122052
rect 133782 122040 133788 122052
rect 124364 122012 133788 122040
rect 124364 122000 124370 122012
rect 133782 122000 133788 122012
rect 133840 122000 133846 122052
rect 143626 122000 143632 122052
rect 143684 122040 143690 122052
rect 153102 122040 153108 122052
rect 143684 122012 153108 122040
rect 143684 122000 143690 122012
rect 153102 122000 153108 122012
rect 153160 122000 153166 122052
rect 162946 122000 162952 122052
rect 163004 122040 163010 122052
rect 172422 122040 172428 122052
rect 163004 122012 172428 122040
rect 163004 122000 163010 122012
rect 172422 122000 172428 122012
rect 172480 122000 172486 122052
rect 172514 122000 172520 122052
rect 172572 122040 172578 122052
rect 172790 122040 172796 122052
rect 172572 122012 172796 122040
rect 172572 122000 172578 122012
rect 172790 122000 172796 122012
rect 172848 122000 172854 122052
rect 182358 122000 182364 122052
rect 182416 122040 182422 122052
rect 191742 122040 191748 122052
rect 182416 122012 191748 122040
rect 182416 122000 182422 122012
rect 191742 122000 191748 122012
rect 191800 122000 191806 122052
rect 240318 122000 240324 122052
rect 240376 122040 240382 122052
rect 241514 122040 241520 122052
rect 240376 122012 241520 122040
rect 240376 122000 240382 122012
rect 241514 122000 241520 122012
rect 241572 122000 241578 122052
rect 326982 122040 326988 122052
rect 326943 122012 326988 122040
rect 326982 122000 326988 122012
rect 327040 122000 327046 122052
rect 367002 122000 367008 122052
rect 367060 122040 367066 122052
rect 503162 122040 503168 122052
rect 367060 122012 503168 122040
rect 367060 122000 367066 122012
rect 503162 122000 503168 122012
rect 503220 122000 503226 122052
rect 86862 121932 86868 121984
rect 86920 121972 86926 121984
rect 95142 121972 95148 121984
rect 86920 121944 95148 121972
rect 86920 121932 86926 121944
rect 95142 121932 95148 121944
rect 95200 121932 95206 121984
rect 95326 121932 95332 121984
rect 95384 121972 95390 121984
rect 101030 121972 101036 121984
rect 95384 121944 101036 121972
rect 95384 121932 95390 121944
rect 101030 121932 101036 121944
rect 101088 121932 101094 121984
rect 376846 121932 376852 121984
rect 376904 121972 376910 121984
rect 386138 121972 386144 121984
rect 376904 121944 386144 121972
rect 376904 121932 376910 121944
rect 386138 121932 386144 121944
rect 386196 121932 386202 121984
rect 393958 121972 393964 121984
rect 393919 121944 393964 121972
rect 393958 121932 393964 121944
rect 394016 121932 394022 121984
rect 404446 121932 404452 121984
rect 404504 121972 404510 121984
rect 413922 121972 413928 121984
rect 404504 121944 413928 121972
rect 404504 121932 404510 121944
rect 413922 121932 413928 121944
rect 413980 121932 413986 121984
rect 415762 121932 415768 121984
rect 415820 121972 415826 121984
rect 424962 121972 424968 121984
rect 415820 121944 424968 121972
rect 415820 121932 415826 121944
rect 424962 121932 424968 121944
rect 425020 121932 425026 121984
rect 440142 121932 440148 121984
rect 440200 121972 440206 121984
rect 511534 121972 511540 121984
rect 440200 121944 511540 121972
rect 440200 121932 440206 121944
rect 511534 121932 511540 121944
rect 511592 121932 511598 121984
rect 95234 121864 95240 121916
rect 95292 121904 95298 121916
rect 105354 121904 105360 121916
rect 95292 121876 105360 121904
rect 95292 121864 95298 121876
rect 105354 121864 105360 121876
rect 105412 121864 105418 121916
rect 469122 121864 469128 121916
rect 469180 121904 469186 121916
rect 503438 121904 503444 121916
rect 469180 121876 503444 121904
rect 469180 121864 469186 121876
rect 503438 121864 503444 121876
rect 503496 121864 503502 121916
rect 79686 121796 79692 121848
rect 79744 121836 79750 121848
rect 84930 121836 84936 121848
rect 79744 121808 84936 121836
rect 79744 121796 79750 121808
rect 84930 121796 84936 121808
rect 84988 121796 84994 121848
rect 90634 121796 90640 121848
rect 90692 121836 90698 121848
rect 129734 121836 129740 121848
rect 90692 121808 129740 121836
rect 90692 121796 90698 121808
rect 129734 121796 129740 121808
rect 129792 121796 129798 121848
rect 338114 121796 338120 121848
rect 338172 121836 338178 121848
rect 342990 121836 342996 121848
rect 338172 121808 342996 121836
rect 338172 121796 338178 121808
rect 342990 121796 342996 121808
rect 343048 121796 343054 121848
rect 484302 121796 484308 121848
rect 484360 121836 484366 121848
rect 498197 121839 498255 121845
rect 498197 121836 498209 121839
rect 484360 121808 498209 121836
rect 484360 121796 484366 121808
rect 498197 121805 498209 121808
rect 498243 121805 498255 121839
rect 498197 121799 498255 121805
rect 498289 121839 498347 121845
rect 498289 121805 498301 121839
rect 498335 121836 498347 121839
rect 505370 121836 505376 121848
rect 498335 121808 505376 121836
rect 498335 121805 498347 121808
rect 498289 121799 498347 121805
rect 505370 121796 505376 121808
rect 505428 121796 505434 121848
rect 78858 121728 78864 121780
rect 78916 121768 78922 121780
rect 82081 121771 82139 121777
rect 82081 121768 82093 121771
rect 78916 121740 82093 121768
rect 78916 121728 78922 121740
rect 82081 121737 82093 121740
rect 82127 121737 82139 121771
rect 82081 121731 82139 121737
rect 82449 121771 82507 121777
rect 82449 121737 82461 121771
rect 82495 121768 82507 121771
rect 84105 121771 84163 121777
rect 84105 121768 84117 121771
rect 82495 121740 84117 121768
rect 82495 121737 82507 121740
rect 82449 121731 82507 121737
rect 84105 121737 84117 121740
rect 84151 121737 84163 121771
rect 84105 121731 84163 121737
rect 92290 121728 92296 121780
rect 92348 121768 92354 121780
rect 123018 121768 123024 121780
rect 92348 121740 123024 121768
rect 92348 121728 92354 121740
rect 123018 121728 123024 121740
rect 123076 121728 123082 121780
rect 330938 121728 330944 121780
rect 330996 121768 331002 121780
rect 336642 121768 336648 121780
rect 330996 121740 336648 121768
rect 330996 121728 331002 121740
rect 336642 121728 336648 121740
rect 336700 121728 336706 121780
rect 480162 121728 480168 121780
rect 480220 121768 480226 121780
rect 502613 121771 502671 121777
rect 502613 121768 502625 121771
rect 480220 121740 502625 121768
rect 480220 121728 480226 121740
rect 502613 121737 502625 121740
rect 502659 121737 502671 121771
rect 502613 121731 502671 121737
rect 78214 121660 78220 121712
rect 78272 121700 78278 121712
rect 111058 121700 111064 121712
rect 78272 121672 111064 121700
rect 78272 121660 78278 121672
rect 111058 121660 111064 121672
rect 111116 121660 111122 121712
rect 338114 121660 338120 121712
rect 338172 121700 338178 121712
rect 338172 121672 338217 121700
rect 338172 121660 338178 121672
rect 491294 121660 491300 121712
rect 491352 121700 491358 121712
rect 492306 121700 492312 121712
rect 491352 121672 492312 121700
rect 491352 121660 491358 121672
rect 492306 121660 492312 121672
rect 492364 121660 492370 121712
rect 493318 121660 493324 121712
rect 493376 121700 493382 121712
rect 498197 121703 498255 121709
rect 498197 121700 498209 121703
rect 493376 121672 498209 121700
rect 493376 121660 493382 121672
rect 498197 121669 498209 121672
rect 498243 121669 498255 121703
rect 498197 121663 498255 121669
rect 498470 121660 498476 121712
rect 498528 121700 498534 121712
rect 499298 121700 499304 121712
rect 498528 121672 499304 121700
rect 498528 121660 498534 121672
rect 499298 121660 499304 121672
rect 499356 121660 499362 121712
rect 499393 121703 499451 121709
rect 499393 121669 499405 121703
rect 499439 121700 499451 121703
rect 507302 121700 507308 121712
rect 499439 121672 507308 121700
rect 499439 121669 499451 121672
rect 499393 121663 499451 121669
rect 507302 121660 507308 121672
rect 507360 121660 507366 121712
rect 9582 121592 9588 121644
rect 9640 121632 9646 121644
rect 175274 121632 175280 121644
rect 9640 121604 175280 121632
rect 9640 121592 9646 121604
rect 175274 121592 175280 121604
rect 175332 121592 175338 121644
rect 399386 121592 399392 121644
rect 399444 121632 399450 121644
rect 498289 121635 498347 121641
rect 498289 121632 498301 121635
rect 399444 121604 498301 121632
rect 399444 121592 399450 121604
rect 498289 121601 498301 121604
rect 498335 121601 498347 121635
rect 498289 121595 498347 121601
rect 498381 121635 498439 121641
rect 498381 121601 498393 121635
rect 498427 121632 498439 121635
rect 506842 121632 506848 121644
rect 498427 121604 506848 121632
rect 498427 121601 498439 121604
rect 498381 121595 498439 121601
rect 506842 121592 506848 121604
rect 506900 121592 506906 121644
rect 3510 121524 3516 121576
rect 3568 121564 3574 121576
rect 277762 121564 277768 121576
rect 3568 121536 277768 121564
rect 3568 121524 3574 121536
rect 277762 121524 277768 121536
rect 277820 121524 277826 121576
rect 377858 121524 377864 121576
rect 377916 121564 377922 121576
rect 507210 121564 507216 121576
rect 377916 121536 507216 121564
rect 377916 121524 377922 121536
rect 507210 121524 507216 121536
rect 507268 121524 507274 121576
rect 79597 121499 79655 121505
rect 79597 121465 79609 121499
rect 79643 121496 79655 121499
rect 79686 121496 79692 121508
rect 79643 121468 79692 121496
rect 79643 121465 79655 121468
rect 79597 121459 79655 121465
rect 79686 121456 79692 121468
rect 79744 121456 79750 121508
rect 81897 121499 81955 121505
rect 81897 121465 81909 121499
rect 81943 121496 81955 121499
rect 445846 121496 445852 121508
rect 81943 121468 445852 121496
rect 81943 121465 81955 121468
rect 81897 121459 81955 121465
rect 445846 121456 445852 121468
rect 445904 121456 445910 121508
rect 496078 121456 496084 121508
rect 496136 121496 496142 121508
rect 501877 121499 501935 121505
rect 501877 121496 501889 121499
rect 496136 121468 501889 121496
rect 496136 121456 496142 121468
rect 501877 121465 501889 121468
rect 501923 121465 501935 121499
rect 501877 121459 501935 121465
rect 507302 121456 507308 121508
rect 507360 121496 507366 121508
rect 510522 121496 510528 121508
rect 507360 121468 510528 121496
rect 507360 121456 507366 121468
rect 510522 121456 510528 121468
rect 510580 121456 510586 121508
rect 9306 121388 9312 121440
rect 9364 121428 9370 121440
rect 494514 121428 494520 121440
rect 9364 121400 494520 121428
rect 9364 121388 9370 121400
rect 494514 121388 494520 121400
rect 494572 121388 494578 121440
rect 499390 121388 499396 121440
rect 499448 121428 499454 121440
rect 501509 121431 501567 121437
rect 501509 121428 501521 121431
rect 499448 121400 501521 121428
rect 499448 121388 499454 121400
rect 501509 121397 501521 121400
rect 501555 121397 501567 121431
rect 501509 121391 501567 121397
rect 509878 121388 509884 121440
rect 509936 121428 509942 121440
rect 511626 121428 511632 121440
rect 509936 121400 511632 121428
rect 509936 121388 509942 121400
rect 511626 121388 511632 121400
rect 511684 121388 511690 121440
rect 8846 121320 8852 121372
rect 8904 121360 8910 121372
rect 454034 121360 454040 121372
rect 8904 121332 454040 121360
rect 8904 121320 8910 121332
rect 454034 121320 454040 121332
rect 454092 121320 454098 121372
rect 456702 121320 456708 121372
rect 456760 121360 456766 121372
rect 502886 121360 502892 121372
rect 456760 121332 502892 121360
rect 456760 121320 456766 121332
rect 502886 121320 502892 121332
rect 502944 121320 502950 121372
rect 42242 121252 42248 121304
rect 42300 121292 42306 121304
rect 465994 121292 466000 121304
rect 42300 121264 466000 121292
rect 42300 121252 42306 121264
rect 465994 121252 466000 121264
rect 466052 121252 466058 121304
rect 488442 121252 488448 121304
rect 488500 121292 488506 121304
rect 499758 121292 499764 121304
rect 488500 121264 499764 121292
rect 488500 121252 488506 121264
rect 499758 121252 499764 121264
rect 499816 121252 499822 121304
rect 502794 121292 502800 121304
rect 499868 121264 502800 121292
rect 24762 121184 24768 121236
rect 24820 121224 24826 121236
rect 427906 121224 427912 121236
rect 24820 121196 427912 121224
rect 24820 121184 24826 121196
rect 427906 121184 427912 121196
rect 427964 121184 427970 121236
rect 431862 121184 431868 121236
rect 431920 121224 431926 121236
rect 499868 121224 499896 121264
rect 502794 121252 502800 121264
rect 502852 121252 502858 121304
rect 431920 121196 499896 121224
rect 431920 121184 431926 121196
rect 499942 121184 499948 121236
rect 500000 121224 500006 121236
rect 501782 121224 501788 121236
rect 500000 121196 501788 121224
rect 500000 121184 500006 121196
rect 501782 121184 501788 121196
rect 501840 121184 501846 121236
rect 3694 121116 3700 121168
rect 3752 121156 3758 121168
rect 173066 121156 173072 121168
rect 3752 121128 173072 121156
rect 3752 121116 3758 121128
rect 173066 121116 173072 121128
rect 173124 121116 173130 121168
rect 189626 121116 189632 121168
rect 189684 121156 189690 121168
rect 580626 121156 580632 121168
rect 189684 121128 580632 121156
rect 189684 121116 189690 121128
rect 580626 121116 580632 121128
rect 580684 121116 580690 121168
rect 82081 121091 82139 121097
rect 82081 121057 82093 121091
rect 82127 121088 82139 121091
rect 85022 121088 85028 121100
rect 82127 121060 85028 121088
rect 82127 121057 82139 121060
rect 82081 121051 82139 121057
rect 85022 121048 85028 121060
rect 85080 121048 85086 121100
rect 392210 121048 392216 121100
rect 392268 121088 392274 121100
rect 499025 121091 499083 121097
rect 499025 121088 499037 121091
rect 392268 121060 499037 121088
rect 392268 121048 392274 121060
rect 499025 121057 499037 121060
rect 499071 121057 499083 121091
rect 499025 121051 499083 121057
rect 500034 121048 500040 121100
rect 500092 121088 500098 121100
rect 501601 121091 501659 121097
rect 501601 121088 501613 121091
rect 500092 121060 501613 121088
rect 500092 121048 500098 121060
rect 501601 121057 501613 121060
rect 501647 121057 501659 121091
rect 501601 121051 501659 121057
rect 501693 121091 501751 121097
rect 501693 121057 501705 121091
rect 501739 121088 501751 121091
rect 511810 121088 511816 121100
rect 501739 121060 511816 121088
rect 501739 121057 501751 121060
rect 501693 121051 501751 121057
rect 511810 121048 511816 121060
rect 511868 121048 511874 121100
rect 33778 120980 33784 121032
rect 33836 121020 33842 121032
rect 127802 121020 127808 121032
rect 33836 120992 127808 121020
rect 33836 120980 33842 120992
rect 127802 120980 127808 120992
rect 127860 120980 127866 121032
rect 144362 120980 144368 121032
rect 144420 121020 144426 121032
rect 506106 121020 506112 121032
rect 144420 120992 506112 121020
rect 144420 120980 144426 120992
rect 506106 120980 506112 120992
rect 506164 120980 506170 121032
rect 3418 120912 3424 120964
rect 3476 120952 3482 120964
rect 146754 120952 146760 120964
rect 3476 120924 146760 120952
rect 3476 120912 3482 120924
rect 146754 120912 146760 120924
rect 146812 120912 146818 120964
rect 165890 120912 165896 120964
rect 165948 120952 165954 120964
rect 505738 120952 505744 120964
rect 165948 120924 505744 120952
rect 165948 120912 165954 120924
rect 505738 120912 505744 120924
rect 505796 120912 505802 120964
rect 9398 120844 9404 120896
rect 9456 120884 9462 120896
rect 337378 120884 337384 120896
rect 9456 120856 337384 120884
rect 9456 120844 9462 120856
rect 337378 120844 337384 120856
rect 337436 120844 337442 120896
rect 349062 120844 349068 120896
rect 349120 120884 349126 120896
rect 511902 120884 511908 120896
rect 349120 120856 511908 120884
rect 349120 120844 349126 120856
rect 511902 120844 511908 120856
rect 511960 120844 511966 120896
rect 42150 120776 42156 120828
rect 42208 120816 42214 120828
rect 163498 120816 163504 120828
rect 42208 120788 163504 120816
rect 42208 120776 42214 120788
rect 163498 120776 163504 120788
rect 163556 120776 163562 120828
rect 239674 120776 239680 120828
rect 239732 120816 239738 120828
rect 506198 120816 506204 120828
rect 239732 120788 506204 120816
rect 239732 120776 239738 120788
rect 506198 120776 506204 120788
rect 506256 120776 506262 120828
rect 77294 120708 77300 120760
rect 77352 120748 77358 120760
rect 313458 120748 313464 120760
rect 77352 120720 313464 120748
rect 77352 120708 77358 120720
rect 313458 120708 313464 120720
rect 313516 120708 313522 120760
rect 318242 120708 318248 120760
rect 318300 120748 318306 120760
rect 580442 120748 580448 120760
rect 318300 120720 580448 120748
rect 318300 120708 318306 120720
rect 580442 120708 580448 120720
rect 580500 120708 580506 120760
rect 79042 120640 79048 120692
rect 79100 120680 79106 120692
rect 150618 120680 150624 120692
rect 79100 120652 150624 120680
rect 79100 120640 79106 120652
rect 150618 120640 150624 120652
rect 150676 120640 150682 120692
rect 274542 120640 274548 120692
rect 274600 120680 274606 120692
rect 496817 120683 496875 120689
rect 496817 120680 496829 120683
rect 274600 120652 496829 120680
rect 274600 120640 274606 120652
rect 496817 120649 496829 120652
rect 496863 120649 496875 120683
rect 498930 120680 498936 120692
rect 496817 120643 496875 120649
rect 496924 120652 498936 120680
rect 82817 120615 82875 120621
rect 82817 120581 82829 120615
rect 82863 120612 82875 120615
rect 84010 120612 84016 120624
rect 82863 120584 84016 120612
rect 82863 120581 82875 120584
rect 82817 120575 82875 120581
rect 84010 120572 84016 120584
rect 84068 120572 84074 120624
rect 84105 120615 84163 120621
rect 84105 120581 84117 120615
rect 84151 120612 84163 120615
rect 118418 120612 118424 120624
rect 84151 120584 118424 120612
rect 84151 120581 84163 120584
rect 84105 120575 84163 120581
rect 118418 120572 118424 120584
rect 118476 120572 118482 120624
rect 284938 120572 284944 120624
rect 284996 120612 285002 120624
rect 496924 120612 496952 120652
rect 498930 120640 498936 120652
rect 498988 120640 498994 120692
rect 499025 120683 499083 120689
rect 499025 120649 499037 120683
rect 499071 120680 499083 120683
rect 507118 120680 507124 120692
rect 499071 120652 507124 120680
rect 499071 120649 499083 120652
rect 499025 120643 499083 120649
rect 507118 120640 507124 120652
rect 507176 120640 507182 120692
rect 284996 120584 496952 120612
rect 497001 120615 497059 120621
rect 284996 120572 285002 120584
rect 497001 120581 497013 120615
rect 497047 120612 497059 120615
rect 506658 120612 506664 120624
rect 497047 120584 506664 120612
rect 497047 120581 497059 120584
rect 497001 120575 497059 120581
rect 506658 120572 506664 120584
rect 506716 120572 506722 120624
rect 80974 120504 80980 120556
rect 81032 120544 81038 120556
rect 110417 120547 110475 120553
rect 110417 120544 110429 120547
rect 81032 120516 110429 120544
rect 81032 120504 81038 120516
rect 110417 120513 110429 120516
rect 110463 120513 110475 120547
rect 110417 120507 110475 120513
rect 304902 120504 304908 120556
rect 304960 120544 304966 120556
rect 509694 120544 509700 120556
rect 304960 120516 509700 120544
rect 304960 120504 304966 120516
rect 509694 120504 509700 120516
rect 509752 120504 509758 120556
rect 82909 120479 82967 120485
rect 82909 120445 82921 120479
rect 82955 120476 82967 120479
rect 106458 120476 106464 120488
rect 82955 120448 106464 120476
rect 82955 120445 82967 120448
rect 82909 120439 82967 120445
rect 106458 120436 106464 120448
rect 106516 120436 106522 120488
rect 329742 120436 329748 120488
rect 329800 120476 329806 120488
rect 501601 120479 501659 120485
rect 501601 120476 501613 120479
rect 329800 120448 501613 120476
rect 329800 120436 329806 120448
rect 501601 120445 501613 120448
rect 501647 120445 501659 120479
rect 501601 120439 501659 120445
rect 393222 120368 393228 120420
rect 393280 120408 393286 120420
rect 510430 120408 510436 120420
rect 393280 120380 510436 120408
rect 393280 120368 393286 120380
rect 510430 120368 510436 120380
rect 510488 120368 510494 120420
rect 31110 120300 31116 120352
rect 31168 120340 31174 120352
rect 401594 120340 401600 120352
rect 31168 120312 401600 120340
rect 31168 120300 31174 120312
rect 401594 120300 401600 120312
rect 401652 120300 401658 120352
rect 501601 120343 501659 120349
rect 501601 120309 501613 120343
rect 501647 120340 501659 120343
rect 508498 120340 508504 120352
rect 501647 120312 508504 120340
rect 501647 120309 501659 120312
rect 501601 120303 501659 120309
rect 508498 120300 508504 120312
rect 508556 120300 508562 120352
rect 15102 120028 15108 120080
rect 15160 120068 15166 120080
rect 137186 120068 137192 120080
rect 15160 120040 137192 120068
rect 15160 120028 15166 120040
rect 137186 120028 137192 120040
rect 137244 120028 137250 120080
rect 149146 120028 149152 120080
rect 149204 120068 149210 120080
rect 150342 120068 150348 120080
rect 149204 120040 150348 120068
rect 149204 120028 149210 120040
rect 150342 120028 150348 120040
rect 150400 120028 150406 120080
rect 199194 120028 199200 120080
rect 199252 120068 199258 120080
rect 200022 120068 200028 120080
rect 199252 120040 200028 120068
rect 199252 120028 199258 120040
rect 200022 120028 200028 120040
rect 200080 120028 200086 120080
rect 201586 120028 201592 120080
rect 201644 120068 201650 120080
rect 225046 120068 225052 120080
rect 201644 120040 225052 120068
rect 201644 120028 201650 120040
rect 225046 120028 225052 120040
rect 225104 120028 225110 120080
rect 244458 120028 244464 120080
rect 244516 120068 244522 120080
rect 245562 120068 245568 120080
rect 244516 120040 245568 120068
rect 244516 120028 244522 120040
rect 245562 120028 245568 120040
rect 245620 120028 245626 120080
rect 251082 120028 251088 120080
rect 251140 120068 251146 120080
rect 496906 120068 496912 120080
rect 251140 120040 496912 120068
rect 251140 120028 251146 120040
rect 496906 120028 496912 120040
rect 496964 120028 496970 120080
rect 84746 119960 84752 120012
rect 84804 120000 84810 120012
rect 242894 120000 242900 120012
rect 84804 119972 242900 120000
rect 84804 119960 84810 119972
rect 242894 119960 242900 119972
rect 242952 119960 242958 120012
rect 261202 119960 261208 120012
rect 261260 120000 261266 120012
rect 262122 120000 262128 120012
rect 261260 119972 262128 120000
rect 261260 119960 261266 119972
rect 262122 119960 262128 119972
rect 262180 119960 262186 120012
rect 265802 119960 265808 120012
rect 265860 120000 265866 120012
rect 511629 120003 511687 120009
rect 511629 120000 511641 120003
rect 265860 119972 511641 120000
rect 265860 119960 265866 119972
rect 511629 119969 511641 119972
rect 511675 119969 511687 120003
rect 511629 119963 511687 119969
rect 22002 119892 22008 119944
rect 22060 119932 22066 119944
rect 156322 119932 156328 119944
rect 22060 119904 156328 119932
rect 22060 119892 22066 119904
rect 156322 119892 156328 119904
rect 156380 119892 156386 119944
rect 179322 119892 179328 119944
rect 179380 119932 179386 119944
rect 430298 119932 430304 119944
rect 179380 119904 430304 119932
rect 179380 119892 179386 119904
rect 430298 119892 430304 119904
rect 430356 119892 430362 119944
rect 437474 119892 437480 119944
rect 437532 119932 437538 119944
rect 438762 119932 438768 119944
rect 437532 119904 438768 119932
rect 437532 119892 437538 119904
rect 438762 119892 438768 119904
rect 438820 119892 438826 119944
rect 461210 119892 461216 119944
rect 461268 119932 461274 119944
rect 508130 119932 508136 119944
rect 461268 119904 508136 119932
rect 461268 119892 461274 119904
rect 508130 119892 508136 119904
rect 508188 119892 508194 119944
rect 17218 119824 17224 119876
rect 17276 119864 17282 119876
rect 270586 119864 270592 119876
rect 17276 119836 270592 119864
rect 17276 119824 17282 119836
rect 270586 119824 270592 119836
rect 270644 119824 270650 119876
rect 275370 119824 275376 119876
rect 275428 119864 275434 119876
rect 522298 119864 522304 119876
rect 275428 119836 522304 119864
rect 275428 119824 275434 119836
rect 522298 119824 522304 119836
rect 522356 119824 522362 119876
rect 71682 119756 71688 119808
rect 71740 119796 71746 119808
rect 234890 119796 234896 119808
rect 71740 119768 234896 119796
rect 71740 119756 71746 119768
rect 234890 119756 234896 119768
rect 234948 119756 234954 119808
rect 242066 119756 242072 119808
rect 242124 119796 242130 119808
rect 495434 119796 495440 119808
rect 242124 119768 495440 119796
rect 242124 119756 242130 119768
rect 495434 119756 495440 119768
rect 495492 119756 495498 119808
rect 51810 119688 51816 119740
rect 51868 119728 51874 119740
rect 306466 119728 306472 119740
rect 51868 119700 306472 119728
rect 51868 119688 51874 119700
rect 306466 119688 306472 119700
rect 306524 119688 306530 119740
rect 311066 119688 311072 119740
rect 311124 119728 311130 119740
rect 349154 119728 349160 119740
rect 311124 119700 349160 119728
rect 311124 119688 311130 119700
rect 349154 119688 349160 119700
rect 349212 119688 349218 119740
rect 352558 119688 352564 119740
rect 352616 119728 352622 119740
rect 356330 119728 356336 119740
rect 352616 119700 356336 119728
rect 352616 119688 352622 119700
rect 356330 119688 356336 119700
rect 356388 119688 356394 119740
rect 363506 119688 363512 119740
rect 363564 119728 363570 119740
rect 519630 119728 519636 119740
rect 363564 119700 519636 119728
rect 363564 119688 363570 119700
rect 519630 119688 519636 119700
rect 519688 119688 519694 119740
rect 59262 119620 59268 119672
rect 59320 119660 59326 119672
rect 227714 119660 227720 119672
rect 59320 119632 227720 119660
rect 59320 119620 59326 119632
rect 227714 119620 227720 119632
rect 227772 119620 227778 119672
rect 230106 119620 230112 119672
rect 230164 119660 230170 119672
rect 489181 119663 489239 119669
rect 489181 119660 489193 119663
rect 230164 119632 489193 119660
rect 230164 119620 230170 119632
rect 489181 119629 489193 119632
rect 489227 119629 489239 119663
rect 489181 119623 489239 119629
rect 489914 119620 489920 119672
rect 489972 119660 489978 119672
rect 491202 119660 491208 119672
rect 489972 119632 491208 119660
rect 489972 119620 489978 119632
rect 491202 119620 491208 119632
rect 491260 119620 491266 119672
rect 80606 119552 80612 119604
rect 80664 119592 80670 119604
rect 86313 119595 86371 119601
rect 86313 119592 86325 119595
rect 80664 119564 86325 119592
rect 80664 119552 80670 119564
rect 86313 119561 86325 119564
rect 86359 119561 86371 119595
rect 86313 119555 86371 119561
rect 103882 119552 103888 119604
rect 103940 119592 103946 119604
rect 104802 119592 104808 119604
rect 103940 119564 104808 119592
rect 103940 119552 103946 119564
rect 104802 119552 104808 119564
rect 104860 119552 104866 119604
rect 106274 119552 106280 119604
rect 106332 119592 106338 119604
rect 107470 119592 107476 119604
rect 106332 119564 107476 119592
rect 106332 119552 106338 119564
rect 107470 119552 107476 119564
rect 107528 119552 107534 119604
rect 107565 119595 107623 119601
rect 107565 119561 107577 119595
rect 107611 119592 107623 119595
rect 382642 119592 382648 119604
rect 107611 119564 382648 119592
rect 107611 119561 107623 119564
rect 107565 119555 107623 119561
rect 382642 119552 382648 119564
rect 382700 119552 382706 119604
rect 391842 119552 391848 119604
rect 391900 119592 391906 119604
rect 473170 119592 473176 119604
rect 391900 119564 473176 119592
rect 391900 119552 391906 119564
rect 473170 119552 473176 119564
rect 473228 119552 473234 119604
rect 479518 119552 479524 119604
rect 479576 119592 479582 119604
rect 509970 119592 509976 119604
rect 479576 119564 509976 119592
rect 479576 119552 479582 119564
rect 509970 119552 509976 119564
rect 510028 119552 510034 119604
rect 28902 119484 28908 119536
rect 28960 119524 28966 119536
rect 194410 119524 194416 119536
rect 28960 119496 194416 119524
rect 28960 119484 28966 119496
rect 194410 119484 194416 119496
rect 194468 119484 194474 119536
rect 211154 119484 211160 119536
rect 211212 119524 211218 119536
rect 212350 119524 212356 119536
rect 211212 119496 212356 119524
rect 211212 119484 211218 119496
rect 212350 119484 212356 119496
rect 212408 119484 212414 119536
rect 212445 119527 212503 119533
rect 212445 119493 212457 119527
rect 212491 119524 212503 119527
rect 509142 119524 509148 119536
rect 212491 119496 509148 119524
rect 212491 119493 212503 119496
rect 212445 119487 212503 119493
rect 509142 119484 509148 119496
rect 509200 119484 509206 119536
rect 46290 119416 46296 119468
rect 46348 119456 46354 119468
rect 82722 119456 82728 119468
rect 46348 119428 82584 119456
rect 82683 119428 82728 119456
rect 46348 119416 46354 119428
rect 20622 119348 20628 119400
rect 20680 119388 20686 119400
rect 82449 119391 82507 119397
rect 82449 119388 82461 119391
rect 20680 119360 82461 119388
rect 20680 119348 20686 119360
rect 82449 119357 82461 119360
rect 82495 119357 82507 119391
rect 82556 119388 82584 119428
rect 82722 119416 82728 119428
rect 82780 119416 82786 119468
rect 425514 119456 425520 119468
rect 82832 119428 425520 119456
rect 82832 119388 82860 119428
rect 425514 119416 425520 119428
rect 425572 119416 425578 119468
rect 463602 119416 463608 119468
rect 463660 119456 463666 119468
rect 471238 119456 471244 119468
rect 463660 119428 471244 119456
rect 463660 119416 463666 119428
rect 471238 119416 471244 119428
rect 471296 119416 471302 119468
rect 476758 119416 476764 119468
rect 476816 119456 476822 119468
rect 510338 119456 510344 119468
rect 476816 119428 510344 119456
rect 476816 119416 476822 119428
rect 510338 119416 510344 119428
rect 510396 119416 510402 119468
rect 82556 119360 82860 119388
rect 83461 119391 83519 119397
rect 82449 119351 82507 119357
rect 83461 119357 83473 119391
rect 83507 119388 83519 119391
rect 91922 119388 91928 119400
rect 83507 119360 91928 119388
rect 83507 119357 83519 119360
rect 83461 119351 83519 119357
rect 91922 119348 91928 119360
rect 91980 119348 91986 119400
rect 94314 119348 94320 119400
rect 94372 119388 94378 119400
rect 473354 119388 473360 119400
rect 94372 119360 473360 119388
rect 94372 119348 94378 119360
rect 473354 119348 473360 119360
rect 473412 119348 473418 119400
rect 489181 119391 489239 119397
rect 489181 119357 489193 119391
rect 489227 119388 489239 119391
rect 492674 119388 492680 119400
rect 489227 119360 492680 119388
rect 489227 119357 489239 119360
rect 489181 119351 489239 119357
rect 492674 119348 492680 119360
rect 492732 119348 492738 119400
rect 492769 119391 492827 119397
rect 492769 119357 492781 119391
rect 492815 119388 492827 119391
rect 571334 119388 571340 119400
rect 492815 119360 571340 119388
rect 492815 119357 492827 119360
rect 492769 119351 492827 119357
rect 571334 119348 571340 119360
rect 571392 119348 571398 119400
rect 38470 119280 38476 119332
rect 38528 119320 38534 119332
rect 151538 119320 151544 119332
rect 38528 119292 151544 119320
rect 38528 119280 38534 119292
rect 151538 119280 151544 119292
rect 151596 119280 151602 119332
rect 161293 119323 161351 119329
rect 161293 119289 161305 119323
rect 161339 119320 161351 119323
rect 365898 119320 365904 119332
rect 161339 119292 365904 119320
rect 161339 119289 161351 119292
rect 161293 119283 161351 119289
rect 365898 119280 365904 119292
rect 365956 119280 365962 119332
rect 373074 119280 373080 119332
rect 373132 119320 373138 119332
rect 373902 119320 373908 119332
rect 373132 119292 373908 119320
rect 373132 119280 373138 119292
rect 373902 119280 373908 119292
rect 373960 119280 373966 119332
rect 380250 119280 380256 119332
rect 380308 119320 380314 119332
rect 441706 119320 441712 119332
rect 380308 119292 441712 119320
rect 380308 119280 380314 119292
rect 441706 119280 441712 119292
rect 441764 119280 441770 119332
rect 467742 119280 467748 119332
rect 467800 119320 467806 119332
rect 480346 119320 480352 119332
rect 467800 119292 480352 119320
rect 467800 119280 467806 119292
rect 480346 119280 480352 119292
rect 480404 119280 480410 119332
rect 487062 119280 487068 119332
rect 487120 119320 487126 119332
rect 501506 119320 501512 119332
rect 487120 119292 501512 119320
rect 487120 119280 487126 119292
rect 501506 119280 501512 119292
rect 501564 119280 501570 119332
rect 82449 119255 82507 119261
rect 82449 119221 82461 119255
rect 82495 119252 82507 119255
rect 83461 119255 83519 119261
rect 83461 119252 83473 119255
rect 82495 119224 83473 119252
rect 82495 119221 82507 119224
rect 82449 119215 82507 119221
rect 83461 119221 83473 119224
rect 83507 119221 83519 119255
rect 83461 119215 83519 119221
rect 83642 119212 83648 119264
rect 83700 119252 83706 119264
rect 87322 119252 87328 119264
rect 83700 119224 87328 119252
rect 83700 119212 83706 119224
rect 87322 119212 87328 119224
rect 87380 119212 87386 119264
rect 102042 119212 102048 119264
rect 102100 119252 102106 119264
rect 107565 119255 107623 119261
rect 107565 119252 107577 119255
rect 102100 119224 107577 119252
rect 102100 119212 102106 119224
rect 107565 119221 107577 119224
rect 107611 119221 107623 119255
rect 107565 119215 107623 119221
rect 113450 119212 113456 119264
rect 113508 119252 113514 119264
rect 114462 119252 114468 119264
rect 113508 119224 114468 119252
rect 113508 119212 113514 119224
rect 114462 119212 114468 119224
rect 114520 119212 114526 119264
rect 114557 119255 114615 119261
rect 114557 119221 114569 119255
rect 114603 119252 114615 119255
rect 232498 119252 232504 119264
rect 114603 119224 232504 119252
rect 114603 119221 114615 119224
rect 114557 119215 114615 119221
rect 232498 119212 232504 119224
rect 232556 119212 232562 119264
rect 240042 119212 240048 119264
rect 240100 119252 240106 119264
rect 249061 119255 249119 119261
rect 249061 119252 249073 119255
rect 240100 119224 249073 119252
rect 240100 119212 240106 119224
rect 249061 119221 249073 119224
rect 249107 119221 249119 119255
rect 249061 119215 249119 119221
rect 249153 119255 249211 119261
rect 249153 119221 249165 119255
rect 249199 119252 249211 119255
rect 449250 119252 449256 119264
rect 249199 119224 449256 119252
rect 249199 119221 249211 119224
rect 249153 119215 249211 119221
rect 449250 119212 449256 119224
rect 449308 119212 449314 119264
rect 487522 119212 487528 119264
rect 487580 119252 487586 119264
rect 492769 119255 492827 119261
rect 492769 119252 492781 119255
rect 487580 119224 492781 119252
rect 487580 119212 487586 119224
rect 492769 119221 492781 119224
rect 492815 119221 492827 119255
rect 492769 119215 492827 119221
rect 92382 119144 92388 119196
rect 92440 119184 92446 119196
rect 208762 119184 208768 119196
rect 92440 119156 208768 119184
rect 92440 119144 92446 119156
rect 208762 119144 208768 119156
rect 208820 119144 208826 119196
rect 211062 119144 211068 119196
rect 211120 119184 211126 119196
rect 212445 119187 212503 119193
rect 212445 119184 212457 119187
rect 211120 119156 212457 119184
rect 211120 119144 211126 119156
rect 212445 119153 212457 119156
rect 212491 119153 212503 119187
rect 212445 119147 212503 119153
rect 218330 119144 218336 119196
rect 218388 119184 218394 119196
rect 219342 119184 219348 119196
rect 218388 119156 219348 119184
rect 218388 119144 218394 119156
rect 219342 119144 219348 119156
rect 219400 119144 219406 119196
rect 222930 119144 222936 119196
rect 222988 119184 222994 119196
rect 416774 119184 416780 119196
rect 222988 119156 416780 119184
rect 222988 119144 222994 119156
rect 416774 119144 416780 119156
rect 416832 119144 416838 119196
rect 500862 119144 500868 119196
rect 500920 119184 500926 119196
rect 501693 119187 501751 119193
rect 501693 119184 501705 119187
rect 500920 119156 501705 119184
rect 500920 119144 500926 119156
rect 501693 119153 501705 119156
rect 501739 119153 501751 119187
rect 501693 119147 501751 119153
rect 91002 119076 91008 119128
rect 91060 119116 91066 119128
rect 196802 119116 196808 119128
rect 91060 119088 196808 119116
rect 91060 119076 91066 119088
rect 196802 119076 196808 119088
rect 196860 119076 196866 119128
rect 206370 119076 206376 119128
rect 206428 119116 206434 119128
rect 396074 119116 396080 119128
rect 206428 119088 396080 119116
rect 206428 119076 206434 119088
rect 396074 119076 396080 119088
rect 396132 119076 396138 119128
rect 402238 119076 402244 119128
rect 402296 119116 402302 119128
rect 451642 119116 451648 119128
rect 402296 119088 451648 119116
rect 402296 119076 402302 119088
rect 451642 119076 451648 119088
rect 451700 119076 451706 119128
rect 78582 119008 78588 119060
rect 78640 119048 78646 119060
rect 161106 119048 161112 119060
rect 78640 119020 161112 119048
rect 78640 119008 78646 119020
rect 161106 119008 161112 119020
rect 161164 119008 161170 119060
rect 180058 119008 180064 119060
rect 180116 119048 180122 119060
rect 360194 119048 360200 119060
rect 180116 119020 360200 119048
rect 180116 119008 180122 119020
rect 360194 119008 360200 119020
rect 360252 119008 360258 119060
rect 384942 119008 384948 119060
rect 385000 119048 385006 119060
rect 447042 119048 447048 119060
rect 385000 119020 447048 119048
rect 385000 119008 385006 119020
rect 447042 119008 447048 119020
rect 447100 119008 447106 119060
rect 106182 118940 106188 118992
rect 106240 118980 106246 118992
rect 203978 118980 203984 118992
rect 106240 118952 203984 118980
rect 106240 118940 106246 118952
rect 203978 118940 203984 118952
rect 204036 118940 204042 118992
rect 233142 118940 233148 118992
rect 233200 118980 233206 118992
rect 301682 118980 301688 118992
rect 233200 118952 301688 118980
rect 233200 118940 233206 118952
rect 301682 118940 301688 118952
rect 301740 118940 301746 118992
rect 313918 118940 313924 118992
rect 313976 118980 313982 118992
rect 332594 118980 332600 118992
rect 313976 118952 332600 118980
rect 313976 118940 313982 118952
rect 332594 118940 332600 118952
rect 332652 118940 332658 118992
rect 355962 118940 355968 118992
rect 356020 118980 356026 118992
rect 509602 118980 509608 118992
rect 356020 118952 509608 118980
rect 356020 118940 356026 118952
rect 509602 118940 509608 118952
rect 509660 118940 509666 118992
rect 72970 118872 72976 118924
rect 73028 118912 73034 118924
rect 125410 118912 125416 118924
rect 73028 118884 125416 118912
rect 73028 118872 73034 118884
rect 125410 118872 125416 118884
rect 125468 118872 125474 118924
rect 246942 118872 246948 118924
rect 247000 118912 247006 118924
rect 248969 118915 249027 118921
rect 248969 118912 248981 118915
rect 247000 118884 248981 118912
rect 247000 118872 247006 118884
rect 248969 118881 248981 118884
rect 249015 118881 249027 118915
rect 248969 118875 249027 118881
rect 249061 118915 249119 118921
rect 249061 118881 249073 118915
rect 249107 118912 249119 118915
rect 375466 118912 375472 118924
rect 249107 118884 375472 118912
rect 249107 118881 249119 118884
rect 249061 118875 249119 118881
rect 375466 118872 375472 118884
rect 375524 118872 375530 118924
rect 407022 118872 407028 118924
rect 407080 118912 407086 118924
rect 423122 118912 423128 118924
rect 407080 118884 423128 118912
rect 407080 118872 407086 118884
rect 423122 118872 423128 118884
rect 423180 118872 423186 118924
rect 113082 118804 113088 118856
rect 113140 118844 113146 118856
rect 114557 118847 114615 118853
rect 114557 118844 114569 118847
rect 113140 118816 114569 118844
rect 113140 118804 113146 118816
rect 114557 118813 114569 118816
rect 114603 118813 114615 118847
rect 114557 118807 114615 118813
rect 120626 118804 120632 118856
rect 120684 118844 120690 118856
rect 169754 118844 169760 118856
rect 120684 118816 169760 118844
rect 120684 118804 120690 118816
rect 169754 118804 169760 118816
rect 169812 118804 169818 118856
rect 222102 118804 222108 118856
rect 222160 118844 222166 118856
rect 226337 118847 226395 118853
rect 226337 118844 226349 118847
rect 222160 118816 226349 118844
rect 222160 118804 222166 118816
rect 226337 118813 226349 118816
rect 226383 118813 226395 118847
rect 226337 118807 226395 118813
rect 237190 118804 237196 118856
rect 237248 118844 237254 118856
rect 304074 118844 304080 118856
rect 237248 118816 304080 118844
rect 237248 118804 237254 118816
rect 304074 118804 304080 118816
rect 304132 118804 304138 118856
rect 350537 118847 350595 118853
rect 350537 118813 350549 118847
rect 350583 118844 350595 118847
rect 433334 118844 433340 118856
rect 350583 118816 433340 118844
rect 350583 118813 350595 118816
rect 350537 118807 350595 118813
rect 433334 118804 433340 118816
rect 433392 118804 433398 118856
rect 435082 118804 435088 118856
rect 435140 118844 435146 118856
rect 436002 118844 436008 118856
rect 435140 118816 436008 118844
rect 435140 118804 435146 118816
rect 436002 118804 436008 118816
rect 436060 118804 436066 118856
rect 107562 118736 107568 118788
rect 107620 118776 107626 118788
rect 132402 118776 132408 118788
rect 107620 118748 132408 118776
rect 107620 118736 107626 118748
rect 132402 118736 132408 118748
rect 132460 118736 132466 118788
rect 201402 118736 201408 118788
rect 201460 118776 201466 118788
rect 268194 118776 268200 118788
rect 201460 118748 268200 118776
rect 201460 118736 201466 118748
rect 268194 118736 268200 118748
rect 268252 118736 268258 118788
rect 280154 118736 280160 118788
rect 280212 118776 280218 118788
rect 310514 118776 310520 118788
rect 280212 118748 310520 118776
rect 280212 118736 280218 118748
rect 310514 118736 310520 118748
rect 310572 118736 310578 118788
rect 344554 118736 344560 118788
rect 344612 118776 344618 118788
rect 419534 118776 419540 118788
rect 344612 118748 419540 118776
rect 344612 118736 344618 118748
rect 419534 118736 419540 118748
rect 419592 118736 419598 118788
rect 225322 118668 225328 118720
rect 225380 118708 225386 118720
rect 226242 118708 226248 118720
rect 225380 118680 226248 118708
rect 225380 118668 225386 118680
rect 226242 118668 226248 118680
rect 226300 118668 226306 118720
rect 226337 118711 226395 118717
rect 226337 118677 226349 118711
rect 226383 118708 226395 118711
rect 263594 118708 263600 118720
rect 226383 118680 261156 118708
rect 226383 118677 226395 118680
rect 226337 118671 226395 118677
rect 156046 118640 156052 118652
rect 156007 118612 156052 118640
rect 156046 118600 156052 118612
rect 156104 118600 156110 118652
rect 261128 118640 261156 118680
rect 262232 118680 263600 118708
rect 262232 118640 262260 118680
rect 263594 118668 263600 118680
rect 263652 118668 263658 118720
rect 307018 118668 307024 118720
rect 307076 118708 307082 118720
rect 315850 118708 315856 118720
rect 307076 118680 315856 118708
rect 307076 118668 307082 118680
rect 315850 118668 315856 118680
rect 315908 118668 315914 118720
rect 349338 118668 349344 118720
rect 349396 118708 349402 118720
rect 350537 118711 350595 118717
rect 350537 118708 350549 118711
rect 349396 118680 350549 118708
rect 349396 118668 349402 118680
rect 350537 118677 350549 118680
rect 350583 118677 350595 118711
rect 350537 118671 350595 118677
rect 368290 118668 368296 118720
rect 368348 118708 368354 118720
rect 369946 118708 369952 118720
rect 368348 118680 369952 118708
rect 368348 118668 368354 118680
rect 369946 118668 369952 118680
rect 370004 118668 370010 118720
rect 261128 118612 262260 118640
rect 81618 118532 81624 118584
rect 81676 118572 81682 118584
rect 258166 118572 258172 118584
rect 81676 118544 258172 118572
rect 81676 118532 81682 118544
rect 258166 118532 258172 118544
rect 258224 118532 258230 118584
rect 502058 118572 502064 118584
rect 502019 118544 502064 118572
rect 502058 118532 502064 118544
rect 502116 118532 502122 118584
rect 83274 118464 83280 118516
rect 83332 118504 83338 118516
rect 267734 118504 267740 118516
rect 83332 118476 267740 118504
rect 83332 118464 83338 118476
rect 267734 118464 267740 118476
rect 267792 118464 267798 118516
rect 81802 118396 81808 118448
rect 81860 118436 81866 118448
rect 269114 118436 269120 118448
rect 81860 118408 269120 118436
rect 81860 118396 81866 118408
rect 269114 118396 269120 118408
rect 269172 118396 269178 118448
rect 83090 118328 83096 118380
rect 83148 118368 83154 118380
rect 287054 118368 287060 118380
rect 83148 118340 287060 118368
rect 83148 118328 83154 118340
rect 287054 118328 287060 118340
rect 287112 118328 287118 118380
rect 500218 118328 500224 118380
rect 500276 118368 500282 118380
rect 504542 118368 504548 118380
rect 500276 118340 504548 118368
rect 500276 118328 500282 118340
rect 504542 118328 504548 118340
rect 504600 118328 504606 118380
rect 80514 118260 80520 118312
rect 80572 118300 80578 118312
rect 304994 118300 305000 118312
rect 80572 118272 305000 118300
rect 80572 118260 80578 118272
rect 304994 118260 305000 118272
rect 305052 118260 305058 118312
rect 413554 118260 413560 118312
rect 413612 118300 413618 118312
rect 413922 118300 413928 118312
rect 413612 118272 413928 118300
rect 413612 118260 413618 118272
rect 413922 118260 413928 118272
rect 413980 118260 413986 118312
rect 422202 118260 422208 118312
rect 422260 118300 422266 118312
rect 503530 118300 503536 118312
rect 422260 118272 503536 118300
rect 422260 118260 422266 118272
rect 503530 118260 503536 118272
rect 503588 118260 503594 118312
rect 78950 118192 78956 118244
rect 79008 118232 79014 118244
rect 320174 118232 320180 118244
rect 79008 118204 320180 118232
rect 79008 118192 79014 118204
rect 320174 118192 320180 118204
rect 320232 118192 320238 118244
rect 398742 118192 398748 118244
rect 398800 118232 398806 118244
rect 503254 118232 503260 118244
rect 398800 118204 503260 118232
rect 398800 118192 398806 118204
rect 503254 118192 503260 118204
rect 503312 118192 503318 118244
rect 82538 118124 82544 118176
rect 82596 118164 82602 118176
rect 84838 118164 84844 118176
rect 82596 118136 84844 118164
rect 82596 118124 82602 118136
rect 84838 118124 84844 118136
rect 84896 118124 84902 118176
rect 244366 118164 244372 118176
rect 86236 118136 244372 118164
rect 82170 118056 82176 118108
rect 82228 118096 82234 118108
rect 86236 118096 86264 118136
rect 244366 118124 244372 118136
rect 244424 118124 244430 118176
rect 249702 118124 249708 118176
rect 249760 118164 249766 118176
rect 503346 118164 503352 118176
rect 249760 118136 503352 118164
rect 249760 118124 249766 118136
rect 503346 118124 503352 118136
rect 503404 118124 503410 118176
rect 82228 118068 86264 118096
rect 86313 118099 86371 118105
rect 82228 118056 82234 118068
rect 86313 118065 86325 118099
rect 86359 118096 86371 118099
rect 132586 118096 132592 118108
rect 86359 118068 132592 118096
rect 86359 118065 86371 118068
rect 86313 118059 86371 118065
rect 132586 118056 132592 118068
rect 132644 118056 132650 118108
rect 220722 118056 220728 118108
rect 220780 118096 220786 118108
rect 504266 118096 504272 118108
rect 220780 118068 504272 118096
rect 220780 118056 220786 118068
rect 504266 118056 504272 118068
rect 504324 118056 504330 118108
rect 81986 117988 81992 118040
rect 82044 118028 82050 118040
rect 514754 118028 514760 118040
rect 82044 118000 514760 118028
rect 82044 117988 82050 118000
rect 514754 117988 514760 118000
rect 514812 117988 514818 118040
rect 82078 117920 82084 117972
rect 82136 117960 82142 117972
rect 536926 117960 536932 117972
rect 82136 117932 536932 117960
rect 82136 117920 82142 117932
rect 536926 117920 536932 117932
rect 536984 117920 536990 117972
rect 500126 117784 500132 117836
rect 500184 117824 500190 117836
rect 503441 117827 503499 117833
rect 503441 117824 503453 117827
rect 500184 117796 503453 117824
rect 500184 117784 500190 117796
rect 503441 117793 503453 117796
rect 503487 117793 503499 117827
rect 503441 117787 503499 117793
rect 492306 117308 492312 117360
rect 492364 117348 492370 117360
rect 496722 117348 496728 117360
rect 492364 117320 496728 117348
rect 492364 117308 492370 117320
rect 496722 117308 496728 117320
rect 496780 117308 496786 117360
rect 490558 117104 490564 117156
rect 490616 117144 490622 117156
rect 493502 117144 493508 117156
rect 490616 117116 493508 117144
rect 490616 117104 490622 117116
rect 493502 117104 493508 117116
rect 493560 117104 493566 117156
rect 82446 116764 82452 116816
rect 82504 116804 82510 116816
rect 161474 116804 161480 116816
rect 82504 116776 161480 116804
rect 82504 116764 82510 116776
rect 161474 116764 161480 116776
rect 161532 116764 161538 116816
rect 322750 116764 322756 116816
rect 322808 116804 322814 116816
rect 511166 116804 511172 116816
rect 322808 116776 511172 116804
rect 322808 116764 322814 116776
rect 511166 116764 511172 116776
rect 511224 116764 511230 116816
rect 83826 116696 83832 116748
rect 83884 116736 83890 116748
rect 372522 116736 372528 116748
rect 83884 116708 372528 116736
rect 83884 116696 83890 116708
rect 372522 116696 372528 116708
rect 372580 116696 372586 116748
rect 401502 116696 401508 116748
rect 401560 116736 401566 116748
rect 502978 116736 502984 116748
rect 401560 116708 502984 116736
rect 401560 116696 401566 116708
rect 502978 116696 502984 116708
rect 503036 116696 503042 116748
rect 136542 116628 136548 116680
rect 136600 116668 136606 116680
rect 505002 116668 505008 116680
rect 136600 116640 505008 116668
rect 136600 116628 136606 116640
rect 505002 116628 505008 116640
rect 505060 116628 505066 116680
rect 79134 116560 79140 116612
rect 79192 116600 79198 116612
rect 451274 116600 451280 116612
rect 79192 116572 451280 116600
rect 79192 116560 79198 116572
rect 451274 116560 451280 116572
rect 451332 116560 451338 116612
rect 415486 116084 415492 116136
rect 415544 116124 415550 116136
rect 415946 116124 415952 116136
rect 415544 116096 415952 116124
rect 415544 116084 415550 116096
rect 415946 116084 415952 116096
rect 416004 116084 416010 116136
rect 161290 116056 161296 116068
rect 161251 116028 161296 116056
rect 161290 116016 161296 116028
rect 161348 116016 161354 116068
rect 153010 115948 153016 116000
rect 153068 115988 153074 116000
rect 153102 115988 153108 116000
rect 153068 115960 153108 115988
rect 153068 115948 153074 115960
rect 153102 115948 153108 115960
rect 153160 115948 153166 116000
rect 509602 115948 509608 116000
rect 509660 115988 509666 116000
rect 511442 115988 511448 116000
rect 509660 115960 511448 115988
rect 509660 115948 509666 115960
rect 511442 115948 511448 115960
rect 511500 115948 511506 116000
rect 131206 115920 131212 115932
rect 131167 115892 131212 115920
rect 131206 115880 131212 115892
rect 131264 115880 131270 115932
rect 155862 115880 155868 115932
rect 155920 115920 155926 115932
rect 156138 115920 156144 115932
rect 155920 115892 156144 115920
rect 155920 115880 155926 115892
rect 156138 115880 156144 115892
rect 156196 115880 156202 115932
rect 161290 115920 161296 115932
rect 161251 115892 161296 115920
rect 161290 115880 161296 115892
rect 161348 115880 161354 115932
rect 179322 115920 179328 115932
rect 179283 115892 179328 115920
rect 179322 115880 179328 115892
rect 179380 115880 179386 115932
rect 244274 115920 244280 115932
rect 244235 115892 244280 115920
rect 244274 115880 244280 115892
rect 244332 115880 244338 115932
rect 258074 115920 258080 115932
rect 258035 115892 258080 115920
rect 258074 115880 258080 115892
rect 258132 115880 258138 115932
rect 445846 115920 445852 115932
rect 445807 115892 445852 115920
rect 445846 115880 445852 115892
rect 445904 115880 445910 115932
rect 153010 115852 153016 115864
rect 152971 115824 153016 115852
rect 153010 115812 153016 115824
rect 153068 115812 153074 115864
rect 511626 115852 511632 115864
rect 511587 115824 511632 115852
rect 511626 115812 511632 115824
rect 511684 115812 511690 115864
rect 278682 115404 278688 115456
rect 278740 115444 278746 115456
rect 502702 115444 502708 115456
rect 278740 115416 502708 115444
rect 278740 115404 278746 115416
rect 502702 115404 502708 115416
rect 502760 115404 502766 115456
rect 186225 115379 186283 115385
rect 186225 115345 186237 115379
rect 186271 115376 186283 115379
rect 504910 115376 504916 115388
rect 186271 115348 504916 115376
rect 186271 115345 186283 115348
rect 186225 115339 186283 115345
rect 504910 115336 504916 115348
rect 504968 115336 504974 115388
rect 183462 115268 183468 115320
rect 183520 115308 183526 115320
rect 504634 115308 504640 115320
rect 183520 115280 504640 115308
rect 183520 115268 183526 115280
rect 504634 115268 504640 115280
rect 504692 115268 504698 115320
rect 80330 115200 80336 115252
rect 80388 115240 80394 115252
rect 552014 115240 552020 115252
rect 80388 115212 552020 115240
rect 80388 115200 80394 115212
rect 552014 115200 552020 115212
rect 552072 115200 552078 115252
rect 393314 115132 393320 115184
rect 393372 115172 393378 115184
rect 394602 115172 394608 115184
rect 393372 115144 394608 115172
rect 393372 115132 393378 115144
rect 394602 115132 394608 115144
rect 394660 115132 394666 115184
rect 500310 114656 500316 114708
rect 500368 114696 500374 114708
rect 507302 114696 507308 114708
rect 500368 114668 507308 114696
rect 500368 114656 500374 114668
rect 507302 114656 507308 114668
rect 507360 114656 507366 114708
rect 110414 114560 110420 114572
rect 110375 114532 110420 114560
rect 110414 114520 110420 114532
rect 110472 114520 110478 114572
rect 186222 114560 186228 114572
rect 186183 114532 186228 114560
rect 186222 114520 186228 114532
rect 186280 114520 186286 114572
rect 272978 114520 272984 114572
rect 273036 114560 273042 114572
rect 273070 114560 273076 114572
rect 273036 114532 273076 114560
rect 273036 114520 273042 114532
rect 273070 114520 273076 114532
rect 273128 114520 273134 114572
rect 524414 114560 524420 114572
rect 524375 114532 524420 114560
rect 524414 114520 524420 114532
rect 524472 114520 524478 114572
rect 532694 114560 532700 114572
rect 532655 114532 532700 114560
rect 532694 114520 532700 114532
rect 532752 114520 532758 114572
rect 155862 114492 155868 114504
rect 155823 114464 155868 114492
rect 155862 114452 155868 114464
rect 155920 114452 155926 114504
rect 511537 114495 511595 114501
rect 511537 114461 511549 114495
rect 511583 114492 511595 114495
rect 511626 114492 511632 114504
rect 511583 114464 511632 114492
rect 511583 114461 511595 114464
rect 511537 114455 511595 114461
rect 511626 114452 511632 114464
rect 511684 114452 511690 114504
rect 110414 114424 110420 114436
rect 110375 114396 110420 114424
rect 110414 114384 110420 114396
rect 110472 114384 110478 114436
rect 487522 114112 487528 114164
rect 487580 114152 487586 114164
rect 492306 114152 492312 114164
rect 487580 114124 492312 114152
rect 487580 114112 487586 114124
rect 492306 114112 492312 114124
rect 492364 114112 492370 114164
rect 348970 113840 348976 113892
rect 349028 113880 349034 113892
rect 502334 113880 502340 113892
rect 349028 113852 502340 113880
rect 349028 113840 349034 113852
rect 502334 113840 502340 113852
rect 502392 113840 502398 113892
rect 79226 113772 79232 113824
rect 79284 113812 79290 113824
rect 454034 113812 454040 113824
rect 79284 113784 454040 113812
rect 79284 113772 79290 113784
rect 454034 113772 454040 113784
rect 454092 113772 454098 113824
rect 82722 113200 82728 113212
rect 82683 113172 82728 113200
rect 82722 113160 82728 113172
rect 82780 113160 82786 113212
rect 505830 113160 505836 113212
rect 505888 113200 505894 113212
rect 506290 113200 506296 113212
rect 505888 113172 506296 113200
rect 505888 113160 505894 113172
rect 506290 113160 506296 113172
rect 506348 113160 506354 113212
rect 89530 113092 89536 113144
rect 89588 113092 89594 113144
rect 89548 113064 89576 113092
rect 89622 113064 89628 113076
rect 89548 113036 89628 113064
rect 89622 113024 89628 113036
rect 89680 113024 89686 113076
rect 110322 112412 110328 112464
rect 110380 112452 110386 112464
rect 505922 112452 505928 112464
rect 110380 112424 505928 112452
rect 110380 112412 110386 112424
rect 505922 112412 505928 112424
rect 505980 112412 505986 112464
rect 481726 111800 481732 111852
rect 481784 111840 481790 111852
rect 487522 111840 487528 111852
rect 481784 111812 487528 111840
rect 481784 111800 481790 111812
rect 487522 111800 487528 111812
rect 487580 111800 487586 111852
rect 506934 111800 506940 111852
rect 506992 111840 506998 111852
rect 509602 111840 509608 111852
rect 506992 111812 509608 111840
rect 506992 111800 506998 111812
rect 509602 111800 509608 111812
rect 509660 111800 509666 111852
rect 80054 111772 80060 111784
rect 80015 111744 80060 111772
rect 80054 111732 80060 111744
rect 80112 111732 80118 111784
rect 82630 111732 82636 111784
rect 82688 111772 82694 111784
rect 82722 111772 82728 111784
rect 82688 111744 82728 111772
rect 82688 111732 82694 111744
rect 82722 111732 82728 111744
rect 82780 111732 82786 111784
rect 83366 111732 83372 111784
rect 83424 111732 83430 111784
rect 83734 111732 83740 111784
rect 83792 111772 83798 111784
rect 83826 111772 83832 111784
rect 83792 111744 83832 111772
rect 83792 111732 83798 111744
rect 83826 111732 83832 111744
rect 83884 111732 83890 111784
rect 83384 111704 83412 111732
rect 83458 111704 83464 111716
rect 83384 111676 83464 111704
rect 83458 111664 83464 111676
rect 83516 111664 83522 111716
rect 508130 111392 508136 111444
rect 508188 111432 508194 111444
rect 509878 111432 509884 111444
rect 508188 111404 509884 111432
rect 508188 111392 508194 111404
rect 509878 111392 509884 111404
rect 509936 111392 509942 111444
rect 304902 111296 304908 111308
rect 304863 111268 304908 111296
rect 304902 111256 304908 111268
rect 304960 111256 304966 111308
rect 440142 111256 440148 111308
rect 440200 111256 440206 111308
rect 295334 111188 295340 111240
rect 295392 111228 295398 111240
rect 304810 111228 304816 111240
rect 295392 111200 304816 111228
rect 295392 111188 295398 111200
rect 304810 111188 304816 111200
rect 304868 111188 304874 111240
rect 372706 111188 372712 111240
rect 372764 111228 372770 111240
rect 382090 111228 382096 111240
rect 372764 111200 382096 111228
rect 372764 111188 372770 111200
rect 382090 111188 382096 111200
rect 382148 111188 382154 111240
rect 411254 111188 411260 111240
rect 411312 111228 411318 111240
rect 420730 111228 420736 111240
rect 411312 111200 420736 111228
rect 411312 111188 411318 111200
rect 420730 111188 420736 111200
rect 420788 111188 420794 111240
rect 81066 111120 81072 111172
rect 81124 111160 81130 111172
rect 263594 111160 263600 111172
rect 81124 111132 263600 111160
rect 81124 111120 81130 111132
rect 263594 111120 263600 111132
rect 263652 111120 263658 111172
rect 276014 111120 276020 111172
rect 276072 111160 276078 111172
rect 285490 111160 285496 111172
rect 276072 111132 285496 111160
rect 276072 111120 276078 111132
rect 285490 111120 285496 111132
rect 285548 111120 285554 111172
rect 314654 111120 314660 111172
rect 314712 111160 314718 111172
rect 323578 111160 323584 111172
rect 314712 111132 323584 111160
rect 314712 111120 314718 111132
rect 323578 111120 323584 111132
rect 323636 111120 323642 111172
rect 353294 111120 353300 111172
rect 353352 111160 353358 111172
rect 362770 111160 362776 111172
rect 353352 111132 362776 111160
rect 353352 111120 353358 111132
rect 362770 111120 362776 111132
rect 362828 111120 362834 111172
rect 430574 111120 430580 111172
rect 430632 111160 430638 111172
rect 440050 111160 440056 111172
rect 430632 111132 440056 111160
rect 430632 111120 430638 111132
rect 440050 111120 440056 111132
rect 440108 111120 440114 111172
rect 440160 111104 440188 111256
rect 79318 111052 79324 111104
rect 79376 111092 79382 111104
rect 436097 111095 436155 111101
rect 436097 111092 436109 111095
rect 79376 111064 436109 111092
rect 79376 111052 79382 111064
rect 436097 111061 436109 111064
rect 436143 111061 436155 111095
rect 436097 111055 436155 111061
rect 440142 111052 440148 111104
rect 440200 111052 440206 111104
rect 378134 111024 378140 111036
rect 378095 110996 378140 111024
rect 378134 110984 378140 110996
rect 378192 110984 378198 111036
rect 117501 110415 117559 110421
rect 117501 110381 117513 110415
rect 117547 110412 117559 110415
rect 117682 110412 117688 110424
rect 117547 110384 117688 110412
rect 117547 110381 117559 110384
rect 117501 110375 117559 110381
rect 117682 110372 117688 110384
rect 117740 110372 117746 110424
rect 505830 109828 505836 109880
rect 505888 109868 505894 109880
rect 506106 109868 506112 109880
rect 505888 109840 506112 109868
rect 505888 109828 505894 109840
rect 506106 109828 506112 109840
rect 506164 109828 506170 109880
rect 481358 109760 481364 109812
rect 481416 109800 481422 109812
rect 481726 109800 481732 109812
rect 481416 109772 481732 109800
rect 481416 109760 481422 109772
rect 481726 109760 481732 109772
rect 481784 109760 481790 109812
rect 85482 109692 85488 109744
rect 85540 109732 85546 109744
rect 505646 109732 505652 109744
rect 85540 109704 505652 109732
rect 85540 109692 85546 109704
rect 505646 109692 505652 109704
rect 505704 109692 505710 109744
rect 272889 109191 272947 109197
rect 272889 109157 272901 109191
rect 272935 109188 272947 109191
rect 272978 109188 272984 109200
rect 272935 109160 272984 109188
rect 272935 109157 272947 109160
rect 272889 109151 272947 109157
rect 272978 109148 272984 109160
rect 273036 109148 273042 109200
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 508958 108984 508964 108996
rect 3292 108956 508964 108984
rect 3292 108944 3298 108956
rect 508958 108944 508964 108956
rect 509016 108944 509022 108996
rect 121362 108876 121368 108928
rect 121420 108916 121426 108928
rect 121546 108916 121552 108928
rect 121420 108888 121552 108916
rect 121420 108876 121426 108888
rect 121546 108876 121552 108888
rect 121604 108876 121610 108928
rect 153010 108916 153016 108928
rect 152971 108888 153016 108916
rect 153010 108876 153016 108888
rect 153068 108876 153074 108928
rect 161290 108916 161296 108928
rect 161251 108888 161296 108916
rect 161290 108876 161296 108888
rect 161348 108876 161354 108928
rect 272886 108916 272892 108928
rect 272847 108888 272892 108916
rect 272886 108876 272892 108888
rect 272944 108876 272950 108928
rect 479610 107448 479616 107500
rect 479668 107488 479674 107500
rect 481358 107488 481364 107500
rect 479668 107460 481364 107488
rect 479668 107448 479674 107460
rect 481358 107448 481364 107460
rect 481416 107448 481422 107500
rect 179322 106400 179328 106412
rect 179283 106372 179328 106400
rect 179322 106360 179328 106372
rect 179380 106360 179386 106412
rect 131206 106332 131212 106344
rect 131167 106304 131212 106332
rect 131206 106292 131212 106304
rect 131264 106292 131270 106344
rect 244274 106332 244280 106344
rect 244235 106304 244280 106332
rect 244274 106292 244280 106304
rect 244332 106292 244338 106344
rect 445846 106332 445852 106344
rect 445807 106304 445852 106332
rect 445846 106292 445852 106304
rect 445904 106292 445910 106344
rect 505738 106292 505744 106344
rect 505796 106332 505802 106344
rect 508130 106332 508136 106344
rect 505796 106304 508136 106332
rect 505796 106292 505802 106304
rect 508130 106292 508136 106304
rect 508188 106292 508194 106344
rect 304902 105516 304908 105528
rect 304863 105488 304908 105516
rect 304902 105476 304908 105488
rect 304960 105476 304966 105528
rect 351730 104932 351736 104984
rect 351788 104972 351794 104984
rect 351914 104972 351920 104984
rect 351788 104944 351920 104972
rect 351788 104932 351794 104944
rect 351914 104932 351920 104944
rect 351972 104932 351978 104984
rect 110414 104904 110420 104916
rect 110375 104876 110420 104904
rect 110414 104864 110420 104876
rect 110472 104864 110478 104916
rect 155865 104907 155923 104913
rect 155865 104873 155877 104907
rect 155911 104904 155923 104907
rect 156046 104904 156052 104916
rect 155911 104876 156052 104904
rect 155911 104873 155923 104876
rect 155865 104867 155923 104873
rect 156046 104864 156052 104876
rect 156104 104864 156110 104916
rect 511534 104904 511540 104916
rect 511495 104876 511540 104904
rect 511534 104864 511540 104876
rect 511592 104864 511598 104916
rect 179322 104836 179328 104848
rect 179283 104808 179328 104836
rect 179322 104796 179328 104808
rect 179380 104796 179386 104848
rect 186222 104836 186228 104848
rect 186183 104808 186228 104836
rect 186222 104796 186228 104808
rect 186280 104796 186286 104848
rect 220722 104836 220728 104848
rect 220683 104808 220728 104836
rect 220722 104796 220728 104808
rect 220780 104796 220786 104848
rect 223574 104836 223580 104848
rect 223535 104808 223580 104836
rect 223574 104796 223580 104808
rect 223632 104796 223638 104848
rect 351730 104836 351736 104848
rect 351691 104808 351736 104836
rect 351730 104796 351736 104808
rect 351788 104796 351794 104848
rect 524414 104836 524420 104848
rect 524375 104808 524420 104836
rect 524414 104796 524420 104808
rect 524472 104796 524478 104848
rect 532694 104836 532700 104848
rect 532655 104808 532700 104836
rect 532694 104796 532700 104808
rect 532752 104796 532758 104848
rect 156138 104728 156144 104780
rect 156196 104768 156202 104780
rect 156233 104771 156291 104777
rect 156233 104768 156245 104771
rect 156196 104740 156245 104768
rect 156196 104728 156202 104740
rect 156233 104737 156245 104740
rect 156279 104737 156291 104771
rect 156233 104731 156291 104737
rect 511626 104728 511632 104780
rect 511684 104768 511690 104780
rect 511721 104771 511779 104777
rect 511721 104768 511733 104771
rect 511684 104740 511733 104768
rect 511684 104728 511690 104740
rect 511721 104737 511733 104740
rect 511767 104737 511779 104771
rect 511721 104731 511779 104737
rect 489178 103096 489184 103148
rect 489236 103136 489242 103148
rect 490558 103136 490564 103148
rect 489236 103108 490564 103136
rect 489236 103096 489242 103108
rect 490558 103096 490564 103108
rect 490616 103096 490622 103148
rect 258074 102932 258080 102944
rect 258035 102904 258080 102932
rect 258074 102892 258080 102904
rect 258132 102892 258138 102944
rect 80054 102184 80060 102196
rect 80015 102156 80060 102184
rect 80054 102144 80060 102156
rect 80112 102144 80118 102196
rect 266078 102144 266084 102196
rect 266136 102184 266142 102196
rect 266262 102184 266268 102196
rect 266136 102156 266268 102184
rect 266136 102144 266142 102156
rect 266262 102144 266268 102156
rect 266320 102144 266326 102196
rect 506934 102184 506940 102196
rect 502352 102156 506940 102184
rect 501230 102076 501236 102128
rect 501288 102116 501294 102128
rect 502352 102116 502380 102156
rect 506934 102144 506940 102156
rect 506992 102144 506998 102196
rect 501288 102088 502380 102116
rect 501288 102076 501294 102088
rect 117498 100824 117504 100836
rect 117459 100796 117504 100824
rect 117498 100784 117504 100796
rect 117556 100784 117562 100836
rect 117498 100648 117504 100700
rect 117556 100688 117562 100700
rect 117774 100688 117780 100700
rect 117556 100660 117780 100688
rect 117556 100648 117562 100660
rect 117774 100648 117780 100660
rect 117832 100648 117838 100700
rect 497458 99832 497464 99884
rect 497516 99872 497522 99884
rect 500310 99872 500316 99884
rect 497516 99844 500316 99872
rect 497516 99832 497522 99844
rect 500310 99832 500316 99844
rect 500368 99832 500374 99884
rect 299290 99424 299296 99476
rect 299348 99424 299354 99476
rect 121454 99356 121460 99408
rect 121512 99396 121518 99408
rect 121638 99396 121644 99408
rect 121512 99368 121644 99396
rect 121512 99356 121518 99368
rect 121638 99356 121644 99368
rect 121696 99356 121702 99408
rect 161198 99356 161204 99408
rect 161256 99396 161262 99408
rect 161382 99396 161388 99408
rect 161256 99368 161388 99396
rect 161256 99356 161262 99368
rect 161382 99356 161388 99368
rect 161440 99356 161446 99408
rect 299308 99340 299336 99424
rect 79686 99288 79692 99340
rect 79744 99328 79750 99340
rect 79962 99328 79968 99340
rect 79744 99300 79968 99328
rect 79744 99288 79750 99300
rect 79962 99288 79968 99300
rect 80020 99288 80026 99340
rect 117501 99331 117559 99337
rect 117501 99297 117513 99331
rect 117547 99328 117559 99331
rect 117774 99328 117780 99340
rect 117547 99300 117780 99328
rect 117547 99297 117559 99300
rect 117501 99291 117559 99297
rect 117774 99288 117780 99300
rect 117832 99288 117838 99340
rect 299290 99288 299296 99340
rect 299348 99288 299354 99340
rect 272610 99220 272616 99272
rect 272668 99260 272674 99272
rect 272978 99260 272984 99272
rect 272668 99232 272984 99260
rect 272668 99220 272674 99232
rect 272978 99220 272984 99232
rect 273036 99220 273042 99272
rect 475378 98404 475384 98456
rect 475436 98444 475442 98456
rect 479610 98444 479616 98456
rect 475436 98416 479616 98444
rect 475436 98404 475442 98416
rect 479610 98404 479616 98416
rect 479668 98404 479674 98456
rect 500310 97996 500316 98048
rect 500368 98036 500374 98048
rect 501230 98036 501236 98048
rect 500368 98008 501236 98036
rect 500368 97996 500374 98008
rect 501230 97996 501236 98008
rect 501288 97996 501294 98048
rect 436094 96744 436100 96756
rect 436055 96716 436100 96744
rect 436094 96704 436100 96716
rect 436152 96704 436158 96756
rect 131206 96608 131212 96620
rect 131167 96580 131212 96608
rect 131206 96568 131212 96580
rect 131264 96568 131270 96620
rect 161198 96568 161204 96620
rect 161256 96608 161262 96620
rect 161290 96608 161296 96620
rect 161256 96580 161296 96608
rect 161256 96568 161262 96580
rect 161290 96568 161296 96580
rect 161348 96568 161354 96620
rect 244274 96608 244280 96620
rect 244235 96580 244280 96608
rect 244274 96568 244280 96580
rect 244332 96568 244338 96620
rect 258074 96608 258080 96620
rect 258035 96580 258080 96608
rect 258074 96568 258080 96580
rect 258132 96568 258138 96620
rect 272978 96608 272984 96620
rect 272939 96580 272984 96608
rect 272978 96568 272984 96580
rect 273036 96568 273042 96620
rect 289538 96568 289544 96620
rect 289596 96608 289602 96620
rect 289722 96608 289728 96620
rect 289596 96580 289728 96608
rect 289596 96568 289602 96580
rect 289722 96568 289728 96580
rect 289780 96568 289786 96620
rect 299290 96608 299296 96620
rect 299251 96580 299296 96608
rect 299290 96568 299296 96580
rect 299348 96568 299354 96620
rect 436094 96568 436100 96620
rect 436152 96608 436158 96620
rect 436278 96608 436284 96620
rect 436152 96580 436284 96608
rect 436152 96568 436158 96580
rect 436278 96568 436284 96580
rect 436336 96568 436342 96620
rect 445846 96608 445852 96620
rect 445807 96580 445852 96608
rect 445846 96568 445852 96580
rect 445904 96568 445910 96620
rect 511718 96540 511724 96552
rect 511679 96512 511724 96540
rect 511718 96500 511724 96512
rect 511776 96500 511782 96552
rect 120258 95276 120264 95328
rect 120316 95316 120322 95328
rect 120350 95316 120356 95328
rect 120316 95288 120356 95316
rect 120316 95276 120322 95288
rect 120350 95276 120356 95288
rect 120408 95276 120414 95328
rect 152918 95208 152924 95260
rect 152976 95248 152982 95260
rect 153102 95248 153108 95260
rect 152976 95220 153108 95248
rect 152976 95208 152982 95220
rect 153102 95208 153108 95220
rect 153160 95208 153166 95260
rect 156230 95248 156236 95260
rect 156191 95220 156236 95248
rect 156230 95208 156236 95220
rect 156288 95208 156294 95260
rect 186222 95248 186228 95260
rect 186183 95220 186228 95248
rect 186222 95208 186228 95220
rect 186280 95208 186286 95260
rect 220722 95248 220728 95260
rect 220683 95220 220728 95248
rect 220722 95208 220728 95220
rect 220780 95208 220786 95260
rect 223574 95248 223580 95260
rect 223535 95220 223580 95248
rect 223574 95208 223580 95220
rect 223632 95208 223638 95260
rect 378134 95248 378140 95260
rect 378095 95220 378140 95248
rect 378134 95208 378140 95220
rect 378192 95208 378198 95260
rect 524414 95248 524420 95260
rect 524375 95220 524420 95248
rect 524414 95208 524420 95220
rect 524472 95208 524478 95260
rect 532694 95248 532700 95260
rect 532655 95220 532700 95248
rect 532694 95208 532700 95220
rect 532752 95208 532758 95260
rect 110414 95180 110420 95192
rect 110375 95152 110420 95180
rect 110414 95140 110420 95152
rect 110472 95140 110478 95192
rect 220538 95180 220544 95192
rect 220499 95152 220544 95180
rect 220538 95140 220544 95152
rect 220596 95140 220602 95192
rect 500218 93888 500224 93900
rect 500179 93860 500224 93888
rect 500218 93848 500224 93860
rect 500276 93848 500282 93900
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 33870 93820 33876 93832
rect 3476 93792 33876 93820
rect 3476 93780 3482 93792
rect 33870 93780 33876 93792
rect 33928 93780 33934 93832
rect 120258 92420 120264 92472
rect 120316 92460 120322 92472
rect 120350 92460 120356 92472
rect 120316 92432 120356 92460
rect 120316 92420 120322 92432
rect 120350 92420 120356 92432
rect 120408 92420 120414 92472
rect 473998 91060 474004 91112
rect 474056 91100 474062 91112
rect 475378 91100 475384 91112
rect 474056 91072 475384 91100
rect 474056 91060 474062 91072
rect 475378 91060 475384 91072
rect 475436 91060 475442 91112
rect 79318 90992 79324 91044
rect 79376 91032 79382 91044
rect 79962 91032 79968 91044
rect 79376 91004 79968 91032
rect 79376 90992 79382 91004
rect 79962 90992 79968 91004
rect 80020 90992 80026 91044
rect 117498 89740 117504 89752
rect 117459 89712 117504 89740
rect 117498 89700 117504 89712
rect 117556 89700 117562 89752
rect 121454 89700 121460 89752
rect 121512 89740 121518 89752
rect 121638 89740 121644 89752
rect 121512 89712 121644 89740
rect 121512 89700 121518 89712
rect 121638 89700 121644 89712
rect 121696 89700 121702 89752
rect 351730 89672 351736 89684
rect 351691 89644 351736 89672
rect 351730 89632 351736 89644
rect 351788 89632 351794 89684
rect 179322 87088 179328 87100
rect 179283 87060 179328 87088
rect 179322 87048 179328 87060
rect 179380 87048 179386 87100
rect 131206 87020 131212 87032
rect 131167 86992 131212 87020
rect 131206 86980 131212 86992
rect 131264 86980 131270 87032
rect 244274 87020 244280 87032
rect 244235 86992 244280 87020
rect 244274 86980 244280 86992
rect 244332 86980 244338 87032
rect 258074 87020 258080 87032
rect 258035 86992 258080 87020
rect 258074 86980 258080 86992
rect 258132 86980 258138 87032
rect 272978 87020 272984 87032
rect 272939 86992 272984 87020
rect 272978 86980 272984 86992
rect 273036 86980 273042 87032
rect 299290 87020 299296 87032
rect 299251 86992 299296 87020
rect 299290 86980 299296 86992
rect 299348 86980 299354 87032
rect 445846 87020 445852 87032
rect 445807 86992 445852 87020
rect 445846 86980 445852 86992
rect 445904 86980 445910 87032
rect 511626 86980 511632 87032
rect 511684 87020 511690 87032
rect 511718 87020 511724 87032
rect 511684 86992 511724 87020
rect 511684 86980 511690 86992
rect 511718 86980 511724 86992
rect 511776 86980 511782 87032
rect 436094 86952 436100 86964
rect 436055 86924 436100 86952
rect 436094 86912 436100 86924
rect 436152 86912 436158 86964
rect 487154 86708 487160 86760
rect 487212 86748 487218 86760
rect 489178 86748 489184 86760
rect 487212 86720 489184 86748
rect 487212 86708 487218 86720
rect 489178 86708 489184 86720
rect 489236 86708 489242 86760
rect 135070 86232 135076 86284
rect 135128 86272 135134 86284
rect 504450 86272 504456 86284
rect 135128 86244 504456 86272
rect 135128 86232 135134 86244
rect 504450 86232 504456 86244
rect 504508 86232 504514 86284
rect 110414 85660 110420 85672
rect 110375 85632 110420 85660
rect 110414 85620 110420 85632
rect 110472 85620 110478 85672
rect 161014 85552 161020 85604
rect 161072 85592 161078 85604
rect 161290 85592 161296 85604
rect 161072 85564 161296 85592
rect 161072 85552 161078 85564
rect 161290 85552 161296 85564
rect 161348 85552 161354 85604
rect 220538 85592 220544 85604
rect 220499 85564 220544 85592
rect 220538 85552 220544 85564
rect 220596 85552 220602 85604
rect 110414 85484 110420 85536
rect 110472 85524 110478 85536
rect 110506 85524 110512 85536
rect 110472 85496 110512 85524
rect 110472 85484 110478 85496
rect 110506 85484 110512 85496
rect 110564 85484 110570 85536
rect 179322 85524 179328 85536
rect 179283 85496 179328 85524
rect 179322 85484 179328 85496
rect 179380 85484 179386 85536
rect 186222 85524 186228 85536
rect 186183 85496 186228 85524
rect 186222 85484 186228 85496
rect 186280 85484 186286 85536
rect 220633 85527 220691 85533
rect 220633 85493 220645 85527
rect 220679 85524 220691 85527
rect 220722 85524 220728 85536
rect 220679 85496 220728 85524
rect 220679 85493 220691 85496
rect 220633 85487 220691 85493
rect 220722 85484 220728 85496
rect 220780 85484 220786 85536
rect 223574 85524 223580 85536
rect 223535 85496 223580 85524
rect 223574 85484 223580 85496
rect 223632 85484 223638 85536
rect 378134 85524 378140 85536
rect 378095 85496 378140 85524
rect 378134 85484 378140 85496
rect 378192 85484 378198 85536
rect 511534 85524 511540 85536
rect 511495 85496 511540 85524
rect 511534 85484 511540 85496
rect 511592 85484 511598 85536
rect 524414 85524 524420 85536
rect 524375 85496 524420 85524
rect 524414 85484 524420 85496
rect 524472 85484 524478 85536
rect 532694 85524 532700 85536
rect 532655 85496 532700 85524
rect 532694 85484 532700 85496
rect 532752 85484 532758 85536
rect 497550 84464 497556 84516
rect 497608 84504 497614 84516
rect 500310 84504 500316 84516
rect 497608 84476 500316 84504
rect 497608 84464 497614 84476
rect 500310 84464 500316 84476
rect 500368 84464 500374 84516
rect 80238 83444 80244 83496
rect 80296 83484 80302 83496
rect 444466 83484 444472 83496
rect 80296 83456 444472 83484
rect 80296 83444 80302 83456
rect 444466 83444 444472 83456
rect 444524 83444 444530 83496
rect 120350 82872 120356 82884
rect 120311 82844 120356 82872
rect 120350 82832 120356 82844
rect 120408 82832 120414 82884
rect 80054 82804 80060 82816
rect 80015 82776 80060 82804
rect 80054 82764 80060 82776
rect 80112 82764 80118 82816
rect 210970 82084 210976 82136
rect 211028 82124 211034 82136
rect 504726 82124 504732 82136
rect 211028 82096 504732 82124
rect 211028 82084 211034 82096
rect 504726 82084 504732 82096
rect 504784 82084 504790 82136
rect 79318 81880 79324 81932
rect 79376 81920 79382 81932
rect 79962 81920 79968 81932
rect 79376 81892 79968 81920
rect 79376 81880 79382 81892
rect 79962 81880 79968 81892
rect 80020 81880 80026 81932
rect 117498 81404 117504 81456
rect 117556 81444 117562 81456
rect 117590 81444 117596 81456
rect 117556 81416 117596 81444
rect 117556 81404 117562 81416
rect 117590 81404 117596 81416
rect 117648 81404 117654 81456
rect 120350 81444 120356 81456
rect 120311 81416 120356 81444
rect 120350 81404 120356 81416
rect 120408 81404 120414 81456
rect 472342 81404 472348 81456
rect 472400 81444 472406 81456
rect 473998 81444 474004 81456
rect 472400 81416 474004 81444
rect 472400 81404 472406 81416
rect 473998 81404 474004 81416
rect 474056 81404 474062 81456
rect 486142 81404 486148 81456
rect 486200 81444 486206 81456
rect 487154 81444 487160 81456
rect 486200 81416 487160 81444
rect 486200 81404 486206 81416
rect 487154 81404 487160 81416
rect 487212 81404 487218 81456
rect 117590 80152 117596 80164
rect 117516 80124 117596 80152
rect 117516 80028 117544 80124
rect 117590 80112 117596 80124
rect 117648 80112 117654 80164
rect 120350 80152 120356 80164
rect 120276 80124 120356 80152
rect 120276 80028 120304 80124
rect 120350 80112 120356 80124
rect 120408 80112 120414 80164
rect 220538 80112 220544 80164
rect 220596 80112 220602 80164
rect 272978 80112 272984 80164
rect 273036 80112 273042 80164
rect 299290 80112 299296 80164
rect 299348 80112 299354 80164
rect 351730 80112 351736 80164
rect 351788 80112 351794 80164
rect 506014 80112 506020 80164
rect 506072 80112 506078 80164
rect 220556 80028 220584 80112
rect 272996 80028 273024 80112
rect 299308 80028 299336 80112
rect 351748 80028 351776 80112
rect 506032 80028 506060 80112
rect 117498 79976 117504 80028
rect 117556 79976 117562 80028
rect 120258 79976 120264 80028
rect 120316 79976 120322 80028
rect 220538 79976 220544 80028
rect 220596 79976 220602 80028
rect 272978 79976 272984 80028
rect 273036 79976 273042 80028
rect 299290 79976 299296 80028
rect 299348 79976 299354 80028
rect 351730 79976 351736 80028
rect 351788 79976 351794 80028
rect 506014 79976 506020 80028
rect 506072 79976 506078 80028
rect 503714 79636 503720 79688
rect 503772 79676 503778 79688
rect 505738 79676 505744 79688
rect 503772 79648 505744 79676
rect 503772 79636 503778 79648
rect 505738 79636 505744 79648
rect 505796 79636 505802 79688
rect 485038 79160 485044 79212
rect 485096 79200 485102 79212
rect 486142 79200 486148 79212
rect 485096 79172 486148 79200
rect 485096 79160 485102 79172
rect 486142 79160 486148 79172
rect 486200 79160 486206 79212
rect 495986 78684 495992 78736
rect 496044 78724 496050 78736
rect 497458 78724 497464 78736
rect 496044 78696 497464 78724
rect 496044 78684 496050 78696
rect 497458 78684 497464 78696
rect 497516 78684 497522 78736
rect 505922 78004 505928 78056
rect 505980 78044 505986 78056
rect 506106 78044 506112 78056
rect 505980 78016 506112 78044
rect 505980 78004 505986 78016
rect 506106 78004 506112 78016
rect 506164 78004 506170 78056
rect 289722 77528 289728 77580
rect 289780 77528 289786 77580
rect 289740 77308 289768 77528
rect 289722 77256 289728 77308
rect 289780 77256 289786 77308
rect 436094 77296 436100 77308
rect 436055 77268 436100 77296
rect 436094 77256 436100 77268
rect 436152 77256 436158 77308
rect 500218 77296 500224 77308
rect 500179 77268 500224 77296
rect 500218 77256 500224 77268
rect 500276 77256 500282 77308
rect 76558 77188 76564 77240
rect 76616 77228 76622 77240
rect 580166 77228 580172 77240
rect 76616 77200 580172 77228
rect 76616 77188 76622 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 244274 77160 244280 77172
rect 244235 77132 244280 77160
rect 244274 77120 244280 77132
rect 244332 77120 244338 77172
rect 258074 77160 258080 77172
rect 258035 77132 258080 77160
rect 258074 77120 258080 77132
rect 258132 77120 258138 77172
rect 445846 77160 445852 77172
rect 445807 77132 445852 77160
rect 445846 77120 445852 77132
rect 445904 77120 445910 77172
rect 470686 77120 470692 77172
rect 470744 77160 470750 77172
rect 472342 77160 472348 77172
rect 470744 77132 472348 77160
rect 470744 77120 470750 77132
rect 472342 77120 472348 77132
rect 472400 77120 472406 77172
rect 494054 76576 494060 76628
rect 494112 76616 494118 76628
rect 495986 76616 495992 76628
rect 494112 76588 495992 76616
rect 494112 76576 494118 76588
rect 495986 76576 495992 76588
rect 496044 76576 496050 76628
rect 155954 75964 155960 76016
rect 156012 76004 156018 76016
rect 156138 76004 156144 76016
rect 156012 75976 156144 76004
rect 156012 75964 156018 75976
rect 156138 75964 156144 75976
rect 156196 75964 156202 76016
rect 161014 75896 161020 75948
rect 161072 75936 161078 75948
rect 161198 75936 161204 75948
rect 161072 75908 161204 75936
rect 161072 75896 161078 75908
rect 161198 75896 161204 75908
rect 161256 75896 161262 75948
rect 179322 75936 179328 75948
rect 179283 75908 179328 75936
rect 179322 75896 179328 75908
rect 179380 75896 179386 75948
rect 186222 75936 186228 75948
rect 186183 75908 186228 75936
rect 186222 75896 186228 75908
rect 186280 75896 186286 75948
rect 220633 75939 220691 75945
rect 220633 75905 220645 75939
rect 220679 75936 220691 75939
rect 220722 75936 220728 75948
rect 220679 75908 220728 75936
rect 220679 75905 220691 75908
rect 220633 75899 220691 75905
rect 220722 75896 220728 75908
rect 220780 75896 220786 75948
rect 223574 75936 223580 75948
rect 223535 75908 223580 75936
rect 223574 75896 223580 75908
rect 223632 75896 223638 75948
rect 378134 75936 378140 75948
rect 378095 75908 378140 75936
rect 378134 75896 378140 75908
rect 378192 75896 378198 75948
rect 511534 75936 511540 75948
rect 511495 75908 511540 75936
rect 511534 75896 511540 75908
rect 511592 75896 511598 75948
rect 524414 75936 524420 75948
rect 524375 75908 524420 75936
rect 524414 75896 524420 75908
rect 524472 75896 524478 75948
rect 532694 75936 532700 75948
rect 532655 75908 532700 75936
rect 532694 75896 532700 75908
rect 532752 75896 532758 75948
rect 110414 75868 110420 75880
rect 110375 75840 110420 75868
rect 110414 75828 110420 75840
rect 110472 75828 110478 75880
rect 497550 74576 497556 74588
rect 496464 74548 497556 74576
rect 494698 74468 494704 74520
rect 494756 74508 494762 74520
rect 496464 74508 496492 74548
rect 497550 74536 497556 74548
rect 497608 74536 497614 74588
rect 494756 74480 496492 74508
rect 494756 74468 494762 74480
rect 80057 73219 80115 73225
rect 80057 73185 80069 73219
rect 80103 73216 80115 73219
rect 80146 73216 80152 73228
rect 80103 73188 80152 73216
rect 80103 73185 80115 73188
rect 80057 73179 80115 73185
rect 80146 73176 80152 73188
rect 80204 73176 80210 73228
rect 492766 73176 492772 73228
rect 492824 73216 492830 73228
rect 494054 73216 494060 73228
rect 492824 73188 494060 73216
rect 492824 73176 492830 73188
rect 494054 73176 494060 73188
rect 494112 73176 494118 73228
rect 503622 73216 503628 73228
rect 498212 73188 503628 73216
rect 496722 73108 496728 73160
rect 496780 73148 496786 73160
rect 498212 73148 498240 73188
rect 503622 73176 503628 73188
rect 503680 73176 503686 73228
rect 496780 73120 498240 73148
rect 496780 73108 496786 73120
rect 499942 73108 499948 73160
rect 500000 73148 500006 73160
rect 500034 73148 500040 73160
rect 500000 73120 500040 73148
rect 500000 73108 500006 73120
rect 500034 73108 500040 73120
rect 500092 73108 500098 73160
rect 500678 73108 500684 73160
rect 500736 73148 500742 73160
rect 500770 73148 500776 73160
rect 500736 73120 500776 73148
rect 500736 73108 500742 73120
rect 500770 73108 500776 73120
rect 500828 73108 500834 73160
rect 482554 71748 482560 71800
rect 482612 71788 482618 71800
rect 485038 71788 485044 71800
rect 482612 71760 485044 71788
rect 482612 71748 482618 71760
rect 485038 71748 485044 71760
rect 485096 71748 485102 71800
rect 155954 70388 155960 70440
rect 156012 70388 156018 70440
rect 155972 70292 156000 70388
rect 156138 70292 156144 70304
rect 155972 70264 156144 70292
rect 156138 70252 156144 70264
rect 156196 70252 156202 70304
rect 79686 69776 79692 69828
rect 79744 69816 79750 69828
rect 79962 69816 79968 69828
rect 79744 69788 79968 69816
rect 79744 69776 79750 69788
rect 79962 69776 79968 69788
rect 80020 69776 80026 69828
rect 470686 69068 470692 69080
rect 469232 69040 470692 69068
rect 467098 68892 467104 68944
rect 467156 68932 467162 68944
rect 469232 68932 469260 69040
rect 470686 69028 470692 69040
rect 470744 69028 470750 69080
rect 492766 69068 492772 69080
rect 491312 69040 492772 69068
rect 491018 68960 491024 69012
rect 491076 69000 491082 69012
rect 491312 69000 491340 69040
rect 492766 69028 492772 69040
rect 492824 69028 492830 69080
rect 491076 68972 491340 69000
rect 491076 68960 491082 68972
rect 467156 68904 469260 68932
rect 467156 68892 467162 68904
rect 244274 67640 244280 67652
rect 244235 67612 244280 67640
rect 244274 67600 244280 67612
rect 244332 67600 244338 67652
rect 258074 67640 258080 67652
rect 258035 67612 258080 67640
rect 258074 67600 258080 67612
rect 258132 67600 258138 67652
rect 445846 67640 445852 67652
rect 445807 67612 445852 67640
rect 445846 67600 445852 67612
rect 445904 67600 445910 67652
rect 436094 67572 436100 67584
rect 436055 67544 436100 67572
rect 436094 67532 436100 67544
rect 436152 67532 436158 67584
rect 494238 66920 494244 66972
rect 494296 66960 494302 66972
rect 496722 66960 496728 66972
rect 494296 66932 496728 66960
rect 494296 66920 494302 66932
rect 496722 66920 496728 66932
rect 496780 66920 496786 66972
rect 80054 66240 80060 66292
rect 80112 66280 80118 66292
rect 80146 66280 80152 66292
rect 80112 66252 80152 66280
rect 80112 66240 80118 66252
rect 80146 66240 80152 66252
rect 80204 66240 80210 66292
rect 110414 66280 110420 66292
rect 110375 66252 110420 66280
rect 110414 66240 110420 66252
rect 110472 66240 110478 66292
rect 152826 66172 152832 66224
rect 152884 66212 152890 66224
rect 152918 66212 152924 66224
rect 152884 66184 152924 66212
rect 152884 66172 152890 66184
rect 152918 66172 152924 66184
rect 152976 66172 152982 66224
rect 155957 66215 156015 66221
rect 155957 66181 155969 66215
rect 156003 66212 156015 66215
rect 156138 66212 156144 66224
rect 156003 66184 156144 66212
rect 156003 66181 156015 66184
rect 155957 66175 156015 66181
rect 156138 66172 156144 66184
rect 156196 66172 156202 66224
rect 179322 66212 179328 66224
rect 179283 66184 179328 66212
rect 179322 66172 179328 66184
rect 179380 66172 179386 66224
rect 186222 66212 186228 66224
rect 186183 66184 186228 66212
rect 186222 66172 186228 66184
rect 186280 66172 186286 66224
rect 220722 66212 220728 66224
rect 220683 66184 220728 66212
rect 220722 66172 220728 66184
rect 220780 66172 220786 66224
rect 223574 66212 223580 66224
rect 223535 66184 223580 66212
rect 223574 66172 223580 66184
rect 223632 66172 223638 66224
rect 378134 66212 378140 66224
rect 378095 66184 378140 66212
rect 378134 66172 378140 66184
rect 378192 66172 378198 66224
rect 511534 66212 511540 66224
rect 511495 66184 511540 66212
rect 511534 66172 511540 66184
rect 511592 66172 511598 66224
rect 524414 66212 524420 66224
rect 524375 66184 524420 66212
rect 524414 66172 524420 66184
rect 524472 66172 524478 66224
rect 532694 66212 532700 66224
rect 532655 66184 532700 66212
rect 532694 66172 532700 66184
rect 532752 66172 532758 66224
rect 482554 64920 482560 64932
rect 480272 64892 482560 64920
rect 161014 64852 161020 64864
rect 160975 64824 161020 64852
rect 161014 64812 161020 64824
rect 161072 64812 161078 64864
rect 478874 64812 478880 64864
rect 478932 64852 478938 64864
rect 480272 64852 480300 64892
rect 482554 64880 482560 64892
rect 482612 64880 482618 64932
rect 487154 64880 487160 64932
rect 487212 64920 487218 64932
rect 491018 64920 491024 64932
rect 487212 64892 491024 64920
rect 487212 64880 487218 64892
rect 491018 64880 491024 64892
rect 491076 64880 491082 64932
rect 478932 64824 480300 64852
rect 478932 64812 478938 64824
rect 519538 64812 519544 64864
rect 519596 64852 519602 64864
rect 580166 64852 580172 64864
rect 519596 64824 580172 64852
rect 519596 64812 519602 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 2774 64540 2780 64592
rect 2832 64580 2838 64592
rect 4890 64580 4896 64592
rect 2832 64552 4896 64580
rect 2832 64540 2838 64552
rect 4890 64540 4896 64552
rect 4948 64540 4954 64592
rect 505830 63520 505836 63572
rect 505888 63560 505894 63572
rect 505922 63560 505928 63572
rect 505888 63532 505928 63560
rect 505888 63520 505894 63532
rect 505922 63520 505928 63532
rect 505980 63520 505986 63572
rect 117314 62092 117320 62144
rect 117372 62132 117378 62144
rect 117590 62132 117596 62144
rect 117372 62104 117596 62132
rect 117372 62092 117378 62104
rect 117590 62092 117596 62104
rect 117648 62092 117654 62144
rect 120074 62092 120080 62144
rect 120132 62132 120138 62144
rect 120350 62132 120356 62144
rect 120132 62104 120356 62132
rect 120132 62092 120138 62104
rect 120350 62092 120356 62104
rect 120408 62092 120414 62144
rect 478874 62132 478880 62144
rect 477512 62104 478880 62132
rect 476022 62024 476028 62076
rect 476080 62064 476086 62076
rect 477512 62064 477540 62104
rect 478874 62092 478880 62104
rect 478932 62092 478938 62144
rect 482278 62092 482284 62144
rect 482336 62132 482342 62144
rect 487154 62132 487160 62144
rect 482336 62104 487160 62132
rect 482336 62092 482342 62104
rect 487154 62092 487160 62104
rect 487212 62092 487218 62144
rect 491938 62092 491944 62144
rect 491996 62132 492002 62144
rect 494238 62132 494244 62144
rect 491996 62104 494244 62132
rect 491996 62092 492002 62104
rect 494238 62092 494244 62104
rect 494296 62092 494302 62144
rect 476080 62036 477540 62064
rect 476080 62024 476086 62036
rect 117590 60840 117596 60852
rect 117516 60812 117596 60840
rect 117516 60716 117544 60812
rect 117590 60800 117596 60812
rect 117648 60800 117654 60852
rect 120350 60840 120356 60852
rect 120276 60812 120356 60840
rect 120276 60716 120304 60812
rect 120350 60800 120356 60812
rect 120408 60800 120414 60852
rect 505830 60732 505836 60784
rect 505888 60732 505894 60784
rect 117498 60664 117504 60716
rect 117556 60664 117562 60716
rect 120258 60664 120264 60716
rect 120316 60664 120322 60716
rect 505848 60636 505876 60732
rect 505922 60636 505928 60648
rect 505848 60608 505928 60636
rect 505922 60596 505928 60608
rect 505980 60596 505986 60648
rect 436094 57984 436100 57996
rect 436055 57956 436100 57984
rect 436094 57944 436100 57956
rect 436152 57944 436158 57996
rect 476022 57984 476028 57996
rect 473372 57956 476028 57984
rect 244274 57916 244280 57928
rect 244235 57888 244280 57916
rect 244274 57876 244280 57888
rect 244332 57876 244338 57928
rect 258074 57916 258080 57928
rect 258035 57888 258080 57916
rect 258074 57876 258080 57888
rect 258132 57876 258138 57928
rect 289538 57876 289544 57928
rect 289596 57916 289602 57928
rect 289722 57916 289728 57928
rect 289596 57888 289728 57916
rect 289596 57876 289602 57888
rect 289722 57876 289728 57888
rect 289780 57876 289786 57928
rect 445846 57916 445852 57928
rect 445807 57888 445852 57916
rect 445846 57876 445852 57888
rect 445904 57876 445910 57928
rect 471974 57876 471980 57928
rect 472032 57916 472038 57928
rect 473372 57916 473400 57956
rect 476022 57944 476028 57956
rect 476080 57944 476086 57996
rect 472032 57888 473400 57916
rect 472032 57876 472038 57888
rect 436094 57848 436100 57860
rect 436055 57820 436100 57848
rect 436094 57808 436100 57820
rect 436152 57808 436158 57860
rect 465718 57604 465724 57656
rect 465776 57644 465782 57656
rect 467098 57644 467104 57656
rect 465776 57616 467104 57644
rect 465776 57604 465782 57616
rect 467098 57604 467104 57616
rect 467156 57604 467162 57656
rect 493594 57468 493600 57520
rect 493652 57508 493658 57520
rect 494698 57508 494704 57520
rect 493652 57480 494704 57508
rect 493652 57468 493658 57480
rect 494698 57468 494704 57480
rect 494756 57468 494762 57520
rect 110414 56720 110420 56772
rect 110472 56720 110478 56772
rect 110432 56636 110460 56720
rect 79594 56584 79600 56636
rect 79652 56624 79658 56636
rect 79686 56624 79692 56636
rect 79652 56596 79692 56624
rect 79652 56584 79658 56596
rect 79686 56584 79692 56596
rect 79744 56584 79750 56636
rect 110414 56584 110420 56636
rect 110472 56584 110478 56636
rect 155954 56624 155960 56636
rect 155915 56596 155960 56624
rect 155954 56584 155960 56596
rect 156012 56584 156018 56636
rect 179322 56624 179328 56636
rect 179283 56596 179328 56624
rect 179322 56584 179328 56596
rect 179380 56584 179386 56636
rect 186222 56624 186228 56636
rect 186183 56596 186228 56624
rect 186222 56584 186228 56596
rect 186280 56584 186286 56636
rect 220722 56624 220728 56636
rect 220683 56596 220728 56624
rect 220722 56584 220728 56596
rect 220780 56584 220786 56636
rect 223574 56624 223580 56636
rect 223535 56596 223580 56624
rect 223574 56584 223580 56596
rect 223632 56584 223638 56636
rect 378134 56624 378140 56636
rect 378095 56596 378140 56624
rect 378134 56584 378140 56596
rect 378192 56584 378198 56636
rect 511534 56624 511540 56636
rect 511495 56596 511540 56624
rect 511534 56584 511540 56596
rect 511592 56584 511598 56636
rect 524414 56624 524420 56636
rect 524375 56596 524420 56624
rect 524414 56584 524420 56596
rect 524472 56584 524478 56636
rect 532694 56624 532700 56636
rect 532655 56596 532700 56624
rect 532694 56584 532700 56596
rect 532752 56584 532758 56636
rect 110414 56488 110420 56500
rect 110375 56460 110420 56488
rect 110414 56448 110420 56460
rect 110472 56448 110478 56500
rect 161017 55267 161075 55273
rect 161017 55233 161029 55267
rect 161063 55264 161075 55267
rect 161382 55264 161388 55276
rect 161063 55236 161388 55264
rect 161063 55233 161075 55236
rect 161017 55227 161075 55233
rect 161382 55224 161388 55236
rect 161440 55224 161446 55276
rect 289538 53864 289544 53916
rect 289596 53904 289602 53916
rect 289722 53904 289728 53916
rect 289596 53876 289728 53904
rect 289596 53864 289602 53876
rect 289722 53864 289728 53876
rect 289780 53864 289786 53916
rect 490282 53864 490288 53916
rect 490340 53904 490346 53916
rect 491938 53904 491944 53916
rect 490340 53876 491944 53904
rect 490340 53864 490346 53876
rect 491938 53864 491944 53876
rect 491996 53864 492002 53916
rect 471974 53836 471980 53848
rect 469232 53808 471980 53836
rect 467098 53660 467104 53712
rect 467156 53700 467162 53712
rect 469232 53700 469260 53808
rect 471974 53796 471980 53808
rect 472032 53796 472038 53848
rect 481266 53796 481272 53848
rect 481324 53836 481330 53848
rect 482278 53836 482284 53848
rect 481324 53808 482284 53836
rect 481324 53796 481330 53808
rect 482278 53796 482284 53808
rect 482336 53796 482342 53848
rect 488534 53728 488540 53780
rect 488592 53768 488598 53780
rect 490282 53768 490288 53780
rect 488592 53740 490288 53768
rect 488592 53728 488598 53740
rect 490282 53728 490288 53740
rect 490340 53728 490346 53780
rect 467156 53672 469260 53700
rect 467156 53660 467162 53672
rect 79594 53388 79600 53440
rect 79652 53428 79658 53440
rect 79962 53428 79968 53440
rect 79652 53400 79968 53428
rect 79652 53388 79658 53400
rect 79962 53388 79968 53400
rect 80020 53388 80026 53440
rect 220538 51116 220544 51128
rect 220372 51088 220544 51116
rect 220372 51060 220400 51088
rect 220538 51076 220544 51088
rect 220596 51076 220602 51128
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 15838 51048 15844 51060
rect 3476 51020 15844 51048
rect 3476 51008 3482 51020
rect 15838 51008 15844 51020
rect 15896 51008 15902 51060
rect 220354 51008 220360 51060
rect 220412 51008 220418 51060
rect 272886 51008 272892 51060
rect 272944 51048 272950 51060
rect 273070 51048 273076 51060
rect 272944 51020 273076 51048
rect 272944 51008 272950 51020
rect 273070 51008 273076 51020
rect 273128 51008 273134 51060
rect 299198 51008 299204 51060
rect 299256 51048 299262 51060
rect 299382 51048 299388 51060
rect 299256 51020 299388 51048
rect 299256 51008 299262 51020
rect 299382 51008 299388 51020
rect 299440 51008 299446 51060
rect 351638 51008 351644 51060
rect 351696 51048 351702 51060
rect 351822 51048 351828 51060
rect 351696 51020 351828 51048
rect 351696 51008 351702 51020
rect 351822 51008 351828 51020
rect 351880 51008 351886 51060
rect 155954 50872 155960 50924
rect 156012 50912 156018 50924
rect 156138 50912 156144 50924
rect 156012 50884 156144 50912
rect 156012 50872 156018 50884
rect 156138 50872 156144 50884
rect 156196 50872 156202 50924
rect 491478 49784 491484 49836
rect 491536 49824 491542 49836
rect 493594 49824 493600 49836
rect 491536 49796 493600 49824
rect 491536 49784 491542 49796
rect 493594 49784 493600 49796
rect 493652 49784 493658 49836
rect 289630 48424 289636 48476
rect 289688 48424 289694 48476
rect 161106 48288 161112 48340
rect 161164 48328 161170 48340
rect 161382 48328 161388 48340
rect 161164 48300 161388 48328
rect 161164 48288 161170 48300
rect 161382 48288 161388 48300
rect 161440 48288 161446 48340
rect 244274 48328 244280 48340
rect 244235 48300 244280 48328
rect 244274 48288 244280 48300
rect 244332 48288 244338 48340
rect 258074 48328 258080 48340
rect 258035 48300 258080 48328
rect 258074 48288 258080 48300
rect 258132 48288 258138 48340
rect 289648 48272 289676 48424
rect 436094 48328 436100 48340
rect 436055 48300 436100 48328
rect 436094 48288 436100 48300
rect 436152 48288 436158 48340
rect 445846 48328 445852 48340
rect 445807 48300 445852 48328
rect 445846 48288 445852 48300
rect 445904 48288 445910 48340
rect 272981 48263 273039 48269
rect 272981 48229 272993 48263
rect 273027 48260 273039 48263
rect 273070 48260 273076 48272
rect 273027 48232 273076 48260
rect 273027 48229 273039 48232
rect 272981 48223 273039 48229
rect 273070 48220 273076 48232
rect 273128 48220 273134 48272
rect 289630 48220 289636 48272
rect 289688 48220 289694 48272
rect 299382 48260 299388 48272
rect 299343 48232 299388 48260
rect 299382 48220 299388 48232
rect 299440 48220 299446 48272
rect 351733 48263 351791 48269
rect 351733 48229 351745 48263
rect 351779 48260 351791 48263
rect 351822 48260 351828 48272
rect 351779 48232 351828 48260
rect 351779 48229 351791 48232
rect 351733 48223 351791 48229
rect 351822 48220 351828 48232
rect 351880 48220 351886 48272
rect 487890 47336 487896 47388
rect 487948 47376 487954 47388
rect 488534 47376 488540 47388
rect 487948 47348 488540 47376
rect 487948 47336 487954 47348
rect 488534 47336 488540 47348
rect 488592 47336 488598 47388
rect 488534 46996 488540 47048
rect 488592 47036 488598 47048
rect 491478 47036 491484 47048
rect 488592 47008 491484 47036
rect 488592 46996 488598 47008
rect 491478 46996 491484 47008
rect 491536 46996 491542 47048
rect 110414 46968 110420 46980
rect 110375 46940 110420 46968
rect 110414 46928 110420 46940
rect 110472 46928 110478 46980
rect 479610 46928 479616 46980
rect 479668 46968 479674 46980
rect 481266 46968 481272 46980
rect 479668 46940 481272 46968
rect 479668 46928 479674 46940
rect 481266 46928 481272 46940
rect 481324 46928 481330 46980
rect 156049 46903 156107 46909
rect 156049 46869 156061 46903
rect 156095 46900 156107 46903
rect 156138 46900 156144 46912
rect 156095 46872 156144 46900
rect 156095 46869 156107 46872
rect 156049 46863 156107 46869
rect 156138 46860 156144 46872
rect 156196 46860 156202 46912
rect 161106 46900 161112 46912
rect 161067 46872 161112 46900
rect 161106 46860 161112 46872
rect 161164 46860 161170 46912
rect 179233 46903 179291 46909
rect 179233 46869 179245 46903
rect 179279 46900 179291 46903
rect 179322 46900 179328 46912
rect 179279 46872 179328 46900
rect 179279 46869 179291 46872
rect 179233 46863 179291 46869
rect 179322 46860 179328 46872
rect 179380 46860 179386 46912
rect 186222 46900 186228 46912
rect 186183 46872 186228 46900
rect 186222 46860 186228 46872
rect 186280 46860 186286 46912
rect 220633 46903 220691 46909
rect 220633 46869 220645 46903
rect 220679 46900 220691 46903
rect 220722 46900 220728 46912
rect 220679 46872 220728 46900
rect 220679 46869 220691 46872
rect 220633 46863 220691 46869
rect 220722 46860 220728 46872
rect 220780 46860 220786 46912
rect 223574 46900 223580 46912
rect 223535 46872 223580 46900
rect 223574 46860 223580 46872
rect 223632 46860 223638 46912
rect 289722 46900 289728 46912
rect 289683 46872 289728 46900
rect 289722 46860 289728 46872
rect 289780 46860 289786 46912
rect 378134 46900 378140 46912
rect 378095 46872 378140 46900
rect 378134 46860 378140 46872
rect 378192 46860 378198 46912
rect 505833 46903 505891 46909
rect 505833 46869 505845 46903
rect 505879 46900 505891 46903
rect 505922 46900 505928 46912
rect 505879 46872 505928 46900
rect 505879 46869 505891 46872
rect 505833 46863 505891 46869
rect 505922 46860 505928 46872
rect 505980 46860 505986 46912
rect 511534 46900 511540 46912
rect 511495 46872 511540 46900
rect 511534 46860 511540 46872
rect 511592 46860 511598 46912
rect 524414 46900 524420 46912
rect 524375 46872 524420 46900
rect 524414 46860 524420 46872
rect 524472 46860 524478 46912
rect 532694 46900 532700 46912
rect 532655 46872 532700 46900
rect 532694 46860 532700 46872
rect 532752 46860 532758 46912
rect 82630 45608 82636 45620
rect 82591 45580 82636 45608
rect 82630 45568 82636 45580
rect 82688 45568 82694 45620
rect 121546 45568 121552 45620
rect 121604 45608 121610 45620
rect 121638 45608 121644 45620
rect 121604 45580 121644 45608
rect 121604 45568 121610 45580
rect 121638 45568 121644 45580
rect 121696 45568 121702 45620
rect 79962 44820 79968 44872
rect 80020 44860 80026 44872
rect 335354 44860 335360 44872
rect 80020 44832 335360 44860
rect 80020 44820 80026 44832
rect 335354 44820 335360 44832
rect 335412 44820 335418 44872
rect 82630 44180 82636 44192
rect 82591 44152 82636 44180
rect 82630 44140 82636 44152
rect 82688 44140 82694 44192
rect 83366 44140 83372 44192
rect 83424 44180 83430 44192
rect 83458 44180 83464 44192
rect 83424 44152 83464 44180
rect 83424 44140 83430 44152
rect 83458 44140 83464 44152
rect 83516 44140 83522 44192
rect 500678 44140 500684 44192
rect 500736 44180 500742 44192
rect 500770 44180 500776 44192
rect 500736 44152 500776 44180
rect 500736 44140 500742 44152
rect 500770 44140 500776 44152
rect 500828 44140 500834 44192
rect 156046 41392 156052 41404
rect 156007 41364 156052 41392
rect 156046 41352 156052 41364
rect 156104 41352 156110 41404
rect 540238 41352 540244 41404
rect 540296 41392 540302 41404
rect 580166 41392 580172 41404
rect 540296 41364 580172 41392
rect 540296 41352 540302 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 505833 41259 505891 41265
rect 505833 41225 505845 41259
rect 505879 41256 505891 41259
rect 505922 41256 505928 41268
rect 505879 41228 505928 41256
rect 505879 41225 505891 41228
rect 505833 41219 505891 41225
rect 505922 41216 505928 41228
rect 505980 41216 505986 41268
rect 486142 40128 486148 40180
rect 486200 40168 486206 40180
rect 487890 40168 487896 40180
rect 486200 40140 487896 40168
rect 486200 40128 486206 40140
rect 487890 40128 487896 40140
rect 487948 40128 487954 40180
rect 487798 39992 487804 40044
rect 487856 40032 487862 40044
rect 488534 40032 488540 40044
rect 487856 40004 488540 40032
rect 487856 39992 487862 40004
rect 488534 39992 488540 40004
rect 488592 39992 488598 40044
rect 117501 39355 117559 39361
rect 117501 39321 117513 39355
rect 117547 39352 117559 39355
rect 117682 39352 117688 39364
rect 117547 39324 117688 39352
rect 117547 39321 117559 39324
rect 117501 39315 117559 39321
rect 117682 39312 117688 39324
rect 117740 39312 117746 39364
rect 120261 39355 120319 39361
rect 120261 39321 120273 39355
rect 120307 39352 120319 39355
rect 120442 39352 120448 39364
rect 120307 39324 120448 39352
rect 120307 39321 120319 39324
rect 120261 39315 120319 39321
rect 120442 39312 120448 39324
rect 120500 39312 120506 39364
rect 459554 39312 459560 39364
rect 459612 39352 459618 39364
rect 465718 39352 465724 39364
rect 459612 39324 465724 39352
rect 459612 39312 459618 39324
rect 465718 39312 465724 39324
rect 465776 39312 465782 39364
rect 272978 38672 272984 38684
rect 272939 38644 272984 38672
rect 272978 38632 272984 38644
rect 273036 38632 273042 38684
rect 299290 38632 299296 38684
rect 299348 38672 299354 38684
rect 299385 38675 299443 38681
rect 299385 38672 299397 38675
rect 299348 38644 299397 38672
rect 299348 38632 299354 38644
rect 299385 38641 299397 38644
rect 299431 38641 299443 38675
rect 351730 38672 351736 38684
rect 351691 38644 351736 38672
rect 299385 38635 299443 38641
rect 351730 38632 351736 38644
rect 351788 38632 351794 38684
rect 244274 38604 244280 38616
rect 244235 38576 244280 38604
rect 244274 38564 244280 38576
rect 244332 38564 244338 38616
rect 258074 38604 258080 38616
rect 258035 38576 258080 38604
rect 258074 38564 258080 38576
rect 258132 38564 258138 38616
rect 436094 38604 436100 38616
rect 436055 38576 436100 38604
rect 436094 38564 436100 38576
rect 436152 38564 436158 38616
rect 445846 38604 445852 38616
rect 445807 38576 445852 38604
rect 445846 38564 445852 38576
rect 445904 38564 445910 38616
rect 476850 38564 476856 38616
rect 476908 38604 476914 38616
rect 479610 38604 479616 38616
rect 476908 38576 479616 38604
rect 476908 38564 476914 38576
rect 479610 38564 479616 38576
rect 479668 38564 479674 38616
rect 505830 38564 505836 38616
rect 505888 38604 505894 38616
rect 505922 38604 505928 38616
rect 505888 38576 505928 38604
rect 505888 38564 505894 38576
rect 505922 38564 505928 38576
rect 505980 38564 505986 38616
rect 88242 37884 88248 37936
rect 88300 37924 88306 37936
rect 505554 37924 505560 37936
rect 88300 37896 505560 37924
rect 88300 37884 88306 37896
rect 505554 37884 505560 37896
rect 505612 37884 505618 37936
rect 110414 37408 110420 37460
rect 110472 37408 110478 37460
rect 110432 37324 110460 37408
rect 110414 37272 110420 37324
rect 110472 37272 110478 37324
rect 161109 37315 161167 37321
rect 161109 37281 161121 37315
rect 161155 37312 161167 37315
rect 161198 37312 161204 37324
rect 161155 37284 161204 37312
rect 161155 37281 161167 37284
rect 161109 37275 161167 37281
rect 161198 37272 161204 37284
rect 161256 37272 161262 37324
rect 179230 37312 179236 37324
rect 179191 37284 179236 37312
rect 179230 37272 179236 37284
rect 179288 37272 179294 37324
rect 186222 37312 186228 37324
rect 186183 37284 186228 37312
rect 186222 37272 186228 37284
rect 186280 37272 186286 37324
rect 220633 37315 220691 37321
rect 220633 37281 220645 37315
rect 220679 37312 220691 37315
rect 220722 37312 220728 37324
rect 220679 37284 220728 37312
rect 220679 37281 220691 37284
rect 220633 37275 220691 37281
rect 220722 37272 220728 37284
rect 220780 37272 220786 37324
rect 223574 37312 223580 37324
rect 223535 37284 223580 37312
rect 223574 37272 223580 37284
rect 223632 37272 223638 37324
rect 289722 37312 289728 37324
rect 289683 37284 289728 37312
rect 289722 37272 289728 37284
rect 289780 37272 289786 37324
rect 361482 37272 361488 37324
rect 361540 37312 361546 37324
rect 362954 37312 362960 37324
rect 361540 37284 362960 37312
rect 361540 37272 361546 37284
rect 362954 37272 362960 37284
rect 363012 37272 363018 37324
rect 378134 37312 378140 37324
rect 378095 37284 378140 37312
rect 378134 37272 378140 37284
rect 378192 37272 378198 37324
rect 524414 37312 524420 37324
rect 524375 37284 524420 37312
rect 524414 37272 524420 37284
rect 524472 37272 524478 37324
rect 532694 37312 532700 37324
rect 532655 37284 532700 37312
rect 532694 37272 532700 37284
rect 532752 37272 532758 37324
rect 220446 37244 220452 37256
rect 220407 37216 220452 37244
rect 220446 37204 220452 37216
rect 220504 37204 220510 37256
rect 110414 37176 110420 37188
rect 110375 37148 110420 37176
rect 110414 37136 110420 37148
rect 110472 37136 110478 37188
rect 484210 36864 484216 36916
rect 484268 36904 484274 36916
rect 486142 36904 486148 36916
rect 484268 36876 486148 36904
rect 484268 36864 484274 36876
rect 486142 36864 486148 36876
rect 486200 36864 486206 36916
rect 457438 36320 457444 36372
rect 457496 36360 457502 36372
rect 459554 36360 459560 36372
rect 457496 36332 459560 36360
rect 457496 36320 457502 36332
rect 459554 36320 459560 36332
rect 459612 36320 459618 36372
rect 3142 35844 3148 35896
rect 3200 35884 3206 35896
rect 6178 35884 6184 35896
rect 3200 35856 6184 35884
rect 3200 35844 3206 35856
rect 6178 35844 6184 35856
rect 6236 35844 6242 35896
rect 83734 35844 83740 35896
rect 83792 35884 83798 35896
rect 83826 35884 83832 35896
rect 83792 35856 83832 35884
rect 83792 35844 83798 35856
rect 83826 35844 83832 35856
rect 83884 35844 83890 35896
rect 161198 32484 161204 32496
rect 161159 32456 161204 32484
rect 161198 32444 161204 32456
rect 161256 32444 161262 32496
rect 351730 31832 351736 31884
rect 351788 31832 351794 31884
rect 152921 31807 152979 31813
rect 152921 31773 152933 31807
rect 152967 31804 152979 31807
rect 153102 31804 153108 31816
rect 152967 31776 153108 31804
rect 152967 31773 152979 31776
rect 152921 31767 152979 31773
rect 153102 31764 153108 31776
rect 153160 31764 153166 31816
rect 351748 31748 351776 31832
rect 156046 31696 156052 31748
rect 156104 31736 156110 31748
rect 156230 31736 156236 31748
rect 156104 31708 156236 31736
rect 156104 31696 156110 31708
rect 156230 31696 156236 31708
rect 156288 31696 156294 31748
rect 351730 31696 351736 31748
rect 351788 31696 351794 31748
rect 505741 29699 505799 29705
rect 505741 29665 505753 29699
rect 505787 29696 505799 29699
rect 505830 29696 505836 29708
rect 505787 29668 505836 29696
rect 505787 29665 505799 29668
rect 505741 29659 505799 29665
rect 505830 29656 505836 29668
rect 505888 29656 505894 29708
rect 436094 29084 436100 29096
rect 436055 29056 436100 29084
rect 436094 29044 436100 29056
rect 436152 29044 436158 29096
rect 511534 29084 511540 29096
rect 511495 29056 511540 29084
rect 511534 29044 511540 29056
rect 511592 29044 511598 29096
rect 152918 29016 152924 29028
rect 152879 28988 152924 29016
rect 152918 28976 152924 28988
rect 152976 28976 152982 29028
rect 244274 29016 244280 29028
rect 244235 28988 244280 29016
rect 244274 28976 244280 28988
rect 244332 28976 244338 29028
rect 258074 29016 258080 29028
rect 258035 28988 258080 29016
rect 258074 28976 258080 28988
rect 258132 28976 258138 29028
rect 425606 28976 425612 29028
rect 425664 29016 425670 29028
rect 427814 29016 427820 29028
rect 425664 28988 427820 29016
rect 425664 28976 425670 28988
rect 427814 28976 427820 28988
rect 427872 28976 427878 29028
rect 445846 29016 445852 29028
rect 445807 28988 445852 29016
rect 445846 28976 445852 28988
rect 445904 28976 445910 29028
rect 484210 29016 484216 29028
rect 481652 28988 484216 29016
rect 156141 28951 156199 28957
rect 156141 28917 156153 28951
rect 156187 28948 156199 28951
rect 156230 28948 156236 28960
rect 156187 28920 156236 28948
rect 156187 28917 156199 28920
rect 156141 28911 156199 28917
rect 156230 28908 156236 28920
rect 156288 28908 156294 28960
rect 161474 28948 161480 28960
rect 161435 28920 161480 28948
rect 161474 28908 161480 28920
rect 161532 28908 161538 28960
rect 436094 28908 436100 28960
rect 436152 28948 436158 28960
rect 436186 28948 436192 28960
rect 436152 28920 436192 28948
rect 436152 28908 436158 28920
rect 436186 28908 436192 28920
rect 436244 28908 436250 28960
rect 480254 28908 480260 28960
rect 480312 28948 480318 28960
rect 481652 28948 481680 28988
rect 484210 28976 484216 28988
rect 484268 28976 484274 29028
rect 480312 28920 481680 28948
rect 480312 28908 480318 28920
rect 110414 27656 110420 27668
rect 110375 27628 110420 27656
rect 110414 27616 110420 27628
rect 110472 27616 110478 27668
rect 117501 27659 117559 27665
rect 117501 27625 117513 27659
rect 117547 27656 117559 27659
rect 117590 27656 117596 27668
rect 117547 27628 117596 27656
rect 117547 27625 117559 27628
rect 117501 27619 117559 27625
rect 117590 27616 117596 27628
rect 117648 27616 117654 27668
rect 120261 27659 120319 27665
rect 120261 27625 120273 27659
rect 120307 27656 120319 27659
rect 120350 27656 120356 27668
rect 120307 27628 120356 27656
rect 120307 27625 120319 27628
rect 120261 27619 120319 27625
rect 120350 27616 120356 27628
rect 120408 27616 120414 27668
rect 161198 27656 161204 27668
rect 161159 27628 161204 27656
rect 161198 27616 161204 27628
rect 161256 27616 161262 27668
rect 220449 27659 220507 27665
rect 220449 27625 220461 27659
rect 220495 27656 220507 27659
rect 220538 27656 220544 27668
rect 220495 27628 220544 27656
rect 220495 27625 220507 27628
rect 220449 27619 220507 27625
rect 220538 27616 220544 27628
rect 220596 27616 220602 27668
rect 152918 27588 152924 27600
rect 152879 27560 152924 27588
rect 152918 27548 152924 27560
rect 152976 27548 152982 27600
rect 178957 27591 179015 27597
rect 178957 27557 178969 27591
rect 179003 27588 179015 27591
rect 179322 27588 179328 27600
rect 179003 27560 179328 27588
rect 179003 27557 179015 27560
rect 178957 27551 179015 27557
rect 179322 27548 179328 27560
rect 179380 27548 179386 27600
rect 186041 27591 186099 27597
rect 186041 27557 186053 27591
rect 186087 27588 186099 27591
rect 186222 27588 186228 27600
rect 186087 27560 186228 27588
rect 186087 27557 186099 27560
rect 186041 27551 186099 27557
rect 186222 27548 186228 27560
rect 186280 27548 186286 27600
rect 220722 27588 220728 27600
rect 220683 27560 220728 27588
rect 220722 27548 220728 27560
rect 220780 27548 220786 27600
rect 223574 27588 223580 27600
rect 223535 27560 223580 27588
rect 223574 27548 223580 27560
rect 223632 27548 223638 27600
rect 289722 27588 289728 27600
rect 289683 27560 289728 27588
rect 289722 27548 289728 27560
rect 289780 27548 289786 27600
rect 299106 27588 299112 27600
rect 299067 27560 299112 27588
rect 299106 27548 299112 27560
rect 299164 27548 299170 27600
rect 362954 27548 362960 27600
rect 363012 27588 363018 27600
rect 363230 27588 363236 27600
rect 363012 27560 363236 27588
rect 363012 27548 363018 27560
rect 363230 27548 363236 27560
rect 363288 27548 363294 27600
rect 378134 27588 378140 27600
rect 378095 27560 378140 27588
rect 378134 27548 378140 27560
rect 378192 27548 378198 27600
rect 454678 27548 454684 27600
rect 454736 27588 454742 27600
rect 457438 27588 457444 27600
rect 454736 27560 457444 27588
rect 454736 27548 454742 27560
rect 457438 27548 457444 27560
rect 457496 27548 457502 27600
rect 511534 27588 511540 27600
rect 511495 27560 511540 27588
rect 511534 27548 511540 27560
rect 511592 27548 511598 27600
rect 524414 27588 524420 27600
rect 524375 27560 524420 27588
rect 524414 27548 524420 27560
rect 524472 27548 524478 27600
rect 532694 27588 532700 27600
rect 532655 27560 532700 27588
rect 532694 27548 532700 27560
rect 532752 27548 532758 27600
rect 478874 24828 478880 24880
rect 478932 24868 478938 24880
rect 480254 24868 480260 24880
rect 478932 24840 480260 24868
rect 478932 24828 478938 24840
rect 480254 24828 480260 24840
rect 480312 24828 480318 24880
rect 117409 22151 117467 22157
rect 117409 22117 117421 22151
rect 117455 22148 117467 22151
rect 117498 22148 117504 22160
rect 117455 22120 117504 22148
rect 117455 22117 117467 22120
rect 117409 22111 117467 22117
rect 117498 22108 117504 22120
rect 117556 22108 117562 22160
rect 272886 22040 272892 22092
rect 272944 22080 272950 22092
rect 273070 22080 273076 22092
rect 272944 22052 273076 22080
rect 272944 22040 272950 22052
rect 273070 22040 273076 22052
rect 273128 22040 273134 22092
rect 161106 20544 161112 20596
rect 161164 20584 161170 20596
rect 161290 20584 161296 20596
rect 161164 20556 161296 20584
rect 161164 20544 161170 20556
rect 161290 20544 161296 20556
rect 161348 20544 161354 20596
rect 478874 19428 478880 19440
rect 477420 19400 478880 19428
rect 156138 19360 156144 19372
rect 156099 19332 156144 19360
rect 156138 19320 156144 19332
rect 156196 19320 156202 19372
rect 131206 19292 131212 19304
rect 131167 19264 131212 19292
rect 131206 19252 131212 19264
rect 131264 19252 131270 19304
rect 244274 19292 244280 19304
rect 244235 19264 244280 19292
rect 244274 19252 244280 19264
rect 244332 19252 244338 19304
rect 258074 19252 258080 19304
rect 258132 19292 258138 19304
rect 258258 19292 258264 19304
rect 258132 19264 258264 19292
rect 258132 19252 258138 19264
rect 258258 19252 258264 19264
rect 258316 19252 258322 19304
rect 351733 19295 351791 19301
rect 351733 19261 351745 19295
rect 351779 19292 351791 19295
rect 351822 19292 351828 19304
rect 351779 19264 351828 19292
rect 351779 19261 351791 19264
rect 351733 19255 351791 19261
rect 351822 19252 351828 19264
rect 351880 19252 351886 19304
rect 427630 19252 427636 19304
rect 427688 19292 427694 19304
rect 427814 19292 427820 19304
rect 427688 19264 427820 19292
rect 427688 19252 427694 19264
rect 427814 19252 427820 19264
rect 427872 19252 427878 19304
rect 436094 19292 436100 19304
rect 436055 19264 436100 19292
rect 436094 19252 436100 19264
rect 436152 19252 436158 19304
rect 445846 19292 445852 19304
rect 445807 19264 445852 19292
rect 445846 19252 445852 19264
rect 445904 19252 445910 19304
rect 474826 19252 474832 19304
rect 474884 19292 474890 19304
rect 477420 19292 477448 19400
rect 478874 19388 478880 19400
rect 478932 19388 478938 19440
rect 474884 19264 477448 19292
rect 474884 19252 474890 19264
rect 463694 19184 463700 19236
rect 463752 19224 463758 19236
rect 467098 19224 467104 19236
rect 463752 19196 467104 19224
rect 463752 19184 463758 19196
rect 467098 19184 467104 19196
rect 467156 19184 467162 19236
rect 505738 19224 505744 19236
rect 505699 19196 505744 19224
rect 505738 19184 505744 19196
rect 505796 19184 505802 19236
rect 475010 18300 475016 18352
rect 475068 18340 475074 18352
rect 476850 18340 476856 18352
rect 475068 18312 476856 18340
rect 475068 18300 475074 18312
rect 476850 18300 476856 18312
rect 476908 18300 476914 18352
rect 110414 18096 110420 18148
rect 110472 18096 110478 18148
rect 110432 18012 110460 18096
rect 110414 17960 110420 18012
rect 110472 17960 110478 18012
rect 152921 18003 152979 18009
rect 152921 17969 152933 18003
rect 152967 18000 152979 18003
rect 153010 18000 153016 18012
rect 152967 17972 153016 18000
rect 152967 17969 152979 17972
rect 152921 17963 152979 17969
rect 153010 17960 153016 17972
rect 153068 17960 153074 18012
rect 161477 18003 161535 18009
rect 161477 17969 161489 18003
rect 161523 18000 161535 18003
rect 161566 18000 161572 18012
rect 161523 17972 161572 18000
rect 161523 17969 161535 17972
rect 161477 17963 161535 17969
rect 161566 17960 161572 17972
rect 161624 17960 161630 18012
rect 220722 18000 220728 18012
rect 220683 17972 220728 18000
rect 220722 17960 220728 17972
rect 220780 17960 220786 18012
rect 223574 18000 223580 18012
rect 223535 17972 223580 18000
rect 223574 17960 223580 17972
rect 223632 17960 223638 18012
rect 299109 18003 299167 18009
rect 299109 17969 299121 18003
rect 299155 18000 299167 18003
rect 299198 18000 299204 18012
rect 299155 17972 299204 18000
rect 299155 17969 299167 17972
rect 299109 17963 299167 17969
rect 299198 17960 299204 17972
rect 299256 17960 299262 18012
rect 378134 18000 378140 18012
rect 378095 17972 378140 18000
rect 378134 17960 378140 17972
rect 378192 17960 378198 18012
rect 511534 18000 511540 18012
rect 511495 17972 511540 18000
rect 511534 17960 511540 17972
rect 511592 17960 511598 18012
rect 524414 18000 524420 18012
rect 524375 17972 524420 18000
rect 524414 17960 524420 17972
rect 524472 17960 524478 18012
rect 340782 17484 340788 17536
rect 340840 17524 340846 17536
rect 505186 17524 505192 17536
rect 340840 17496 505192 17524
rect 340840 17484 340846 17496
rect 505186 17484 505192 17496
rect 505244 17484 505250 17536
rect 119522 17416 119528 17468
rect 119580 17456 119586 17468
rect 504174 17456 504180 17468
rect 119580 17428 504180 17456
rect 119580 17416 119586 17428
rect 504174 17416 504180 17428
rect 504232 17416 504238 17468
rect 99190 17348 99196 17400
rect 99248 17388 99254 17400
rect 504818 17388 504824 17400
rect 99248 17360 504824 17388
rect 99248 17348 99254 17360
rect 504818 17348 504824 17360
rect 504876 17348 504882 17400
rect 96522 17280 96528 17332
rect 96580 17320 96586 17332
rect 503898 17320 503904 17332
rect 96580 17292 503904 17320
rect 96580 17280 96586 17292
rect 503898 17280 503904 17292
rect 503956 17280 503962 17332
rect 56410 17212 56416 17264
rect 56468 17252 56474 17264
rect 506014 17252 506020 17264
rect 56468 17224 506020 17252
rect 56468 17212 56474 17224
rect 506014 17212 506020 17224
rect 506072 17212 506078 17264
rect 452654 17144 452660 17196
rect 452712 17184 452718 17196
rect 454678 17184 454684 17196
rect 452712 17156 454684 17184
rect 452712 17144 452718 17156
rect 454678 17144 454684 17156
rect 454736 17144 454742 17196
rect 471330 16600 471336 16652
rect 471388 16640 471394 16652
rect 474826 16640 474832 16652
rect 471388 16612 474832 16640
rect 471388 16600 471394 16612
rect 474826 16600 474832 16612
rect 474884 16600 474890 16652
rect 259362 15988 259368 16040
rect 259420 16028 259426 16040
rect 401594 16028 401600 16040
rect 259420 16000 401600 16028
rect 259420 15988 259426 16000
rect 401594 15988 401600 16000
rect 401652 15988 401658 16040
rect 293862 15920 293868 15972
rect 293920 15960 293926 15972
rect 505462 15960 505468 15972
rect 293920 15932 505468 15960
rect 293920 15920 293926 15932
rect 505462 15920 505468 15932
rect 505520 15920 505526 15972
rect 158622 15852 158628 15904
rect 158680 15892 158686 15904
rect 504082 15892 504088 15904
rect 158680 15864 504088 15892
rect 158680 15852 158686 15864
rect 504082 15852 504088 15864
rect 504140 15852 504146 15904
rect 117406 15212 117412 15224
rect 117367 15184 117412 15212
rect 117406 15172 117412 15184
rect 117464 15172 117470 15224
rect 120074 15172 120080 15224
rect 120132 15212 120138 15224
rect 120166 15212 120172 15224
rect 120132 15184 120172 15212
rect 120132 15172 120138 15184
rect 120166 15172 120172 15184
rect 120224 15172 120230 15224
rect 461854 15172 461860 15224
rect 461912 15212 461918 15224
rect 463694 15212 463700 15224
rect 461912 15184 463700 15212
rect 461912 15172 461918 15184
rect 463694 15172 463700 15184
rect 463752 15172 463758 15224
rect 295242 14832 295248 14884
rect 295300 14872 295306 14884
rect 302234 14872 302240 14884
rect 295300 14844 302240 14872
rect 295300 14832 295306 14844
rect 302234 14832 302240 14844
rect 302292 14832 302298 14884
rect 256602 14764 256608 14816
rect 256660 14804 256666 14816
rect 313274 14804 313280 14816
rect 256660 14776 313280 14804
rect 256660 14764 256666 14776
rect 313274 14764 313280 14776
rect 313332 14764 313338 14816
rect 272886 14696 272892 14748
rect 272944 14736 272950 14748
rect 333974 14736 333980 14748
rect 272944 14708 333980 14736
rect 272944 14696 272950 14708
rect 333974 14696 333980 14708
rect 334032 14696 334038 14748
rect 341889 14739 341947 14745
rect 341889 14705 341901 14739
rect 341935 14736 341947 14739
rect 474734 14736 474740 14748
rect 341935 14708 474740 14736
rect 341935 14705 341947 14708
rect 341889 14699 341947 14705
rect 474734 14696 474740 14708
rect 474792 14696 474798 14748
rect 226242 14628 226248 14680
rect 226300 14668 226306 14680
rect 365714 14668 365720 14680
rect 226300 14640 365720 14668
rect 226300 14628 226306 14640
rect 365714 14628 365720 14640
rect 365772 14628 365778 14680
rect 156138 14600 156144 14612
rect 156099 14572 156144 14600
rect 156138 14560 156144 14572
rect 156196 14560 156202 14612
rect 200022 14560 200028 14612
rect 200080 14600 200086 14612
rect 351914 14600 351920 14612
rect 200080 14572 351920 14600
rect 200080 14560 200086 14572
rect 351914 14560 351920 14572
rect 351972 14560 351978 14612
rect 81250 14492 81256 14544
rect 81308 14532 81314 14544
rect 367094 14532 367100 14544
rect 81308 14504 367100 14532
rect 81308 14492 81314 14504
rect 367094 14492 367100 14504
rect 367152 14492 367158 14544
rect 375190 14492 375196 14544
rect 375248 14532 375254 14544
rect 405734 14532 405740 14544
rect 375248 14504 405740 14532
rect 375248 14492 375254 14504
rect 405734 14492 405740 14504
rect 405792 14492 405798 14544
rect 79410 14424 79416 14476
rect 79468 14464 79474 14476
rect 412634 14464 412640 14476
rect 79468 14436 412640 14464
rect 79468 14424 79474 14436
rect 412634 14424 412640 14436
rect 412692 14424 412698 14476
rect 332502 13608 332508 13660
rect 332560 13648 332566 13660
rect 501966 13648 501972 13660
rect 332560 13620 501972 13648
rect 332560 13608 332566 13620
rect 501966 13608 501972 13620
rect 502024 13608 502030 13660
rect 335262 13540 335268 13592
rect 335320 13580 335326 13592
rect 527453 13583 527511 13589
rect 527453 13580 527465 13583
rect 335320 13552 527465 13580
rect 335320 13540 335326 13552
rect 527453 13549 527465 13552
rect 527499 13549 527511 13583
rect 527453 13543 527511 13549
rect 193122 13472 193128 13524
rect 193180 13512 193186 13524
rect 386414 13512 386420 13524
rect 193180 13484 386420 13512
rect 193180 13472 193186 13484
rect 386414 13472 386420 13484
rect 386472 13472 386478 13524
rect 245473 13447 245531 13453
rect 245473 13413 245485 13447
rect 245519 13444 245531 13447
rect 498194 13444 498200 13456
rect 245519 13416 498200 13444
rect 245519 13413 245531 13416
rect 245473 13407 245531 13413
rect 498194 13404 498200 13416
rect 498252 13404 498258 13456
rect 78674 13336 78680 13388
rect 78732 13376 78738 13388
rect 358814 13376 358820 13388
rect 78732 13348 358820 13376
rect 78732 13336 78738 13348
rect 358814 13336 358820 13348
rect 358872 13336 358878 13388
rect 371142 13336 371148 13388
rect 371200 13376 371206 13388
rect 541713 13379 541771 13385
rect 541713 13376 541725 13379
rect 371200 13348 541725 13376
rect 371200 13336 371206 13348
rect 541713 13345 541725 13348
rect 541759 13345 541771 13379
rect 541713 13339 541771 13345
rect 184842 13268 184848 13320
rect 184900 13308 184906 13320
rect 470594 13308 470600 13320
rect 184900 13280 470600 13308
rect 184900 13268 184906 13280
rect 470594 13268 470600 13280
rect 470652 13268 470658 13320
rect 220446 13200 220452 13252
rect 220504 13240 220510 13252
rect 284294 13240 284300 13252
rect 220504 13212 284300 13240
rect 220504 13200 220510 13212
rect 284294 13200 284300 13212
rect 284352 13200 284358 13252
rect 289630 13200 289636 13252
rect 289688 13240 289694 13252
rect 576854 13240 576860 13252
rect 289688 13212 576860 13240
rect 289688 13200 289694 13212
rect 576854 13200 576860 13212
rect 576912 13200 576918 13252
rect 79870 13132 79876 13184
rect 79928 13172 79934 13184
rect 377674 13172 377680 13184
rect 79928 13144 377680 13172
rect 79928 13132 79934 13144
rect 377674 13132 377680 13144
rect 377732 13132 377738 13184
rect 109954 13064 109960 13116
rect 110012 13104 110018 13116
rect 110322 13104 110328 13116
rect 110012 13076 110328 13104
rect 110012 13064 110018 13076
rect 110322 13064 110328 13076
rect 110380 13064 110386 13116
rect 219342 13064 219348 13116
rect 219400 13104 219406 13116
rect 565814 13104 565820 13116
rect 219400 13076 565820 13104
rect 219400 13064 219406 13076
rect 565814 13064 565820 13076
rect 565872 13064 565878 13116
rect 220541 12563 220599 12569
rect 220541 12529 220553 12563
rect 220587 12560 220599 12563
rect 220722 12560 220728 12572
rect 220587 12532 220728 12560
rect 220587 12529 220599 12532
rect 220541 12523 220599 12529
rect 220722 12520 220728 12532
rect 220780 12520 220786 12572
rect 393041 12563 393099 12569
rect 393041 12529 393053 12563
rect 393087 12560 393099 12563
rect 393222 12560 393228 12572
rect 393087 12532 393228 12560
rect 393087 12529 393099 12532
rect 393041 12523 393099 12529
rect 393222 12520 393228 12532
rect 393280 12520 393286 12572
rect 119522 12492 119528 12504
rect 119448 12464 119528 12492
rect 119448 12436 119476 12464
rect 119522 12452 119528 12464
rect 119580 12452 119586 12504
rect 135070 12492 135076 12504
rect 134904 12464 135076 12492
rect 134904 12436 134932 12464
rect 135070 12452 135076 12464
rect 135128 12452 135134 12504
rect 153010 12492 153016 12504
rect 152752 12464 153016 12492
rect 152752 12436 152780 12464
rect 153010 12452 153016 12464
rect 153068 12452 153074 12504
rect 221737 12495 221795 12501
rect 221737 12461 221749 12495
rect 221783 12492 221795 12495
rect 222102 12492 222108 12504
rect 221783 12464 222108 12492
rect 221783 12461 221795 12464
rect 221737 12455 221795 12461
rect 222102 12452 222108 12464
rect 222160 12452 222166 12504
rect 289722 12492 289728 12504
rect 289683 12464 289728 12492
rect 289722 12452 289728 12464
rect 289780 12452 289786 12504
rect 369946 12452 369952 12504
rect 370004 12452 370010 12504
rect 371234 12452 371240 12504
rect 371292 12452 371298 12504
rect 372614 12452 372620 12504
rect 372672 12452 372678 12504
rect 378134 12452 378140 12504
rect 378192 12452 378198 12504
rect 461854 12492 461860 12504
rect 459572 12464 461860 12492
rect 99006 12384 99012 12436
rect 99064 12424 99070 12436
rect 99190 12424 99196 12436
rect 99064 12396 99196 12424
rect 99064 12384 99070 12396
rect 99190 12384 99196 12396
rect 99248 12384 99254 12436
rect 106458 12384 106464 12436
rect 106516 12424 106522 12436
rect 107378 12424 107384 12436
rect 106516 12396 107384 12424
rect 106516 12384 106522 12396
rect 107378 12384 107384 12396
rect 107436 12384 107442 12436
rect 119430 12384 119436 12436
rect 119488 12384 119494 12436
rect 128354 12384 128360 12436
rect 128412 12424 128418 12436
rect 128998 12424 129004 12436
rect 128412 12396 129004 12424
rect 128412 12384 128418 12396
rect 128998 12384 129004 12396
rect 129056 12384 129062 12436
rect 134886 12384 134892 12436
rect 134944 12384 134950 12436
rect 152734 12384 152740 12436
rect 152792 12384 152798 12436
rect 196066 12384 196072 12436
rect 196124 12424 196130 12436
rect 196802 12424 196808 12436
rect 196124 12396 196808 12424
rect 196124 12384 196130 12396
rect 196802 12384 196808 12396
rect 196860 12384 196866 12436
rect 349154 12384 349160 12436
rect 349212 12424 349218 12436
rect 350258 12424 350264 12436
rect 349212 12396 350264 12424
rect 349212 12384 349218 12396
rect 350258 12384 350264 12396
rect 350316 12384 350322 12436
rect 351914 12384 351920 12436
rect 351972 12424 351978 12436
rect 352466 12424 352472 12436
rect 351972 12396 352472 12424
rect 351972 12384 351978 12396
rect 352466 12384 352472 12396
rect 352524 12384 352530 12436
rect 360194 12384 360200 12436
rect 360252 12424 360258 12436
rect 360930 12424 360936 12436
rect 360252 12396 360936 12424
rect 360252 12384 360258 12396
rect 360930 12384 360936 12396
rect 360988 12384 360994 12436
rect 367094 12384 367100 12436
rect 367152 12424 367158 12436
rect 368014 12424 368020 12436
rect 367152 12396 368020 12424
rect 367152 12384 367158 12396
rect 368014 12384 368020 12396
rect 368072 12384 368078 12436
rect 369964 12356 369992 12452
rect 370406 12356 370412 12368
rect 369964 12328 370412 12356
rect 370406 12316 370412 12328
rect 370464 12316 370470 12368
rect 371252 12356 371280 12452
rect 371602 12356 371608 12368
rect 371252 12328 371608 12356
rect 371602 12316 371608 12328
rect 371660 12316 371666 12368
rect 372632 12356 372660 12452
rect 372798 12356 372804 12368
rect 372632 12328 372804 12356
rect 372798 12316 372804 12328
rect 372856 12316 372862 12368
rect 378152 12356 378180 12452
rect 426434 12384 426440 12436
rect 426492 12424 426498 12436
rect 427538 12424 427544 12436
rect 426492 12396 427544 12424
rect 426492 12384 426498 12396
rect 427538 12384 427544 12396
rect 427596 12384 427602 12436
rect 458266 12384 458272 12436
rect 458324 12424 458330 12436
rect 459572 12424 459600 12464
rect 461854 12452 461860 12464
rect 461912 12452 461918 12504
rect 482830 12452 482836 12504
rect 482888 12492 482894 12504
rect 487798 12492 487804 12504
rect 482888 12464 487804 12492
rect 482888 12452 482894 12464
rect 487798 12452 487804 12464
rect 487856 12452 487862 12504
rect 511534 12492 511540 12504
rect 511460 12464 511540 12492
rect 511460 12436 511488 12464
rect 511534 12452 511540 12464
rect 511592 12452 511598 12504
rect 524414 12452 524420 12504
rect 524472 12452 524478 12504
rect 458324 12396 459600 12424
rect 458324 12384 458330 12396
rect 511442 12384 511448 12436
rect 511500 12384 511506 12436
rect 523034 12384 523040 12436
rect 523092 12424 523098 12436
rect 523862 12424 523868 12436
rect 523092 12396 523868 12424
rect 523092 12384 523098 12396
rect 523862 12384 523868 12396
rect 523920 12384 523926 12436
rect 378778 12356 378784 12368
rect 378152 12328 378784 12356
rect 378778 12316 378784 12328
rect 378836 12316 378842 12368
rect 524432 12356 524460 12452
rect 529934 12384 529940 12436
rect 529992 12424 529998 12436
rect 531038 12424 531044 12436
rect 529992 12396 531044 12424
rect 529992 12384 529998 12396
rect 531038 12384 531044 12396
rect 531096 12384 531102 12436
rect 534074 12384 534080 12436
rect 534132 12424 534138 12436
rect 534534 12424 534540 12436
rect 534132 12396 534540 12424
rect 534132 12384 534138 12396
rect 534534 12384 534540 12396
rect 534592 12384 534598 12436
rect 538214 12384 538220 12436
rect 538272 12424 538278 12436
rect 539318 12424 539324 12436
rect 538272 12396 539324 12424
rect 538272 12384 538278 12396
rect 539318 12384 539324 12396
rect 539376 12384 539382 12436
rect 542354 12384 542360 12436
rect 542412 12424 542418 12436
rect 542906 12424 542912 12436
rect 542412 12396 542912 12424
rect 542412 12384 542418 12396
rect 542906 12384 542912 12396
rect 542964 12384 542970 12436
rect 525058 12356 525064 12368
rect 524432 12328 525064 12356
rect 525058 12316 525064 12328
rect 525116 12316 525122 12368
rect 527450 12356 527456 12368
rect 527411 12328 527456 12356
rect 527450 12316 527456 12328
rect 527508 12316 527514 12368
rect 181346 12112 181352 12164
rect 181404 12152 181410 12164
rect 245654 12152 245660 12164
rect 181404 12124 245660 12152
rect 181404 12112 181410 12124
rect 245654 12112 245660 12124
rect 245712 12112 245718 12164
rect 138474 12044 138480 12096
rect 138532 12084 138538 12096
rect 251174 12084 251180 12096
rect 138532 12056 251180 12084
rect 138532 12044 138538 12056
rect 251174 12044 251180 12056
rect 251232 12044 251238 12096
rect 325602 12044 325608 12096
rect 325660 12084 325666 12096
rect 429930 12084 429936 12096
rect 325660 12056 429936 12084
rect 325660 12044 325666 12056
rect 429930 12044 429936 12056
rect 429988 12044 429994 12096
rect 154482 11976 154488 12028
rect 154540 12016 154546 12028
rect 230474 12016 230480 12028
rect 154540 11988 230480 12016
rect 154540 11976 154546 11988
rect 230474 11976 230480 11988
rect 230532 11976 230538 12028
rect 249610 11976 249616 12028
rect 249668 12016 249674 12028
rect 462038 12016 462044 12028
rect 249668 11988 462044 12016
rect 249668 11976 249674 11988
rect 462038 11976 462044 11988
rect 462096 11976 462102 12028
rect 216490 11908 216496 11960
rect 216548 11948 216554 11960
rect 506014 11948 506020 11960
rect 216548 11920 506020 11948
rect 216548 11908 216554 11920
rect 506014 11908 506020 11920
rect 506072 11908 506078 11960
rect 76558 11840 76564 11892
rect 76616 11880 76622 11892
rect 76834 11880 76840 11892
rect 76616 11852 76840 11880
rect 76616 11840 76622 11852
rect 76834 11840 76840 11852
rect 76892 11840 76898 11892
rect 155126 11840 155132 11892
rect 155184 11880 155190 11892
rect 477494 11880 477500 11892
rect 155184 11852 477500 11880
rect 155184 11840 155190 11852
rect 477494 11840 477500 11852
rect 477552 11840 477558 11892
rect 104802 11772 104808 11824
rect 104860 11812 104866 11824
rect 495342 11812 495348 11824
rect 104860 11784 495348 11812
rect 104860 11772 104866 11784
rect 495342 11772 495348 11784
rect 495400 11772 495406 11824
rect 84010 11704 84016 11756
rect 84068 11744 84074 11756
rect 509602 11744 509608 11756
rect 84068 11716 509608 11744
rect 84068 11704 84074 11716
rect 509602 11704 509608 11716
rect 509660 11704 509666 11756
rect 245470 11540 245476 11552
rect 245431 11512 245476 11540
rect 245470 11500 245476 11512
rect 245528 11500 245534 11552
rect 475010 11064 475016 11076
rect 471992 11036 475016 11064
rect 471606 10956 471612 11008
rect 471664 10996 471670 11008
rect 471992 10996 472020 11036
rect 475010 11024 475016 11036
rect 475068 11024 475074 11076
rect 471664 10968 472020 10996
rect 471664 10956 471670 10968
rect 445754 10888 445760 10940
rect 445812 10928 445818 10940
rect 452654 10928 452660 10940
rect 445812 10900 452660 10928
rect 445812 10888 445818 10900
rect 452654 10888 452660 10900
rect 452712 10888 452718 10940
rect 84102 10548 84108 10600
rect 84160 10588 84166 10600
rect 309134 10588 309140 10600
rect 84160 10560 309140 10588
rect 84160 10548 84166 10560
rect 309134 10548 309140 10560
rect 309192 10548 309198 10600
rect 354582 10548 354588 10600
rect 354640 10588 354646 10600
rect 546586 10588 546592 10600
rect 354640 10560 546592 10588
rect 354640 10548 354646 10560
rect 546586 10548 546592 10560
rect 546644 10548 546650 10600
rect 115842 10480 115848 10532
rect 115900 10520 115906 10532
rect 137278 10520 137284 10532
rect 115900 10492 137284 10520
rect 115900 10480 115906 10492
rect 137278 10480 137284 10492
rect 137336 10480 137342 10532
rect 173802 10480 173808 10532
rect 173860 10520 173866 10532
rect 191834 10520 191840 10532
rect 173860 10492 191840 10520
rect 173860 10480 173866 10492
rect 191834 10480 191840 10492
rect 191892 10480 191898 10532
rect 194410 10480 194416 10532
rect 194468 10520 194474 10532
rect 467834 10520 467840 10532
rect 194468 10492 467840 10520
rect 194468 10480 194474 10492
rect 467834 10480 467840 10492
rect 467892 10480 467898 10532
rect 79778 10412 79784 10464
rect 79836 10452 79842 10464
rect 383562 10452 383568 10464
rect 79836 10424 383568 10452
rect 79836 10412 79842 10424
rect 383562 10412 383568 10424
rect 383620 10412 383626 10464
rect 491202 10412 491208 10464
rect 491260 10452 491266 10464
rect 571426 10452 571432 10464
rect 491260 10424 571432 10452
rect 491260 10412 491266 10424
rect 571426 10412 571432 10424
rect 571484 10412 571490 10464
rect 79502 10344 79508 10396
rect 79560 10384 79566 10396
rect 404906 10384 404912 10396
rect 79560 10356 404912 10384
rect 79560 10344 79566 10356
rect 404906 10344 404912 10356
rect 404964 10344 404970 10396
rect 438762 10344 438768 10396
rect 438820 10384 438826 10396
rect 581086 10384 581092 10396
rect 438820 10356 581092 10384
rect 438820 10344 438826 10356
rect 581086 10344 581092 10356
rect 581144 10344 581150 10396
rect 135162 10276 135168 10328
rect 135220 10316 135226 10328
rect 491386 10316 491392 10328
rect 135220 10288 491392 10316
rect 135220 10276 135226 10288
rect 491386 10276 491392 10288
rect 491444 10276 491450 10328
rect 186038 9772 186044 9784
rect 185999 9744 186044 9772
rect 186038 9732 186044 9744
rect 186096 9732 186102 9784
rect 351730 9772 351736 9784
rect 351691 9744 351736 9772
rect 351730 9732 351736 9744
rect 351788 9732 351794 9784
rect 436094 9772 436100 9784
rect 436055 9744 436100 9772
rect 436094 9732 436100 9744
rect 436152 9732 436158 9784
rect 131206 9704 131212 9716
rect 131167 9676 131212 9704
rect 131206 9664 131212 9676
rect 131264 9664 131270 9716
rect 156141 9707 156199 9713
rect 156141 9673 156153 9707
rect 156187 9704 156199 9707
rect 156230 9704 156236 9716
rect 156187 9676 156236 9704
rect 156187 9673 156199 9676
rect 156141 9667 156199 9673
rect 156230 9664 156236 9676
rect 156288 9664 156294 9716
rect 161474 9664 161480 9716
rect 161532 9704 161538 9716
rect 161566 9704 161572 9716
rect 161532 9676 161572 9704
rect 161532 9664 161538 9676
rect 161566 9664 161572 9676
rect 161624 9664 161630 9716
rect 178954 9704 178960 9716
rect 178915 9676 178960 9704
rect 178954 9664 178960 9676
rect 179012 9664 179018 9716
rect 220538 9704 220544 9716
rect 220499 9676 220544 9704
rect 220538 9664 220544 9676
rect 220596 9664 220602 9716
rect 221734 9704 221740 9716
rect 221695 9676 221740 9704
rect 221734 9664 221740 9676
rect 221792 9664 221798 9716
rect 244274 9704 244280 9716
rect 244235 9676 244280 9704
rect 244274 9664 244280 9676
rect 244332 9664 244338 9716
rect 341886 9704 341892 9716
rect 341847 9676 341892 9704
rect 341886 9664 341892 9676
rect 341944 9664 341950 9716
rect 393038 9704 393044 9716
rect 392999 9676 393044 9704
rect 393038 9664 393044 9676
rect 393096 9664 393102 9716
rect 445846 9704 445852 9716
rect 445807 9676 445852 9704
rect 445846 9664 445852 9676
rect 445904 9664 445910 9716
rect 532697 9707 532755 9713
rect 532697 9673 532709 9707
rect 532743 9704 532755 9707
rect 533430 9704 533436 9716
rect 532743 9676 533436 9704
rect 532743 9673 532755 9676
rect 532697 9667 532755 9673
rect 533430 9664 533436 9676
rect 533488 9664 533494 9716
rect 541710 9704 541716 9716
rect 541671 9676 541716 9704
rect 541710 9664 541716 9676
rect 541768 9664 541774 9716
rect 99466 9596 99472 9648
rect 99524 9636 99530 9648
rect 100481 9639 100539 9645
rect 100481 9636 100493 9639
rect 99524 9608 100493 9636
rect 99524 9596 99530 9608
rect 100481 9605 100493 9608
rect 100527 9605 100539 9639
rect 134886 9636 134892 9648
rect 134847 9608 134892 9636
rect 100481 9599 100539 9605
rect 134886 9596 134892 9608
rect 134944 9596 134950 9648
rect 186038 9636 186044 9648
rect 185999 9608 186044 9636
rect 186038 9596 186044 9608
rect 186096 9596 186102 9648
rect 195606 9596 195612 9648
rect 195664 9596 195670 9648
rect 245470 9596 245476 9648
rect 245528 9636 245534 9648
rect 245654 9636 245660 9648
rect 245528 9608 245660 9636
rect 245528 9596 245534 9608
rect 245654 9596 245660 9608
rect 245712 9596 245718 9648
rect 258074 9596 258080 9648
rect 258132 9636 258138 9648
rect 258629 9639 258687 9645
rect 258629 9636 258641 9639
rect 258132 9608 258641 9636
rect 258132 9596 258138 9608
rect 258629 9605 258641 9608
rect 258675 9605 258687 9639
rect 351730 9636 351736 9648
rect 351691 9608 351736 9636
rect 258629 9599 258687 9605
rect 351730 9596 351736 9608
rect 351788 9596 351794 9648
rect 370406 9636 370412 9648
rect 370367 9608 370412 9636
rect 370406 9596 370412 9608
rect 370464 9596 370470 9648
rect 371602 9636 371608 9648
rect 371563 9608 371608 9636
rect 371602 9596 371608 9608
rect 371660 9596 371666 9648
rect 372798 9636 372804 9648
rect 372759 9608 372804 9636
rect 372798 9596 372804 9608
rect 372856 9596 372862 9648
rect 377582 9636 377588 9648
rect 377543 9608 377588 9636
rect 377582 9596 377588 9608
rect 377640 9596 377646 9648
rect 378778 9636 378784 9648
rect 378739 9608 378784 9636
rect 378778 9596 378784 9608
rect 378836 9596 378842 9648
rect 427814 9596 427820 9648
rect 427872 9636 427878 9648
rect 428737 9639 428795 9645
rect 428737 9636 428749 9639
rect 427872 9608 428749 9636
rect 427872 9596 427878 9608
rect 428737 9605 428749 9608
rect 428783 9605 428795 9639
rect 428737 9599 428795 9605
rect 436094 9596 436100 9648
rect 436152 9636 436158 9648
rect 437017 9639 437075 9645
rect 437017 9636 437029 9639
rect 436152 9608 437029 9636
rect 436152 9596 436158 9608
rect 437017 9605 437029 9608
rect 437063 9605 437075 9639
rect 437017 9599 437075 9605
rect 525058 9596 525064 9648
rect 525116 9596 525122 9648
rect 527450 9596 527456 9648
rect 527508 9596 527514 9648
rect 195624 9512 195652 9596
rect 525076 9512 525104 9596
rect 527468 9512 527496 9596
rect 195606 9460 195612 9512
rect 195664 9460 195670 9512
rect 525058 9460 525064 9512
rect 525116 9460 525122 9512
rect 527450 9460 527456 9512
rect 527508 9460 527514 9512
rect 83826 9392 83832 9444
rect 83884 9432 83890 9444
rect 171778 9432 171784 9444
rect 83884 9404 171784 9432
rect 83884 9392 83890 9404
rect 171778 9392 171784 9404
rect 171836 9392 171842 9444
rect 81710 9324 81716 9376
rect 81768 9364 81774 9376
rect 222930 9364 222936 9376
rect 81768 9336 222936 9364
rect 81768 9324 81774 9336
rect 222930 9324 222936 9336
rect 222988 9324 222994 9376
rect 126606 9256 126612 9308
rect 126664 9296 126670 9308
rect 287146 9296 287152 9308
rect 126664 9268 287152 9296
rect 126664 9256 126670 9268
rect 287146 9256 287152 9268
rect 287204 9256 287210 9308
rect 83458 9188 83464 9240
rect 83516 9228 83522 9240
rect 308582 9228 308588 9240
rect 83516 9200 308588 9228
rect 83516 9188 83522 9200
rect 308582 9188 308588 9200
rect 308640 9188 308646 9240
rect 413922 9188 413928 9240
rect 413980 9228 413986 9240
rect 501230 9228 501236 9240
rect 413980 9200 501236 9228
rect 413980 9188 413986 9200
rect 501230 9188 501236 9200
rect 501288 9188 501294 9240
rect 81434 9120 81440 9172
rect 81492 9160 81498 9172
rect 358538 9160 358544 9172
rect 81492 9132 358544 9160
rect 81492 9120 81498 9132
rect 358538 9120 358544 9132
rect 358596 9120 358602 9172
rect 436002 9120 436008 9172
rect 436060 9160 436066 9172
rect 526254 9160 526260 9172
rect 436060 9132 526260 9160
rect 436060 9120 436066 9132
rect 526254 9120 526260 9132
rect 526312 9120 526318 9172
rect 150342 9052 150348 9104
rect 150400 9092 150406 9104
rect 540514 9092 540520 9104
rect 150400 9064 540520 9092
rect 150400 9052 150406 9064
rect 540514 9052 540520 9064
rect 540572 9052 540578 9104
rect 89530 8984 89536 9036
rect 89588 9024 89594 9036
rect 519078 9024 519084 9036
rect 89588 8996 519084 9024
rect 89588 8984 89594 8996
rect 519078 8984 519084 8996
rect 519136 8984 519142 9036
rect 108942 8916 108948 8968
rect 109000 8956 109006 8968
rect 551186 8956 551192 8968
rect 109000 8928 551192 8956
rect 109000 8916 109006 8928
rect 551186 8916 551192 8928
rect 551244 8916 551250 8968
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 508682 8276 508688 8288
rect 3476 8248 508688 8276
rect 3476 8236 3482 8248
rect 508682 8236 508688 8248
rect 508740 8236 508746 8288
rect 117130 8168 117136 8220
rect 117188 8208 117194 8220
rect 253934 8208 253940 8220
rect 117188 8180 253940 8208
rect 117188 8168 117194 8180
rect 253934 8168 253940 8180
rect 253992 8168 253998 8220
rect 262122 8168 262128 8220
rect 262180 8208 262186 8220
rect 400214 8208 400220 8220
rect 262180 8180 400220 8208
rect 262180 8168 262186 8180
rect 400214 8168 400220 8180
rect 400272 8168 400278 8220
rect 113542 8100 113548 8152
rect 113600 8140 113606 8152
rect 327074 8140 327080 8152
rect 113600 8112 327080 8140
rect 113600 8100 113606 8112
rect 327074 8100 327080 8112
rect 327132 8100 327138 8152
rect 171042 8032 171048 8084
rect 171100 8072 171106 8084
rect 457254 8072 457260 8084
rect 171100 8044 457260 8072
rect 171100 8032 171106 8044
rect 457254 8032 457260 8044
rect 457312 8032 457318 8084
rect 102778 7964 102784 8016
rect 102836 8004 102842 8016
rect 408494 8004 408500 8016
rect 102836 7976 408500 8004
rect 102836 7964 102842 7976
rect 408494 7964 408500 7976
rect 408552 7964 408558 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 340874 7936 340880 7948
rect 33928 7908 340880 7936
rect 33928 7896 33934 7908
rect 340874 7896 340880 7908
rect 340932 7896 340938 7948
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 329834 7868 329840 7880
rect 18380 7840 329840 7868
rect 18380 7828 18386 7840
rect 329834 7828 329840 7840
rect 329892 7828 329898 7880
rect 124214 7760 124220 7812
rect 124272 7800 124278 7812
rect 438854 7800 438860 7812
rect 124272 7772 438860 7800
rect 124272 7760 124278 7772
rect 438854 7760 438860 7772
rect 438912 7760 438918 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 346394 7732 346400 7744
rect 21968 7704 346400 7732
rect 21968 7692 21974 7704
rect 346394 7692 346400 7704
rect 346452 7692 346458 7744
rect 357342 7692 357348 7744
rect 357400 7732 357406 7744
rect 402974 7732 402980 7744
rect 357400 7704 402980 7732
rect 357400 7692 357406 7704
rect 402974 7692 402980 7704
rect 403032 7692 403038 7744
rect 44542 7624 44548 7676
rect 44600 7664 44606 7676
rect 396166 7664 396172 7676
rect 44600 7636 396172 7664
rect 44600 7624 44606 7636
rect 396166 7624 396172 7636
rect 396224 7624 396230 7676
rect 401594 7624 401600 7676
rect 401652 7664 401658 7676
rect 402514 7664 402520 7676
rect 401652 7636 402520 7664
rect 401652 7624 401658 7636
rect 402514 7624 402520 7636
rect 402572 7624 402578 7676
rect 419534 7624 419540 7676
rect 419592 7664 419598 7676
rect 420362 7664 420368 7676
rect 419592 7636 420368 7664
rect 419592 7624 419598 7636
rect 420362 7624 420368 7636
rect 420420 7624 420426 7676
rect 433334 7624 433340 7676
rect 433392 7664 433398 7676
rect 434622 7664 434628 7676
rect 433392 7636 434628 7664
rect 433392 7624 433398 7636
rect 434622 7624 434628 7636
rect 434680 7624 434686 7676
rect 459462 7624 459468 7676
rect 459520 7664 459526 7676
rect 529842 7664 529848 7676
rect 459520 7636 529848 7664
rect 459520 7624 459526 7636
rect 529842 7624 529848 7636
rect 529900 7624 529906 7676
rect 50522 7556 50528 7608
rect 50580 7596 50586 7608
rect 484394 7596 484400 7608
rect 50580 7568 484400 7596
rect 50580 7556 50586 7568
rect 484394 7556 484400 7568
rect 484452 7556 484458 7608
rect 520274 7556 520280 7608
rect 520332 7596 520338 7608
rect 521470 7596 521476 7608
rect 520332 7568 521476 7596
rect 520332 7556 520338 7568
rect 521470 7556 521476 7568
rect 521528 7556 521534 7608
rect 536834 7556 536840 7608
rect 536892 7596 536898 7608
rect 538122 7596 538128 7608
rect 536892 7568 538128 7596
rect 536892 7556 536898 7568
rect 538122 7556 538128 7568
rect 538180 7556 538186 7608
rect 81526 7488 81532 7540
rect 81584 7528 81590 7540
rect 183738 7528 183744 7540
rect 81584 7500 183744 7528
rect 81584 7488 81590 7500
rect 183738 7488 183744 7500
rect 183796 7488 183802 7540
rect 287054 7488 287060 7540
rect 287112 7528 287118 7540
rect 288342 7528 288348 7540
rect 287112 7500 288348 7528
rect 287112 7488 287118 7500
rect 288342 7488 288348 7500
rect 288400 7488 288406 7540
rect 365714 7488 365720 7540
rect 365772 7528 365778 7540
rect 366910 7528 366916 7540
rect 365772 7500 366916 7528
rect 365772 7488 365778 7500
rect 366910 7488 366916 7500
rect 366968 7488 366974 7540
rect 478046 7352 478052 7404
rect 478104 7392 478110 7404
rect 482830 7392 482836 7404
rect 478104 7364 482836 7392
rect 478104 7352 478110 7364
rect 482830 7352 482836 7364
rect 482888 7352 482894 7404
rect 500034 7216 500040 7268
rect 500092 7256 500098 7268
rect 500678 7256 500684 7268
rect 500092 7228 500684 7256
rect 500092 7216 500098 7228
rect 500678 7216 500684 7228
rect 500736 7216 500742 7268
rect 469306 7148 469312 7200
rect 469364 7188 469370 7200
rect 471606 7188 471612 7200
rect 469364 7160 471612 7188
rect 469364 7148 469370 7160
rect 471606 7148 471612 7160
rect 471664 7148 471670 7200
rect 76558 6876 76564 6928
rect 76616 6916 76622 6928
rect 76926 6916 76932 6928
rect 76616 6888 76932 6916
rect 76616 6876 76622 6888
rect 76926 6876 76932 6888
rect 76984 6876 76990 6928
rect 82630 6876 82636 6928
rect 82688 6876 82694 6928
rect 120166 6876 120172 6928
rect 120224 6916 120230 6928
rect 120258 6916 120264 6928
rect 120224 6888 120264 6916
rect 120224 6876 120230 6888
rect 120258 6876 120264 6888
rect 120316 6876 120322 6928
rect 82538 6672 82544 6724
rect 82596 6712 82602 6724
rect 82648 6712 82676 6876
rect 110414 6808 110420 6860
rect 110472 6848 110478 6860
rect 111153 6851 111211 6857
rect 111153 6848 111165 6851
rect 110472 6820 111165 6848
rect 110472 6808 110478 6820
rect 111153 6817 111165 6820
rect 111199 6817 111211 6851
rect 111153 6811 111211 6817
rect 117406 6808 117412 6860
rect 117464 6848 117470 6860
rect 118234 6848 118240 6860
rect 117464 6820 118240 6848
rect 117464 6808 117470 6820
rect 118234 6808 118240 6820
rect 118292 6808 118298 6860
rect 395430 6808 395436 6860
rect 395488 6848 395494 6860
rect 510890 6848 510896 6860
rect 395488 6820 510896 6848
rect 395488 6808 395494 6820
rect 510890 6808 510896 6820
rect 510948 6808 510954 6860
rect 382366 6740 382372 6792
rect 382424 6780 382430 6792
rect 511074 6780 511080 6792
rect 382424 6752 511080 6780
rect 382424 6740 382430 6752
rect 511074 6740 511080 6752
rect 511132 6740 511138 6792
rect 82596 6684 82676 6712
rect 82596 6672 82602 6684
rect 376386 6672 376392 6724
rect 376444 6712 376450 6724
rect 507762 6712 507768 6724
rect 376444 6684 507768 6712
rect 376444 6672 376450 6684
rect 507762 6672 507768 6684
rect 507820 6672 507826 6724
rect 77018 6604 77024 6656
rect 77076 6644 77082 6656
rect 159910 6644 159916 6656
rect 77076 6616 159916 6644
rect 77076 6604 77082 6616
rect 159910 6604 159916 6616
rect 159968 6604 159974 6656
rect 345474 6604 345480 6656
rect 345532 6644 345538 6656
rect 509510 6644 509516 6656
rect 345532 6616 509516 6644
rect 345532 6604 345538 6616
rect 509510 6604 509516 6616
rect 509568 6604 509574 6656
rect 78306 6536 78312 6588
rect 78364 6576 78370 6588
rect 261018 6576 261024 6588
rect 78364 6548 261024 6576
rect 78364 6536 78370 6548
rect 261018 6536 261024 6548
rect 261076 6536 261082 6588
rect 346670 6536 346676 6588
rect 346728 6576 346734 6588
rect 510982 6576 510988 6588
rect 346728 6548 510988 6576
rect 346728 6536 346734 6548
rect 510982 6536 510988 6548
rect 511040 6536 511046 6588
rect 78490 6468 78496 6520
rect 78548 6508 78554 6520
rect 281258 6508 281264 6520
rect 78548 6480 281264 6508
rect 78548 6468 78554 6480
rect 281258 6468 281264 6480
rect 281316 6468 281322 6520
rect 299198 6468 299204 6520
rect 299256 6508 299262 6520
rect 520274 6508 520280 6520
rect 299256 6480 520280 6508
rect 299256 6468 299262 6480
rect 520274 6468 520280 6480
rect 520332 6468 520338 6520
rect 99282 6400 99288 6452
rect 99340 6440 99346 6452
rect 409690 6440 409696 6452
rect 99340 6412 409696 6440
rect 99340 6400 99346 6412
rect 409690 6400 409696 6412
rect 409748 6400 409754 6452
rect 410886 6400 410892 6452
rect 410944 6440 410950 6452
rect 502426 6440 502432 6452
rect 410944 6412 502432 6440
rect 410944 6400 410950 6412
rect 502426 6400 502432 6412
rect 502484 6400 502490 6452
rect 78398 6332 78404 6384
rect 78456 6372 78462 6384
rect 417970 6372 417976 6384
rect 78456 6344 417976 6372
rect 78456 6332 78462 6344
rect 417970 6332 417976 6344
rect 418028 6332 418034 6384
rect 423950 6332 423956 6384
rect 424008 6372 424014 6384
rect 509418 6372 509424 6384
rect 424008 6344 509424 6372
rect 424008 6332 424014 6344
rect 509418 6332 509424 6344
rect 509476 6332 509482 6384
rect 74350 6264 74356 6316
rect 74408 6304 74414 6316
rect 472710 6304 472716 6316
rect 74408 6276 472716 6304
rect 74408 6264 74414 6276
rect 472710 6264 472716 6276
rect 472768 6264 472774 6316
rect 497734 6264 497740 6316
rect 497792 6304 497798 6316
rect 510798 6304 510804 6316
rect 497792 6276 510804 6304
rect 497792 6264 497798 6276
rect 510798 6264 510804 6276
rect 510856 6264 510862 6316
rect 77754 6196 77760 6248
rect 77812 6236 77818 6248
rect 502426 6236 502432 6248
rect 77812 6208 502432 6236
rect 77812 6196 77818 6208
rect 502426 6196 502432 6208
rect 502484 6196 502490 6248
rect 74442 6128 74448 6180
rect 74500 6168 74506 6180
rect 516778 6168 516784 6180
rect 74500 6140 516784 6168
rect 74500 6128 74506 6140
rect 516778 6128 516784 6140
rect 516836 6128 516842 6180
rect 432322 6060 432328 6112
rect 432380 6100 432386 6112
rect 505738 6100 505744 6112
rect 432380 6072 505744 6100
rect 432380 6060 432386 6072
rect 505738 6060 505744 6072
rect 505796 6060 505802 6112
rect 451366 5992 451372 6044
rect 451424 6032 451430 6044
rect 508314 6032 508320 6044
rect 451424 6004 508320 6032
rect 451424 5992 451430 6004
rect 508314 5992 508320 6004
rect 508372 5992 508378 6044
rect 471238 5652 471244 5704
rect 471296 5692 471302 5704
rect 478046 5692 478052 5704
rect 471296 5664 478052 5692
rect 471296 5652 471302 5664
rect 478046 5652 478052 5664
rect 478104 5652 478110 5704
rect 469214 5516 469220 5568
rect 469272 5556 469278 5568
rect 471330 5556 471336 5568
rect 469272 5528 471336 5556
rect 469272 5516 469278 5528
rect 471330 5516 471336 5528
rect 471388 5516 471394 5568
rect 499942 5516 499948 5568
rect 500000 5556 500006 5568
rect 500126 5556 500132 5568
rect 500000 5528 500132 5556
rect 500000 5516 500006 5528
rect 500126 5516 500132 5528
rect 500184 5516 500190 5568
rect 256234 5448 256240 5500
rect 256292 5488 256298 5500
rect 296714 5488 296720 5500
rect 256292 5460 296720 5488
rect 256292 5448 256298 5460
rect 296714 5448 296720 5460
rect 296772 5448 296778 5500
rect 297818 5448 297824 5500
rect 297876 5488 297882 5500
rect 418154 5488 418160 5500
rect 297876 5460 418160 5488
rect 297876 5448 297882 5460
rect 418154 5448 418160 5460
rect 418212 5448 418218 5500
rect 442902 5448 442908 5500
rect 442960 5488 442966 5500
rect 467926 5488 467932 5500
rect 442960 5460 467932 5488
rect 442960 5448 442966 5460
rect 467926 5448 467932 5460
rect 467984 5448 467990 5500
rect 213822 5380 213828 5432
rect 213880 5420 213886 5432
rect 294322 5420 294328 5432
rect 213880 5392 294328 5420
rect 213880 5380 213886 5392
rect 294322 5380 294328 5392
rect 294380 5380 294386 5432
rect 300302 5380 300308 5432
rect 300360 5420 300366 5432
rect 445754 5420 445760 5432
rect 300360 5392 445760 5420
rect 300360 5380 300366 5392
rect 445754 5380 445760 5392
rect 445812 5380 445818 5432
rect 245562 5312 245568 5364
rect 245620 5352 245626 5364
rect 394234 5352 394240 5364
rect 245620 5324 394240 5352
rect 245620 5312 245626 5324
rect 394234 5312 394240 5324
rect 394292 5312 394298 5364
rect 415670 5312 415676 5364
rect 415728 5352 415734 5364
rect 491294 5352 491300 5364
rect 415728 5324 491300 5352
rect 415728 5312 415734 5324
rect 491294 5312 491300 5324
rect 491352 5312 491358 5364
rect 176562 5244 176568 5296
rect 176620 5284 176626 5296
rect 183554 5284 183560 5296
rect 176620 5256 183560 5284
rect 176620 5244 176626 5256
rect 183554 5244 183560 5256
rect 183612 5244 183618 5296
rect 201586 5244 201592 5296
rect 201644 5284 201650 5296
rect 357434 5284 357440 5296
rect 201644 5256 357440 5284
rect 201644 5244 201650 5256
rect 357434 5244 357440 5256
rect 357492 5244 357498 5296
rect 373902 5244 373908 5296
rect 373960 5284 373966 5296
rect 476298 5284 476304 5296
rect 373960 5256 476304 5284
rect 373960 5244 373966 5256
rect 476298 5244 476304 5256
rect 476356 5244 476362 5296
rect 127802 5176 127808 5228
rect 127860 5216 127866 5228
rect 281534 5216 281540 5228
rect 127860 5188 281540 5216
rect 127860 5176 127866 5188
rect 281534 5176 281540 5188
rect 281592 5176 281598 5228
rect 291930 5176 291936 5228
rect 291988 5216 291994 5228
rect 458266 5216 458272 5228
rect 291988 5188 458272 5216
rect 291988 5176 291994 5188
rect 458266 5176 458272 5188
rect 458324 5176 458330 5228
rect 107470 5108 107476 5160
rect 107528 5148 107534 5160
rect 312170 5148 312176 5160
rect 107528 5120 312176 5148
rect 107528 5108 107534 5120
rect 312170 5108 312176 5120
rect 312228 5108 312234 5160
rect 337102 5108 337108 5160
rect 337160 5148 337166 5160
rect 481634 5148 481640 5160
rect 337160 5120 481640 5148
rect 337160 5108 337166 5120
rect 481634 5108 481640 5120
rect 481692 5108 481698 5160
rect 114462 5040 114468 5092
rect 114520 5080 114526 5092
rect 187234 5080 187240 5092
rect 114520 5052 187240 5080
rect 114520 5040 114526 5052
rect 187234 5040 187240 5052
rect 187292 5040 187298 5092
rect 262214 5040 262220 5092
rect 262272 5080 262278 5092
rect 469214 5080 469220 5092
rect 262272 5052 469220 5080
rect 262272 5040 262278 5052
rect 469214 5040 469220 5052
rect 469272 5040 469278 5092
rect 118602 4972 118608 5024
rect 118660 5012 118666 5024
rect 205082 5012 205088 5024
rect 118660 4984 205088 5012
rect 118660 4972 118666 4984
rect 205082 4972 205088 4984
rect 205140 4972 205146 5024
rect 212350 4972 212356 5024
rect 212408 5012 212414 5024
rect 233694 5012 233700 5024
rect 212408 4984 233700 5012
rect 212408 4972 212414 4984
rect 233694 4972 233700 4984
rect 233752 4972 233758 5024
rect 251450 4972 251456 5024
rect 251508 5012 251514 5024
rect 469306 5012 469312 5024
rect 251508 4984 469312 5012
rect 251508 4972 251514 4984
rect 469306 4972 469312 4984
rect 469364 4972 469370 5024
rect 84838 4904 84844 4956
rect 84896 4944 84902 4956
rect 140866 4944 140872 4956
rect 84896 4916 140872 4944
rect 84896 4904 84902 4916
rect 140866 4904 140872 4916
rect 140924 4904 140930 4956
rect 144454 4904 144460 4956
rect 144512 4944 144518 4956
rect 374641 4947 374699 4953
rect 374641 4944 374653 4947
rect 144512 4916 374653 4944
rect 144512 4904 144518 4916
rect 374641 4913 374653 4916
rect 374687 4913 374699 4947
rect 374641 4907 374699 4913
rect 387794 4904 387800 4956
rect 387852 4944 387858 4956
rect 471238 4944 471244 4956
rect 387852 4916 471244 4944
rect 387852 4904 387858 4916
rect 471238 4904 471244 4916
rect 471296 4904 471302 4956
rect 101950 4836 101956 4888
rect 102008 4876 102014 4888
rect 426342 4876 426348 4888
rect 102008 4848 426348 4876
rect 102008 4836 102014 4848
rect 426342 4836 426348 4848
rect 426400 4836 426406 4888
rect 433242 4836 433248 4888
rect 433300 4876 433306 4888
rect 475102 4876 475108 4888
rect 433300 4848 475108 4876
rect 433300 4836 433306 4848
rect 475102 4836 475108 4848
rect 475160 4836 475166 4888
rect 81894 4768 81900 4820
rect 81952 4808 81958 4820
rect 522666 4808 522672 4820
rect 81952 4780 522672 4808
rect 81952 4768 81958 4780
rect 522666 4768 522672 4780
rect 522724 4768 522730 4820
rect 333606 4700 333612 4752
rect 333664 4740 333670 4752
rect 444374 4740 444380 4752
rect 333664 4712 444380 4740
rect 333664 4700 333670 4712
rect 444374 4700 444380 4712
rect 444432 4700 444438 4752
rect 351733 4675 351791 4681
rect 351733 4641 351745 4675
rect 351779 4672 351791 4675
rect 362126 4672 362132 4684
rect 351779 4644 362132 4672
rect 351779 4641 351791 4644
rect 351733 4635 351791 4641
rect 362126 4632 362132 4644
rect 362184 4632 362190 4684
rect 374641 4675 374699 4681
rect 374641 4641 374653 4675
rect 374687 4672 374699 4675
rect 385034 4672 385040 4684
rect 374687 4644 385040 4672
rect 374687 4641 374699 4644
rect 374641 4635 374699 4641
rect 385034 4632 385040 4644
rect 385092 4632 385098 4684
rect 408494 4632 408500 4684
rect 408552 4672 408558 4684
rect 455414 4672 455420 4684
rect 408552 4644 455420 4672
rect 408552 4632 408558 4644
rect 455414 4632 455420 4644
rect 455472 4632 455478 4684
rect 379974 4564 379980 4616
rect 380032 4604 380038 4616
rect 419626 4604 419632 4616
rect 380032 4576 419632 4604
rect 380032 4564 380038 4576
rect 419626 4564 419632 4576
rect 419684 4564 419690 4616
rect 494977 4335 495035 4341
rect 494977 4301 494989 4335
rect 495023 4332 495035 4335
rect 500126 4332 500132 4344
rect 495023 4304 500132 4332
rect 495023 4301 495035 4304
rect 494977 4295 495035 4301
rect 500126 4292 500132 4304
rect 500184 4292 500190 4344
rect 494698 4224 494704 4276
rect 494756 4264 494762 4276
rect 495618 4264 495624 4276
rect 494756 4236 495624 4264
rect 494756 4224 494762 4236
rect 495618 4224 495624 4236
rect 495676 4224 495682 4276
rect 94409 4199 94467 4205
rect 94409 4165 94421 4199
rect 94455 4196 94467 4199
rect 99285 4199 99343 4205
rect 99285 4196 99297 4199
rect 94455 4168 94636 4196
rect 94455 4165 94467 4168
rect 94409 4159 94467 4165
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 9030 4128 9036 4140
rect 624 4100 9036 4128
rect 624 4088 630 4100
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 32674 4088 32680 4140
rect 32732 4128 32738 4140
rect 51718 4128 51724 4140
rect 32732 4100 51724 4128
rect 32732 4088 32738 4100
rect 51718 4088 51724 4100
rect 51776 4088 51782 4140
rect 76650 4088 76656 4140
rect 76708 4128 76714 4140
rect 77110 4128 77116 4140
rect 76708 4100 77116 4128
rect 76708 4088 76714 4100
rect 77110 4088 77116 4100
rect 77168 4088 77174 4140
rect 84930 4088 84936 4140
rect 84988 4128 84994 4140
rect 85482 4128 85488 4140
rect 84988 4100 85488 4128
rect 84988 4088 84994 4100
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 87322 4088 87328 4140
rect 87380 4128 87386 4140
rect 88242 4128 88248 4140
rect 87380 4100 88248 4128
rect 87380 4088 87386 4100
rect 88242 4088 88248 4100
rect 88300 4088 88306 4140
rect 88337 4131 88395 4137
rect 88337 4097 88349 4131
rect 88383 4128 88395 4131
rect 94501 4131 94559 4137
rect 94501 4128 94513 4131
rect 88383 4100 94513 4128
rect 88383 4097 88395 4100
rect 88337 4091 88395 4097
rect 94501 4097 94513 4100
rect 94547 4097 94559 4131
rect 94608 4128 94636 4168
rect 95620 4168 96660 4196
rect 95620 4128 95648 4168
rect 94608 4100 95648 4128
rect 94501 4091 94559 4097
rect 95694 4088 95700 4140
rect 95752 4128 95758 4140
rect 96522 4128 96528 4140
rect 95752 4100 96528 4128
rect 95752 4088 95758 4100
rect 96522 4088 96528 4100
rect 96580 4088 96586 4140
rect 96632 4128 96660 4168
rect 98012 4168 99297 4196
rect 98012 4128 98040 4168
rect 99285 4165 99297 4168
rect 99331 4165 99343 4199
rect 99285 4159 99343 4165
rect 112257 4199 112315 4205
rect 112257 4165 112269 4199
rect 112303 4196 112315 4199
rect 118329 4199 118387 4205
rect 118329 4196 118341 4199
rect 112303 4168 118341 4196
rect 112303 4165 112315 4168
rect 112257 4159 112315 4165
rect 118329 4165 118341 4168
rect 118375 4165 118387 4199
rect 118329 4159 118387 4165
rect 162946 4156 162952 4208
rect 163004 4196 163010 4208
rect 164694 4196 164700 4208
rect 163004 4168 164700 4196
rect 163004 4156 163010 4168
rect 164694 4156 164700 4168
rect 164752 4156 164758 4208
rect 405642 4156 405648 4208
rect 405700 4196 405706 4208
rect 413830 4196 413836 4208
rect 405700 4168 413836 4196
rect 405700 4156 405706 4168
rect 413830 4156 413836 4168
rect 413888 4156 413894 4208
rect 414014 4156 414020 4208
rect 414072 4196 414078 4208
rect 424962 4196 424968 4208
rect 414072 4168 424968 4196
rect 414072 4156 414078 4168
rect 424962 4156 424968 4168
rect 425020 4156 425026 4208
rect 495066 4156 495072 4208
rect 495124 4196 495130 4208
rect 495526 4196 495532 4208
rect 495124 4168 495532 4196
rect 495124 4156 495130 4168
rect 495526 4156 495532 4168
rect 495584 4156 495590 4208
rect 500052 4168 501000 4196
rect 96632 4100 98040 4128
rect 98086 4088 98092 4140
rect 98144 4128 98150 4140
rect 99098 4128 99104 4140
rect 98144 4100 99104 4128
rect 98144 4088 98150 4100
rect 99098 4088 99104 4100
rect 99156 4088 99162 4140
rect 99193 4131 99251 4137
rect 99193 4097 99205 4131
rect 99239 4128 99251 4131
rect 352558 4128 352564 4140
rect 99239 4100 352564 4128
rect 99239 4097 99251 4100
rect 99193 4091 99251 4097
rect 352558 4088 352564 4100
rect 352616 4088 352622 4140
rect 354950 4088 354956 4140
rect 355008 4128 355014 4140
rect 355962 4128 355968 4140
rect 355008 4100 355968 4128
rect 355008 4088 355014 4100
rect 355962 4088 355968 4100
rect 356020 4088 356026 4140
rect 364518 4088 364524 4140
rect 364576 4128 364582 4140
rect 365622 4128 365628 4140
rect 364576 4100 365628 4128
rect 364576 4088 364582 4100
rect 365622 4088 365628 4100
rect 365680 4088 365686 4140
rect 365714 4088 365720 4140
rect 365772 4128 365778 4140
rect 367002 4128 367008 4140
rect 365772 4100 367008 4128
rect 365772 4088 365778 4100
rect 367002 4088 367008 4100
rect 367060 4088 367066 4140
rect 373994 4088 374000 4140
rect 374052 4128 374058 4140
rect 375190 4128 375196 4140
rect 374052 4100 375196 4128
rect 374052 4088 374058 4100
rect 375190 4088 375196 4100
rect 375248 4088 375254 4140
rect 381170 4088 381176 4140
rect 381228 4128 381234 4140
rect 500052 4128 500080 4168
rect 381228 4100 500080 4128
rect 381228 4088 381234 4100
rect 500126 4088 500132 4140
rect 500184 4128 500190 4140
rect 500862 4128 500868 4140
rect 500184 4100 500868 4128
rect 500184 4088 500190 4100
rect 500862 4088 500868 4100
rect 500920 4088 500926 4140
rect 500972 4128 501000 4168
rect 501598 4128 501604 4140
rect 500972 4100 501604 4128
rect 501598 4088 501604 4100
rect 501656 4088 501662 4140
rect 502518 4088 502524 4140
rect 502576 4128 502582 4140
rect 503622 4128 503628 4140
rect 502576 4100 503628 4128
rect 502576 4088 502582 4100
rect 503622 4088 503628 4100
rect 503680 4088 503686 4140
rect 507670 4088 507676 4140
rect 507728 4128 507734 4140
rect 508406 4128 508412 4140
rect 507728 4100 508412 4128
rect 507728 4088 507734 4100
rect 508406 4088 508412 4100
rect 508464 4088 508470 4140
rect 511258 4088 511264 4140
rect 511316 4128 511322 4140
rect 511994 4128 512000 4140
rect 511316 4100 512000 4128
rect 511316 4088 511322 4100
rect 511994 4088 512000 4100
rect 512052 4088 512058 4140
rect 42150 4020 42156 4072
rect 42208 4060 42214 4072
rect 64138 4060 64144 4072
rect 42208 4032 64144 4060
rect 42208 4020 42214 4032
rect 64138 4020 64144 4032
rect 64196 4020 64202 4072
rect 76742 4020 76748 4072
rect 76800 4060 76806 4072
rect 340690 4060 340696 4072
rect 76800 4032 340696 4060
rect 76800 4020 76806 4032
rect 340690 4020 340696 4032
rect 340748 4020 340754 4072
rect 347866 4020 347872 4072
rect 347924 4060 347930 4072
rect 348970 4060 348976 4072
rect 347924 4032 348976 4060
rect 347924 4020 347930 4032
rect 348970 4020 348976 4032
rect 349028 4020 349034 4072
rect 349065 4063 349123 4069
rect 349065 4029 349077 4063
rect 349111 4060 349123 4063
rect 509326 4060 509332 4072
rect 349111 4032 509332 4060
rect 349111 4029 349123 4032
rect 349065 4023 349123 4029
rect 509326 4020 509332 4032
rect 509384 4020 509390 4072
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 304997 3995 305055 4001
rect 304997 3992 305009 3995
rect 43404 3964 305009 3992
rect 43404 3952 43410 3964
rect 304997 3961 305009 3964
rect 305043 3961 305055 3995
rect 304997 3955 305055 3961
rect 326341 3995 326399 4001
rect 326341 3961 326353 3995
rect 326387 3992 326399 3995
rect 506566 3992 506572 4004
rect 326387 3964 506572 3992
rect 326387 3961 326399 3964
rect 326341 3955 326399 3961
rect 506566 3952 506572 3964
rect 506624 3952 506630 4004
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 51810 3924 51816 3936
rect 30340 3896 51816 3924
rect 30340 3884 30346 3896
rect 51810 3884 51816 3896
rect 51868 3884 51874 3936
rect 52822 3884 52828 3936
rect 52880 3924 52886 3936
rect 57238 3924 57244 3936
rect 52880 3896 57244 3924
rect 52880 3884 52886 3896
rect 57238 3884 57244 3896
rect 57296 3884 57302 3936
rect 76834 3884 76840 3936
rect 76892 3924 76898 3936
rect 351362 3924 351368 3936
rect 76892 3896 351368 3924
rect 76892 3884 76898 3896
rect 351362 3884 351368 3896
rect 351420 3884 351426 3936
rect 385862 3884 385868 3936
rect 385920 3924 385926 3936
rect 506474 3924 506480 3936
rect 385920 3896 506480 3924
rect 385920 3884 385926 3896
rect 506474 3884 506480 3896
rect 506532 3884 506538 3936
rect 26694 3816 26700 3868
rect 26752 3856 26758 3868
rect 50338 3856 50344 3868
rect 26752 3828 50344 3856
rect 26752 3816 26758 3828
rect 50338 3816 50344 3828
rect 50396 3816 50402 3868
rect 80422 3816 80428 3868
rect 80480 3856 80486 3868
rect 208581 3859 208639 3865
rect 208581 3856 208593 3859
rect 80480 3828 208593 3856
rect 80480 3816 80486 3828
rect 208581 3825 208593 3828
rect 208627 3825 208639 3859
rect 208581 3819 208639 3825
rect 208670 3816 208676 3868
rect 208728 3856 208734 3868
rect 209682 3856 209688 3868
rect 208728 3828 209688 3856
rect 208728 3816 208734 3828
rect 209682 3816 209688 3828
rect 209740 3816 209746 3868
rect 209866 3816 209872 3868
rect 209924 3856 209930 3868
rect 210970 3856 210976 3868
rect 209924 3828 210976 3856
rect 209924 3816 209930 3828
rect 210970 3816 210976 3828
rect 211028 3816 211034 3868
rect 215846 3816 215852 3868
rect 215904 3856 215910 3868
rect 216582 3856 216588 3868
rect 215904 3828 216588 3856
rect 215904 3816 215910 3828
rect 216582 3816 216588 3828
rect 216640 3816 216646 3868
rect 217042 3816 217048 3868
rect 217100 3856 217106 3868
rect 217962 3856 217968 3868
rect 217100 3828 217968 3856
rect 217100 3816 217106 3828
rect 217962 3816 217968 3828
rect 218020 3816 218026 3868
rect 226518 3816 226524 3868
rect 226576 3856 226582 3868
rect 227622 3856 227628 3868
rect 226576 3828 227628 3856
rect 226576 3816 226582 3828
rect 227622 3816 227628 3828
rect 227680 3816 227686 3868
rect 227714 3816 227720 3868
rect 227772 3856 227778 3868
rect 498841 3859 498899 3865
rect 498841 3856 498853 3859
rect 227772 3828 498853 3856
rect 227772 3816 227778 3828
rect 498841 3825 498853 3828
rect 498887 3825 498899 3859
rect 498841 3819 498899 3825
rect 498930 3816 498936 3868
rect 498988 3856 498994 3868
rect 501690 3856 501696 3868
rect 498988 3828 501696 3856
rect 498988 3816 498994 3828
rect 501690 3816 501696 3828
rect 501748 3816 501754 3868
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 31018 3788 31024 3800
rect 25556 3760 31024 3788
rect 25556 3748 25562 3760
rect 31018 3748 31024 3760
rect 31076 3748 31082 3800
rect 39758 3748 39764 3800
rect 39816 3788 39822 3800
rect 313918 3788 313924 3800
rect 39816 3760 313924 3788
rect 39816 3748 39822 3760
rect 313918 3748 313924 3760
rect 313976 3748 313982 3800
rect 315758 3748 315764 3800
rect 315816 3788 315822 3800
rect 502242 3788 502248 3800
rect 315816 3760 502248 3788
rect 315816 3748 315822 3760
rect 502242 3748 502248 3760
rect 502300 3748 502306 3800
rect 538858 3748 538864 3800
rect 538916 3788 538922 3800
rect 548886 3788 548892 3800
rect 538916 3760 548892 3788
rect 538916 3748 538922 3760
rect 548886 3748 548892 3760
rect 548944 3748 548950 3800
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 59998 3720 60004 3732
rect 31536 3692 60004 3720
rect 31536 3680 31542 3692
rect 59998 3680 60004 3692
rect 60056 3680 60062 3732
rect 69293 3723 69351 3729
rect 69293 3689 69305 3723
rect 69339 3720 69351 3723
rect 73798 3720 73804 3732
rect 69339 3692 73804 3720
rect 69339 3689 69351 3692
rect 69293 3683 69351 3689
rect 73798 3680 73804 3692
rect 73856 3680 73862 3732
rect 89714 3680 89720 3732
rect 89772 3720 89778 3732
rect 91002 3720 91008 3732
rect 89772 3692 91008 3720
rect 89772 3680 89778 3692
rect 91002 3680 91008 3692
rect 91060 3680 91066 3732
rect 93302 3680 93308 3732
rect 93360 3720 93366 3732
rect 99193 3723 99251 3729
rect 99193 3720 99205 3723
rect 93360 3692 99205 3720
rect 93360 3680 93366 3692
rect 99193 3689 99205 3692
rect 99239 3689 99251 3723
rect 99193 3683 99251 3689
rect 101582 3680 101588 3732
rect 101640 3720 101646 3732
rect 102042 3720 102048 3732
rect 101640 3692 102048 3720
rect 101640 3680 101646 3692
rect 102042 3680 102048 3692
rect 102100 3680 102106 3732
rect 103514 3680 103520 3732
rect 103572 3720 103578 3732
rect 103974 3720 103980 3732
rect 103572 3692 103980 3720
rect 103572 3680 103578 3692
rect 103974 3680 103980 3692
rect 104032 3680 104038 3732
rect 105170 3680 105176 3732
rect 105228 3720 105234 3732
rect 106182 3720 106188 3732
rect 105228 3692 106188 3720
rect 105228 3680 105234 3692
rect 106182 3680 106188 3692
rect 106240 3680 106246 3732
rect 106366 3680 106372 3732
rect 106424 3720 106430 3732
rect 107562 3720 107568 3732
rect 106424 3692 107568 3720
rect 106424 3680 106430 3692
rect 107562 3680 107568 3692
rect 107620 3680 107626 3732
rect 109037 3723 109095 3729
rect 109037 3689 109049 3723
rect 109083 3720 109095 3723
rect 112257 3723 112315 3729
rect 112257 3720 112269 3723
rect 109083 3692 112269 3720
rect 109083 3689 109095 3692
rect 109037 3683 109095 3689
rect 112257 3689 112269 3692
rect 112303 3689 112315 3723
rect 112257 3683 112315 3689
rect 112346 3680 112352 3732
rect 112404 3720 112410 3732
rect 113082 3720 113088 3732
rect 112404 3692 113088 3720
rect 112404 3680 112410 3692
rect 113082 3680 113088 3692
rect 113140 3680 113146 3732
rect 115750 3680 115756 3732
rect 115808 3720 115814 3732
rect 116854 3720 116860 3732
rect 115808 3692 116860 3720
rect 115808 3680 115814 3692
rect 116854 3680 116860 3692
rect 116912 3680 116918 3732
rect 118329 3723 118387 3729
rect 118329 3689 118341 3723
rect 118375 3720 118387 3723
rect 393314 3720 393320 3732
rect 118375 3692 393320 3720
rect 118375 3689 118387 3692
rect 118329 3683 118387 3689
rect 393314 3680 393320 3692
rect 393372 3680 393378 3732
rect 393866 3680 393872 3732
rect 393924 3720 393930 3732
rect 567838 3720 567844 3732
rect 393924 3692 567844 3720
rect 393924 3680 393930 3692
rect 567838 3680 567844 3692
rect 567896 3680 567902 3732
rect 29086 3612 29092 3664
rect 29144 3652 29150 3664
rect 42058 3652 42064 3664
rect 29144 3624 42064 3652
rect 29144 3612 29150 3624
rect 42058 3612 42064 3624
rect 42116 3612 42122 3664
rect 45738 3612 45744 3664
rect 45796 3652 45802 3664
rect 393961 3655 394019 3661
rect 393961 3652 393973 3655
rect 45796 3624 393973 3652
rect 45796 3612 45802 3624
rect 393961 3621 393973 3624
rect 394007 3621 394019 3655
rect 393961 3615 394019 3621
rect 397822 3612 397828 3664
rect 397880 3652 397886 3664
rect 398742 3652 398748 3664
rect 397880 3624 398748 3652
rect 397880 3612 397886 3624
rect 398742 3612 398748 3624
rect 398800 3612 398806 3664
rect 399018 3612 399024 3664
rect 399076 3652 399082 3664
rect 400122 3652 400128 3664
rect 399076 3624 400128 3652
rect 399076 3612 399082 3624
rect 400122 3612 400128 3624
rect 400180 3612 400186 3664
rect 406102 3612 406108 3664
rect 406160 3652 406166 3664
rect 407022 3652 407028 3664
rect 406160 3624 407028 3652
rect 406160 3612 406166 3624
rect 407022 3612 407028 3624
rect 407080 3612 407086 3664
rect 412082 3612 412088 3664
rect 412140 3652 412146 3664
rect 415486 3652 415492 3664
rect 412140 3624 415492 3652
rect 412140 3612 412146 3624
rect 415486 3612 415492 3624
rect 415544 3612 415550 3664
rect 415581 3655 415639 3661
rect 415581 3621 415593 3655
rect 415627 3652 415639 3655
rect 430117 3655 430175 3661
rect 430117 3652 430129 3655
rect 415627 3624 430129 3652
rect 415627 3621 415639 3624
rect 415581 3615 415639 3621
rect 430117 3621 430129 3624
rect 430163 3621 430175 3655
rect 430117 3615 430175 3621
rect 431126 3612 431132 3664
rect 431184 3652 431190 3664
rect 431862 3652 431868 3664
rect 431184 3624 431868 3652
rect 431184 3612 431190 3624
rect 431862 3612 431868 3624
rect 431920 3612 431926 3664
rect 439406 3612 439412 3664
rect 439464 3652 439470 3664
rect 440142 3652 440148 3664
rect 439464 3624 440148 3652
rect 439464 3612 439470 3624
rect 440142 3612 440148 3624
rect 440200 3612 440206 3664
rect 444190 3612 444196 3664
rect 444248 3652 444254 3664
rect 500221 3655 500279 3661
rect 500221 3652 500233 3655
rect 444248 3624 500233 3652
rect 444248 3612 444254 3624
rect 500221 3621 500233 3624
rect 500267 3621 500279 3655
rect 500221 3615 500279 3621
rect 519630 3612 519636 3664
rect 519688 3652 519694 3664
rect 528646 3652 528652 3664
rect 519688 3624 528652 3652
rect 519688 3612 519694 3624
rect 528646 3612 528652 3624
rect 528704 3612 528710 3664
rect 531958 3612 531964 3664
rect 532016 3652 532022 3664
rect 532016 3624 532464 3652
rect 532016 3612 532022 3624
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 46290 3584 46296 3596
rect 17368 3556 46296 3584
rect 17368 3544 17374 3556
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 53098 3584 53104 3596
rect 46860 3556 53104 3584
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4798 3516 4804 3528
rect 2924 3488 4804 3516
rect 2924 3476 2930 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 12342 3516 12348 3528
rect 11296 3488 12348 3516
rect 11296 3476 11302 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 17218 3516 17224 3528
rect 12452 3488 17224 3516
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 12452 3448 12480 3488
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20622 3516 20628 3528
rect 19576 3488 20628 3516
rect 19576 3476 19582 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 46860 3516 46888 3556
rect 53098 3544 53104 3556
rect 53156 3544 53162 3596
rect 55214 3544 55220 3596
rect 55272 3584 55278 3596
rect 56410 3584 56416 3596
rect 55272 3556 56416 3584
rect 55272 3544 55278 3556
rect 56410 3544 56416 3556
rect 56468 3544 56474 3596
rect 59998 3544 60004 3596
rect 60056 3584 60062 3596
rect 71038 3584 71044 3596
rect 60056 3556 71044 3584
rect 60056 3544 60062 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 77662 3544 77668 3596
rect 77720 3584 77726 3596
rect 504818 3584 504824 3596
rect 77720 3556 504824 3584
rect 77720 3544 77726 3556
rect 504818 3544 504824 3556
rect 504876 3544 504882 3596
rect 522298 3544 522304 3596
rect 522356 3584 522362 3596
rect 532234 3584 532240 3596
rect 522356 3556 532240 3584
rect 522356 3544 522362 3556
rect 532234 3544 532240 3556
rect 532292 3544 532298 3596
rect 532436 3584 532464 3624
rect 540330 3612 540336 3664
rect 540388 3652 540394 3664
rect 582190 3652 582196 3664
rect 540388 3624 582196 3652
rect 540388 3612 540394 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 532436 3556 571380 3584
rect 23164 3488 46888 3516
rect 23164 3476 23170 3488
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 48958 3516 48964 3528
rect 46992 3488 48964 3516
rect 46992 3476 46998 3488
rect 48958 3476 48964 3488
rect 49016 3476 49022 3528
rect 51626 3476 51632 3528
rect 51684 3516 51690 3528
rect 52362 3516 52368 3528
rect 51684 3488 52368 3516
rect 51684 3476 51690 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 58802 3476 58808 3528
rect 58860 3516 58866 3528
rect 59262 3516 59268 3528
rect 58860 3488 59268 3516
rect 58860 3476 58866 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 61378 3516 61384 3528
rect 59372 3488 61384 3516
rect 8904 3420 12480 3448
rect 8904 3408 8910 3420
rect 24302 3408 24308 3460
rect 24360 3448 24366 3460
rect 59372 3448 59400 3488
rect 61378 3476 61384 3488
rect 61436 3476 61442 3528
rect 62390 3476 62396 3528
rect 62448 3516 62454 3528
rect 63402 3516 63408 3528
rect 62448 3488 63408 3516
rect 62448 3476 62454 3488
rect 63402 3476 63408 3488
rect 63460 3476 63466 3528
rect 63586 3476 63592 3528
rect 63644 3516 63650 3528
rect 64690 3516 64696 3528
rect 63644 3488 64696 3516
rect 63644 3476 63650 3488
rect 64690 3476 64696 3488
rect 64748 3476 64754 3528
rect 69293 3519 69351 3525
rect 69293 3516 69305 3519
rect 64800 3488 69305 3516
rect 24360 3420 59400 3448
rect 24360 3408 24366 3420
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 35802 3380 35808 3392
rect 35032 3352 35808 3380
rect 35032 3340 35038 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 38470 3380 38476 3392
rect 37424 3352 38476 3380
rect 37424 3340 37430 3352
rect 38470 3340 38476 3352
rect 38528 3340 38534 3392
rect 46198 3380 46204 3392
rect 38580 3352 46204 3380
rect 1670 3272 1676 3324
rect 1728 3312 1734 3324
rect 1728 3284 7604 3312
rect 1728 3272 1734 3284
rect 7576 3244 7604 3284
rect 7650 3272 7656 3324
rect 7708 3312 7714 3324
rect 9122 3312 9128 3324
rect 7708 3284 9128 3312
rect 7708 3272 7714 3284
rect 9122 3272 9128 3284
rect 9180 3272 9186 3324
rect 36170 3272 36176 3324
rect 36228 3312 36234 3324
rect 38580 3312 38608 3352
rect 46198 3340 46204 3352
rect 46256 3340 46262 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 64800 3380 64828 3488
rect 69293 3485 69305 3488
rect 69339 3485 69351 3519
rect 69293 3479 69351 3485
rect 69474 3476 69480 3528
rect 69532 3516 69538 3528
rect 70210 3516 70216 3528
rect 69532 3488 70216 3516
rect 69532 3476 69538 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 70670 3476 70676 3528
rect 70728 3516 70734 3528
rect 71682 3516 71688 3528
rect 70728 3488 71688 3516
rect 70728 3476 70734 3488
rect 71682 3476 71688 3488
rect 71740 3476 71746 3528
rect 71866 3476 71872 3528
rect 71924 3516 71930 3528
rect 72970 3516 72976 3528
rect 71924 3488 72976 3516
rect 71924 3476 71930 3488
rect 72970 3476 72976 3488
rect 73028 3476 73034 3528
rect 77478 3476 77484 3528
rect 77536 3516 77542 3528
rect 554774 3516 554780 3528
rect 77536 3488 554780 3516
rect 77536 3476 77542 3488
rect 554774 3476 554780 3488
rect 554832 3476 554838 3528
rect 77570 3408 77576 3460
rect 77628 3448 77634 3460
rect 569034 3448 569040 3460
rect 77628 3420 569040 3448
rect 77628 3408 77634 3420
rect 569034 3408 569040 3420
rect 569092 3408 569098 3460
rect 571352 3448 571380 3556
rect 571426 3544 571432 3596
rect 571484 3584 571490 3596
rect 572622 3584 572628 3596
rect 571484 3556 572628 3584
rect 571484 3544 571490 3556
rect 572622 3544 572628 3556
rect 572680 3544 572686 3596
rect 576210 3448 576216 3460
rect 571352 3420 576216 3448
rect 576210 3408 576216 3420
rect 576268 3408 576274 3460
rect 61252 3352 64828 3380
rect 61252 3340 61258 3352
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 209501 3383 209559 3389
rect 209501 3380 209513 3383
rect 68336 3352 209513 3380
rect 68336 3340 68342 3352
rect 209501 3349 209513 3352
rect 209547 3349 209559 3383
rect 209501 3343 209559 3349
rect 219529 3383 219587 3389
rect 219529 3349 219541 3383
rect 219575 3380 219587 3383
rect 249061 3383 249119 3389
rect 249061 3380 249073 3383
rect 219575 3352 249073 3380
rect 219575 3349 219587 3352
rect 219529 3343 219587 3349
rect 249061 3349 249073 3352
rect 249107 3349 249119 3383
rect 249061 3343 249119 3349
rect 249150 3340 249156 3392
rect 249208 3380 249214 3392
rect 249702 3380 249708 3392
rect 249208 3352 249708 3380
rect 249208 3340 249214 3352
rect 249702 3340 249708 3352
rect 249760 3340 249766 3392
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 251082 3380 251088 3392
rect 250404 3352 251088 3380
rect 250404 3340 250410 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 252646 3340 252652 3392
rect 252704 3380 252710 3392
rect 253842 3380 253848 3392
rect 252704 3352 253848 3380
rect 252704 3340 252710 3352
rect 253842 3340 253848 3352
rect 253900 3340 253906 3392
rect 258721 3383 258779 3389
rect 258721 3349 258733 3383
rect 258767 3380 258779 3383
rect 283561 3383 283619 3389
rect 283561 3380 283573 3383
rect 258767 3352 283573 3380
rect 258767 3349 258779 3352
rect 258721 3343 258779 3349
rect 283561 3349 283573 3352
rect 283607 3349 283619 3383
rect 283561 3343 283619 3349
rect 283650 3340 283656 3392
rect 283708 3380 283714 3392
rect 284202 3380 284208 3392
rect 283708 3352 284208 3380
rect 283708 3340 283714 3352
rect 284202 3340 284208 3352
rect 284260 3340 284266 3392
rect 285950 3340 285956 3392
rect 286008 3380 286014 3392
rect 286962 3380 286968 3392
rect 286008 3352 286968 3380
rect 286008 3340 286014 3352
rect 286962 3340 286968 3352
rect 287020 3340 287026 3392
rect 293126 3340 293132 3392
rect 293184 3380 293190 3392
rect 293862 3380 293868 3392
rect 293184 3352 293868 3380
rect 293184 3340 293190 3352
rect 293862 3340 293868 3352
rect 293920 3340 293926 3392
rect 295518 3340 295524 3392
rect 295576 3380 295582 3392
rect 296622 3380 296628 3392
rect 295576 3352 296628 3380
rect 295576 3340 295582 3352
rect 296622 3340 296628 3352
rect 296680 3340 296686 3392
rect 303798 3340 303804 3392
rect 303856 3380 303862 3392
rect 304902 3380 304908 3392
rect 303856 3352 304908 3380
rect 303856 3340 303862 3352
rect 304902 3340 304908 3352
rect 304960 3340 304966 3392
rect 304997 3383 305055 3389
rect 304997 3349 305009 3383
rect 305043 3380 305055 3383
rect 307754 3380 307760 3392
rect 305043 3352 307760 3380
rect 305043 3349 305055 3352
rect 304997 3343 305055 3349
rect 307754 3340 307760 3352
rect 307812 3340 307818 3392
rect 321646 3340 321652 3392
rect 321704 3380 321710 3392
rect 322750 3380 322756 3392
rect 321704 3352 322756 3380
rect 321704 3340 321710 3352
rect 322750 3340 322756 3352
rect 322808 3340 322814 3392
rect 324038 3340 324044 3392
rect 324096 3380 324102 3392
rect 326341 3383 326399 3389
rect 326341 3380 326353 3383
rect 324096 3352 326353 3380
rect 324096 3340 324102 3352
rect 326341 3349 326353 3352
rect 326387 3349 326399 3383
rect 326341 3343 326399 3349
rect 326430 3340 326436 3392
rect 326488 3380 326494 3392
rect 326982 3380 326988 3392
rect 326488 3352 326988 3380
rect 326488 3340 326494 3352
rect 326982 3340 326988 3352
rect 327040 3340 327046 3392
rect 327626 3340 327632 3392
rect 327684 3380 327690 3392
rect 328362 3380 328368 3392
rect 327684 3352 328368 3380
rect 327684 3340 327690 3352
rect 328362 3340 328368 3352
rect 328420 3340 328426 3392
rect 328822 3340 328828 3392
rect 328880 3380 328886 3392
rect 329742 3380 329748 3392
rect 328880 3352 329748 3380
rect 328880 3340 328886 3352
rect 329742 3340 329748 3352
rect 329800 3340 329806 3392
rect 330018 3340 330024 3392
rect 330076 3380 330082 3392
rect 331122 3380 331128 3392
rect 330076 3352 331128 3380
rect 330076 3340 330082 3352
rect 331122 3340 331128 3352
rect 331180 3340 331186 3392
rect 331214 3340 331220 3392
rect 331272 3380 331278 3392
rect 332502 3380 332508 3392
rect 331272 3352 332508 3380
rect 331272 3340 331278 3352
rect 332502 3340 332508 3352
rect 332560 3340 332566 3392
rect 339494 3340 339500 3392
rect 339552 3380 339558 3392
rect 340782 3380 340788 3392
rect 339552 3352 340788 3380
rect 339552 3340 339558 3352
rect 340782 3340 340788 3352
rect 340840 3340 340846 3392
rect 344278 3340 344284 3392
rect 344336 3380 344342 3392
rect 349065 3383 349123 3389
rect 349065 3380 349077 3383
rect 344336 3352 349077 3380
rect 344336 3340 344342 3352
rect 349065 3349 349077 3352
rect 349111 3349 349123 3383
rect 349065 3343 349123 3349
rect 388254 3340 388260 3392
rect 388312 3380 388318 3392
rect 490653 3383 490711 3389
rect 490653 3380 490665 3383
rect 388312 3352 490665 3380
rect 388312 3340 388318 3352
rect 490653 3349 490665 3352
rect 490699 3349 490711 3383
rect 490653 3343 490711 3349
rect 500221 3383 500279 3389
rect 500221 3349 500233 3383
rect 500267 3380 500279 3383
rect 505094 3380 505100 3392
rect 500267 3352 505100 3380
rect 500267 3349 500279 3352
rect 500221 3343 500279 3349
rect 505094 3340 505100 3352
rect 505152 3340 505158 3392
rect 36228 3284 38608 3312
rect 36228 3272 36234 3284
rect 54018 3272 54024 3324
rect 54076 3312 54082 3324
rect 291286 3312 291292 3324
rect 54076 3284 291292 3312
rect 54076 3272 54082 3284
rect 291286 3272 291292 3284
rect 291344 3272 291350 3324
rect 297361 3315 297419 3321
rect 297361 3281 297373 3315
rect 297407 3312 297419 3315
rect 307018 3312 307024 3324
rect 297407 3284 307024 3312
rect 297407 3281 297419 3284
rect 297361 3275 297419 3281
rect 307018 3272 307024 3284
rect 307076 3272 307082 3324
rect 307386 3272 307392 3324
rect 307444 3312 307450 3324
rect 493318 3312 493324 3324
rect 307444 3284 493324 3312
rect 307444 3272 307450 3284
rect 493318 3272 493324 3284
rect 493376 3272 493382 3324
rect 494146 3272 494152 3324
rect 494204 3312 494210 3324
rect 494204 3284 503208 3312
rect 494204 3272 494210 3284
rect 9214 3244 9220 3256
rect 7576 3216 9220 3244
rect 9214 3204 9220 3216
rect 9272 3204 9278 3256
rect 77386 3204 77392 3256
rect 77444 3244 77450 3256
rect 248969 3247 249027 3253
rect 248969 3244 248981 3247
rect 77444 3216 214788 3244
rect 77444 3204 77450 3216
rect 65978 3136 65984 3188
rect 66036 3176 66042 3188
rect 69658 3176 69664 3188
rect 66036 3148 69664 3176
rect 66036 3136 66042 3148
rect 69658 3136 69664 3148
rect 69716 3136 69722 3188
rect 78122 3136 78128 3188
rect 78180 3176 78186 3188
rect 208489 3179 208547 3185
rect 208489 3176 208501 3179
rect 78180 3148 208501 3176
rect 78180 3136 78186 3148
rect 208489 3145 208501 3148
rect 208535 3145 208547 3179
rect 208489 3139 208547 3145
rect 208581 3179 208639 3185
rect 208581 3145 208593 3179
rect 208627 3176 208639 3179
rect 214650 3176 214656 3188
rect 208627 3148 214656 3176
rect 208627 3145 208639 3148
rect 208581 3139 208639 3145
rect 214650 3136 214656 3148
rect 214708 3136 214714 3188
rect 214760 3176 214788 3216
rect 220004 3216 248981 3244
rect 220004 3176 220032 3216
rect 248969 3213 248981 3216
rect 249015 3213 249027 3247
rect 248969 3207 249027 3213
rect 265802 3204 265808 3256
rect 265860 3244 265866 3256
rect 266262 3244 266268 3256
rect 265860 3216 266268 3244
rect 265860 3204 265866 3216
rect 266262 3204 266268 3216
rect 266320 3204 266326 3256
rect 266372 3216 269252 3244
rect 214760 3148 220032 3176
rect 220081 3179 220139 3185
rect 220081 3145 220093 3179
rect 220127 3176 220139 3179
rect 220817 3179 220875 3185
rect 220817 3176 220829 3179
rect 220127 3148 220829 3176
rect 220127 3145 220139 3148
rect 220081 3139 220139 3145
rect 220817 3145 220829 3148
rect 220863 3145 220875 3179
rect 255038 3176 255044 3188
rect 220817 3139 220875 3145
rect 246316 3148 255044 3176
rect 74258 3068 74264 3120
rect 74316 3108 74322 3120
rect 75178 3108 75184 3120
rect 74316 3080 75184 3108
rect 74316 3068 74322 3080
rect 75178 3068 75184 3080
rect 75236 3068 75242 3120
rect 85022 3068 85028 3120
rect 85080 3108 85086 3120
rect 99285 3111 99343 3117
rect 85080 3080 88472 3108
rect 85080 3068 85086 3080
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 13722 3040 13728 3052
rect 12492 3012 13728 3040
rect 12492 3000 12498 3012
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 22002 3040 22008 3052
rect 20772 3012 22008 3040
rect 20772 3000 20778 3012
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 77202 3000 77208 3052
rect 77260 3040 77266 3052
rect 88337 3043 88395 3049
rect 88337 3040 88349 3043
rect 77260 3012 88349 3040
rect 77260 3000 77266 3012
rect 88337 3009 88349 3012
rect 88383 3009 88395 3043
rect 88444 3040 88472 3080
rect 99285 3077 99297 3111
rect 99331 3108 99343 3111
rect 118697 3111 118755 3117
rect 118697 3108 118709 3111
rect 99331 3080 118709 3108
rect 99331 3077 99343 3080
rect 99285 3071 99343 3077
rect 118697 3077 118709 3080
rect 118743 3077 118755 3111
rect 118697 3071 118755 3077
rect 129734 3068 129740 3120
rect 129792 3108 129798 3120
rect 130194 3108 130200 3120
rect 129792 3080 130200 3108
rect 129792 3068 129798 3080
rect 130194 3068 130200 3080
rect 130252 3068 130258 3120
rect 132405 3111 132463 3117
rect 132405 3077 132417 3111
rect 132451 3108 132463 3111
rect 133877 3111 133935 3117
rect 133877 3108 133889 3111
rect 132451 3080 133889 3108
rect 132451 3077 132463 3080
rect 132405 3071 132463 3077
rect 133877 3077 133889 3080
rect 133923 3077 133935 3111
rect 133877 3071 133935 3077
rect 136082 3068 136088 3120
rect 136140 3108 136146 3120
rect 136542 3108 136548 3120
rect 136140 3080 136548 3108
rect 136140 3068 136146 3080
rect 136542 3068 136548 3080
rect 136600 3068 136606 3120
rect 136652 3080 139624 3108
rect 94409 3043 94467 3049
rect 94409 3040 94421 3043
rect 88444 3012 94421 3040
rect 88337 3003 88395 3009
rect 94409 3009 94421 3012
rect 94455 3009 94467 3043
rect 94409 3003 94467 3009
rect 94501 3043 94559 3049
rect 94501 3009 94513 3043
rect 94547 3040 94559 3043
rect 122837 3043 122895 3049
rect 122837 3040 122849 3043
rect 94547 3012 122849 3040
rect 94547 3009 94559 3012
rect 94501 3003 94559 3009
rect 122837 3009 122849 3012
rect 122883 3009 122895 3043
rect 122837 3003 122895 3009
rect 122926 3000 122932 3052
rect 122984 3040 122990 3052
rect 128173 3043 128231 3049
rect 128173 3040 128185 3043
rect 122984 3012 128185 3040
rect 122984 3000 122990 3012
rect 128173 3009 128185 3012
rect 128219 3009 128231 3043
rect 128173 3003 128231 3009
rect 128449 3043 128507 3049
rect 128449 3009 128461 3043
rect 128495 3040 128507 3043
rect 136652 3040 136680 3080
rect 128495 3012 136680 3040
rect 136729 3043 136787 3049
rect 128495 3009 128507 3012
rect 128449 3003 128507 3009
rect 136729 3009 136741 3043
rect 136775 3040 136787 3043
rect 139596 3040 139624 3080
rect 139670 3068 139676 3120
rect 139728 3108 139734 3120
rect 140682 3108 140688 3120
rect 139728 3080 140688 3108
rect 139728 3068 139734 3080
rect 140682 3068 140688 3080
rect 140740 3068 140746 3120
rect 142154 3068 142160 3120
rect 142212 3108 142218 3120
rect 143258 3108 143264 3120
rect 142212 3080 143264 3108
rect 142212 3068 142218 3080
rect 143258 3068 143264 3080
rect 143316 3068 143322 3120
rect 145650 3068 145656 3120
rect 145708 3108 145714 3120
rect 146202 3108 146208 3120
rect 145708 3080 146208 3108
rect 145708 3068 145714 3080
rect 146202 3068 146208 3080
rect 146260 3068 146266 3120
rect 146386 3068 146392 3120
rect 146444 3108 146450 3120
rect 146846 3108 146852 3120
rect 146444 3080 146852 3108
rect 146444 3068 146450 3080
rect 146846 3068 146852 3080
rect 146904 3068 146910 3120
rect 153194 3068 153200 3120
rect 153252 3108 153258 3120
rect 153930 3108 153936 3120
rect 153252 3080 153936 3108
rect 153252 3068 153258 3080
rect 153930 3068 153936 3080
rect 153988 3068 153994 3120
rect 157245 3111 157303 3117
rect 157245 3077 157257 3111
rect 157291 3108 157303 3111
rect 157337 3111 157395 3117
rect 157337 3108 157349 3111
rect 157291 3080 157349 3108
rect 157291 3077 157303 3080
rect 157245 3071 157303 3077
rect 157337 3077 157349 3080
rect 157383 3077 157395 3111
rect 157337 3071 157395 3077
rect 166905 3111 166963 3117
rect 166905 3077 166917 3111
rect 166951 3108 166963 3111
rect 166951 3080 179276 3108
rect 166951 3077 166963 3080
rect 166905 3071 166963 3077
rect 154025 3043 154083 3049
rect 154025 3040 154037 3043
rect 136775 3012 139532 3040
rect 139596 3012 154037 3040
rect 136775 3009 136787 3012
rect 136729 3003 136787 3009
rect 77754 2932 77760 2984
rect 77812 2972 77818 2984
rect 99374 2972 99380 2984
rect 77812 2944 99380 2972
rect 77812 2932 77818 2944
rect 99374 2932 99380 2944
rect 99432 2932 99438 2984
rect 108942 2932 108948 2984
rect 109000 2972 109006 2984
rect 118694 2972 118700 2984
rect 109000 2944 118700 2972
rect 109000 2932 109006 2944
rect 118694 2932 118700 2944
rect 118752 2932 118758 2984
rect 118789 2975 118847 2981
rect 118789 2941 118801 2975
rect 118835 2972 118847 2975
rect 128265 2975 128323 2981
rect 128265 2972 128277 2975
rect 118835 2944 128277 2972
rect 118835 2941 118847 2944
rect 118789 2935 118847 2941
rect 128265 2941 128277 2944
rect 128311 2941 128323 2975
rect 128265 2935 128323 2941
rect 128357 2975 128415 2981
rect 128357 2941 128369 2975
rect 128403 2972 128415 2975
rect 139504 2972 139532 3012
rect 154025 3009 154037 3012
rect 154071 3009 154083 3043
rect 154025 3003 154083 3009
rect 154117 3043 154175 3049
rect 154117 3009 154129 3043
rect 154163 3040 154175 3043
rect 154163 3012 157472 3040
rect 154163 3009 154175 3012
rect 154117 3003 154175 3009
rect 142801 2975 142859 2981
rect 142801 2972 142813 2975
rect 128403 2944 139440 2972
rect 139504 2944 142813 2972
rect 128403 2941 128415 2944
rect 128357 2935 128415 2941
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 8938 2904 8944 2916
rect 4120 2876 8944 2904
rect 4120 2864 4126 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 85114 2864 85120 2916
rect 85172 2904 85178 2916
rect 139412 2904 139440 2944
rect 142801 2941 142813 2944
rect 142847 2941 142859 2975
rect 157444 2972 157472 3012
rect 157518 3000 157524 3052
rect 157576 3040 157582 3052
rect 158622 3040 158628 3052
rect 157576 3012 158628 3040
rect 157576 3000 157582 3012
rect 158622 3000 158628 3012
rect 158680 3000 158686 3052
rect 164694 3000 164700 3052
rect 164752 3040 164758 3052
rect 165522 3040 165528 3052
rect 164752 3012 165528 3040
rect 164752 3000 164758 3012
rect 165522 3000 165528 3012
rect 165580 3000 165586 3052
rect 167178 3000 167184 3052
rect 167236 3040 167242 3052
rect 168190 3040 168196 3052
rect 167236 3012 168196 3040
rect 167236 3000 167242 3012
rect 168190 3000 168196 3012
rect 168248 3000 168254 3052
rect 172974 3000 172980 3052
rect 173032 3040 173038 3052
rect 173802 3040 173808 3052
rect 173032 3012 173808 3040
rect 173032 3000 173038 3012
rect 173802 3000 173808 3012
rect 173860 3000 173866 3052
rect 176654 3000 176660 3052
rect 176712 3040 176718 3052
rect 177758 3040 177764 3052
rect 176712 3012 177764 3040
rect 176712 3000 176718 3012
rect 177758 3000 177764 3012
rect 177816 3000 177822 3052
rect 165890 2972 165896 2984
rect 157444 2944 165896 2972
rect 142801 2935 142859 2941
rect 165890 2932 165896 2944
rect 165948 2932 165954 2984
rect 179248 2972 179276 3080
rect 179414 3068 179420 3120
rect 179472 3108 179478 3120
rect 180150 3108 180156 3120
rect 179472 3080 180156 3108
rect 179472 3068 179478 3080
rect 180150 3068 180156 3080
rect 180208 3068 180214 3120
rect 182542 3068 182548 3120
rect 182600 3108 182606 3120
rect 183462 3108 183468 3120
rect 182600 3080 183468 3108
rect 182600 3068 182606 3080
rect 183462 3068 183468 3080
rect 183520 3068 183526 3120
rect 187694 3068 187700 3120
rect 187752 3108 187758 3120
rect 188430 3108 188436 3120
rect 187752 3080 188436 3108
rect 187752 3068 187758 3080
rect 188430 3068 188436 3080
rect 188488 3068 188494 3120
rect 189626 3068 189632 3120
rect 189684 3108 189690 3120
rect 190362 3108 190368 3120
rect 189684 3080 190368 3108
rect 189684 3068 189690 3080
rect 190362 3068 190368 3080
rect 190420 3068 190426 3120
rect 192018 3068 192024 3120
rect 192076 3108 192082 3120
rect 193122 3108 193128 3120
rect 192076 3080 193128 3108
rect 192076 3068 192082 3080
rect 193122 3068 193128 3080
rect 193180 3068 193186 3120
rect 197998 3068 198004 3120
rect 198056 3108 198062 3120
rect 198642 3108 198648 3120
rect 198056 3080 198648 3108
rect 198056 3068 198062 3080
rect 198642 3068 198648 3080
rect 198700 3068 198706 3120
rect 199194 3068 199200 3120
rect 199252 3108 199258 3120
rect 199930 3108 199936 3120
rect 199252 3080 199936 3108
rect 199252 3068 199258 3080
rect 199930 3068 199936 3080
rect 199988 3068 199994 3120
rect 200390 3068 200396 3120
rect 200448 3108 200454 3120
rect 201402 3108 201408 3120
rect 200448 3080 201408 3108
rect 200448 3068 200454 3080
rect 201402 3068 201408 3080
rect 201460 3068 201466 3120
rect 201494 3068 201500 3120
rect 201552 3108 201558 3120
rect 202690 3108 202696 3120
rect 201552 3080 202696 3108
rect 201552 3068 201558 3080
rect 202690 3068 202696 3080
rect 202748 3068 202754 3120
rect 209501 3111 209559 3117
rect 209501 3077 209513 3111
rect 209547 3108 209559 3111
rect 219529 3111 219587 3117
rect 219529 3108 219541 3111
rect 209547 3080 219541 3108
rect 209547 3077 209559 3080
rect 209501 3071 209559 3077
rect 219529 3077 219541 3080
rect 219575 3077 219587 3111
rect 219529 3071 219587 3077
rect 219912 3080 231992 3108
rect 211065 3043 211123 3049
rect 211065 3009 211077 3043
rect 211111 3040 211123 3043
rect 219912 3040 219940 3080
rect 211111 3012 219940 3040
rect 220817 3043 220875 3049
rect 211111 3009 211123 3012
rect 211065 3003 211123 3009
rect 220817 3009 220829 3043
rect 220863 3040 220875 3043
rect 229097 3043 229155 3049
rect 229097 3040 229109 3043
rect 220863 3012 229109 3040
rect 220863 3009 220875 3012
rect 220817 3003 220875 3009
rect 229097 3009 229109 3012
rect 229143 3009 229155 3043
rect 231964 3040 231992 3080
rect 232498 3068 232504 3120
rect 232556 3108 232562 3120
rect 233142 3108 233148 3120
rect 232556 3080 233148 3108
rect 232556 3068 232562 3080
rect 233142 3068 233148 3080
rect 233200 3068 233206 3120
rect 235994 3068 236000 3120
rect 236052 3108 236058 3120
rect 237190 3108 237196 3120
rect 236052 3080 237196 3108
rect 236052 3068 236058 3080
rect 237190 3068 237196 3080
rect 237248 3068 237254 3120
rect 239582 3068 239588 3120
rect 239640 3108 239646 3120
rect 240042 3108 240048 3120
rect 239640 3080 240048 3108
rect 239640 3068 239646 3080
rect 240042 3068 240048 3080
rect 240100 3068 240106 3120
rect 240778 3068 240784 3120
rect 240836 3108 240842 3120
rect 241422 3108 241428 3120
rect 240836 3080 241428 3108
rect 240836 3068 240842 3080
rect 241422 3068 241428 3080
rect 241480 3068 241486 3120
rect 241974 3068 241980 3120
rect 242032 3108 242038 3120
rect 242802 3108 242808 3120
rect 242032 3080 242808 3108
rect 242032 3068 242038 3080
rect 242802 3068 242808 3080
rect 242860 3068 242866 3120
rect 234798 3040 234804 3052
rect 231964 3012 234804 3040
rect 229097 3003 229155 3009
rect 234798 3000 234804 3012
rect 234856 3000 234862 3052
rect 234893 3043 234951 3049
rect 234893 3009 234905 3043
rect 234939 3040 234951 3043
rect 246316 3040 246344 3148
rect 255038 3136 255044 3148
rect 255096 3136 255102 3188
rect 234939 3012 246344 3040
rect 248969 3043 249027 3049
rect 234939 3009 234951 3012
rect 234893 3003 234951 3009
rect 248969 3009 248981 3043
rect 249015 3040 249027 3043
rect 266372 3040 266400 3216
rect 269224 3176 269252 3216
rect 274082 3204 274088 3256
rect 274140 3244 274146 3256
rect 274542 3244 274548 3256
rect 274140 3216 274548 3244
rect 274140 3204 274146 3216
rect 274542 3204 274548 3216
rect 274600 3204 274606 3256
rect 277670 3204 277676 3256
rect 277728 3244 277734 3256
rect 278682 3244 278688 3256
rect 277728 3216 278688 3244
rect 277728 3204 277734 3216
rect 278682 3204 278688 3216
rect 278740 3204 278746 3256
rect 287146 3204 287152 3256
rect 287204 3244 287210 3256
rect 479518 3244 479524 3256
rect 287204 3216 479524 3244
rect 287204 3204 287210 3216
rect 479518 3204 479524 3216
rect 479576 3204 479582 3256
rect 483474 3204 483480 3256
rect 483532 3244 483538 3256
rect 484302 3244 484308 3256
rect 483532 3216 484308 3244
rect 483532 3204 483538 3216
rect 484302 3204 484308 3216
rect 484360 3204 484366 3256
rect 485774 3204 485780 3256
rect 485832 3244 485838 3256
rect 487062 3244 487068 3256
rect 485832 3216 487068 3244
rect 485832 3204 485838 3216
rect 487062 3204 487068 3216
rect 487120 3204 487126 3256
rect 490561 3247 490619 3253
rect 490561 3213 490573 3247
rect 490607 3244 490619 3247
rect 502981 3247 503039 3253
rect 502981 3244 502993 3247
rect 490607 3216 502993 3244
rect 490607 3213 490619 3216
rect 490561 3207 490619 3213
rect 502981 3213 502993 3216
rect 503027 3213 503039 3247
rect 502981 3207 503039 3213
rect 276474 3176 276480 3188
rect 269224 3148 276480 3176
rect 276474 3136 276480 3148
rect 276532 3136 276538 3188
rect 305086 3136 305092 3188
rect 305144 3176 305150 3188
rect 476758 3176 476764 3188
rect 305144 3148 476764 3176
rect 305144 3136 305150 3148
rect 476758 3136 476764 3148
rect 476816 3136 476822 3188
rect 477494 3136 477500 3188
rect 477552 3176 477558 3188
rect 498841 3179 498899 3185
rect 477552 3148 496860 3176
rect 477552 3136 477558 3148
rect 283561 3111 283619 3117
rect 283561 3077 283573 3111
rect 283607 3108 283619 3111
rect 297361 3111 297419 3117
rect 297361 3108 297373 3111
rect 283607 3080 297373 3108
rect 283607 3077 283619 3080
rect 283561 3071 283619 3077
rect 297361 3077 297373 3080
rect 297407 3077 297419 3111
rect 297361 3071 297419 3077
rect 356146 3068 356152 3120
rect 356204 3108 356210 3120
rect 387794 3108 387800 3120
rect 356204 3080 387800 3108
rect 356204 3068 356210 3080
rect 387794 3068 387800 3080
rect 387852 3068 387858 3120
rect 393961 3111 394019 3117
rect 393961 3077 393973 3111
rect 394007 3108 394019 3111
rect 402238 3108 402244 3120
rect 394007 3080 402244 3108
rect 394007 3077 394019 3080
rect 393961 3071 394019 3077
rect 402238 3068 402244 3080
rect 402296 3068 402302 3120
rect 411162 3068 411168 3120
rect 411220 3108 411226 3120
rect 415581 3111 415639 3117
rect 415581 3108 415593 3111
rect 411220 3080 415593 3108
rect 411220 3068 411226 3080
rect 415581 3077 415593 3080
rect 415627 3077 415639 3111
rect 415581 3071 415639 3077
rect 421558 3068 421564 3120
rect 421616 3108 421622 3120
rect 422202 3108 422208 3120
rect 421616 3080 422208 3108
rect 421616 3068 421622 3080
rect 422202 3068 422208 3080
rect 422260 3068 422266 3120
rect 430117 3111 430175 3117
rect 430117 3077 430129 3111
rect 430163 3108 430175 3111
rect 440602 3108 440608 3120
rect 430163 3080 440608 3108
rect 430163 3077 430175 3080
rect 430117 3071 430175 3077
rect 440602 3068 440608 3080
rect 440660 3068 440666 3120
rect 447778 3068 447784 3120
rect 447836 3108 447842 3120
rect 496725 3111 496783 3117
rect 496725 3108 496737 3111
rect 447836 3080 496737 3108
rect 447836 3068 447842 3080
rect 496725 3077 496737 3080
rect 496771 3077 496783 3111
rect 496832 3108 496860 3148
rect 498841 3145 498853 3179
rect 498887 3176 498899 3179
rect 503070 3176 503076 3188
rect 498887 3148 503076 3176
rect 498887 3145 498899 3148
rect 498841 3139 498899 3145
rect 503070 3136 503076 3148
rect 503128 3136 503134 3188
rect 503180 3176 503208 3284
rect 503257 3247 503315 3253
rect 503257 3213 503269 3247
rect 503303 3244 503315 3247
rect 510706 3244 510712 3256
rect 503303 3216 510712 3244
rect 503303 3213 503315 3216
rect 503257 3207 503315 3213
rect 510706 3204 510712 3216
rect 510764 3204 510770 3256
rect 507946 3176 507952 3188
rect 503180 3148 507952 3176
rect 507946 3136 507952 3148
rect 508004 3136 508010 3188
rect 508038 3108 508044 3120
rect 496832 3080 508044 3108
rect 496725 3071 496783 3077
rect 508038 3068 508044 3080
rect 508096 3068 508102 3120
rect 249015 3012 266400 3040
rect 249015 3009 249027 3012
rect 248969 3003 249027 3009
rect 296714 3000 296720 3052
rect 296772 3040 296778 3052
rect 297910 3040 297916 3052
rect 296772 3012 297916 3040
rect 296772 3000 296778 3012
rect 297910 3000 297916 3012
rect 297968 3000 297974 3052
rect 450170 3000 450176 3052
rect 450228 3040 450234 3052
rect 509234 3040 509240 3052
rect 450228 3012 509240 3040
rect 450228 3000 450234 3012
rect 509234 3000 509240 3012
rect 509292 3000 509298 3052
rect 201497 2975 201555 2981
rect 201497 2972 201509 2975
rect 179248 2944 180564 2972
rect 158714 2904 158720 2916
rect 85172 2876 136864 2904
rect 139412 2876 158720 2904
rect 85172 2864 85178 2876
rect 76926 2796 76932 2848
rect 76984 2836 76990 2848
rect 133782 2836 133788 2848
rect 76984 2808 133788 2836
rect 76984 2796 76990 2808
rect 133782 2796 133788 2808
rect 133840 2796 133846 2848
rect 133877 2839 133935 2845
rect 133877 2805 133889 2839
rect 133923 2836 133935 2839
rect 136729 2839 136787 2845
rect 136729 2836 136741 2839
rect 133923 2808 136741 2836
rect 133923 2805 133935 2808
rect 133877 2799 133935 2805
rect 136729 2805 136741 2808
rect 136775 2805 136787 2839
rect 136836 2836 136864 2876
rect 158714 2864 158720 2876
rect 158772 2864 158778 2916
rect 180536 2904 180564 2944
rect 193232 2944 201509 2972
rect 193232 2904 193260 2944
rect 201497 2941 201509 2944
rect 201543 2941 201555 2975
rect 201497 2935 201555 2941
rect 249061 2975 249119 2981
rect 249061 2941 249073 2975
rect 249107 2972 249119 2975
rect 258721 2975 258779 2981
rect 258721 2972 258733 2975
rect 249107 2944 258733 2972
rect 249107 2941 249119 2944
rect 249061 2935 249119 2941
rect 258721 2941 258733 2944
rect 258767 2941 258779 2975
rect 258721 2935 258779 2941
rect 451274 2932 451280 2984
rect 451332 2972 451338 2984
rect 452470 2972 452476 2984
rect 451332 2944 452476 2972
rect 451332 2932 451338 2944
rect 452470 2932 452476 2944
rect 452528 2932 452534 2984
rect 456058 2932 456064 2984
rect 456116 2972 456122 2984
rect 456702 2972 456708 2984
rect 456116 2944 456708 2972
rect 456116 2932 456122 2944
rect 456702 2932 456708 2944
rect 456760 2932 456766 2984
rect 466822 2932 466828 2984
rect 466880 2972 466886 2984
rect 467742 2972 467748 2984
rect 466880 2944 467748 2972
rect 466880 2932 466886 2944
rect 467742 2932 467748 2944
rect 467800 2932 467806 2984
rect 471514 2932 471520 2984
rect 471572 2972 471578 2984
rect 506382 2972 506388 2984
rect 471572 2944 506388 2972
rect 471572 2932 471578 2944
rect 506382 2932 506388 2944
rect 506440 2932 506446 2984
rect 180536 2876 193260 2904
rect 208489 2907 208547 2913
rect 208489 2873 208501 2907
rect 208535 2904 208547 2907
rect 220081 2907 220139 2913
rect 220081 2904 220093 2907
rect 208535 2876 220093 2904
rect 208535 2873 208547 2876
rect 208489 2867 208547 2873
rect 220081 2873 220093 2876
rect 220127 2873 220139 2907
rect 220081 2867 220139 2873
rect 229097 2907 229155 2913
rect 229097 2873 229109 2907
rect 229143 2904 229155 2907
rect 234893 2907 234951 2913
rect 234893 2904 234905 2907
rect 229143 2876 234905 2904
rect 229143 2873 229155 2876
rect 229097 2867 229155 2873
rect 234893 2873 234905 2876
rect 234939 2873 234951 2907
rect 234893 2867 234951 2873
rect 471146 2864 471152 2916
rect 471204 2904 471210 2916
rect 484578 2904 484584 2916
rect 471204 2876 484584 2904
rect 471204 2864 471210 2876
rect 484578 2864 484584 2876
rect 484636 2864 484642 2916
rect 489362 2864 489368 2916
rect 489420 2904 489426 2916
rect 510614 2904 510620 2916
rect 489420 2876 510620 2904
rect 489420 2864 489426 2876
rect 510614 2864 510620 2876
rect 510672 2864 510678 2916
rect 571978 2864 571984 2916
rect 572036 2904 572042 2916
rect 578602 2904 578608 2916
rect 572036 2876 578608 2904
rect 572036 2864 572042 2876
rect 578602 2864 578608 2876
rect 578660 2864 578666 2916
rect 142062 2836 142068 2848
rect 136836 2808 142068 2836
rect 136729 2799 136787 2805
rect 142062 2796 142068 2808
rect 142120 2796 142126 2848
rect 142801 2839 142859 2845
rect 142801 2805 142813 2839
rect 142847 2836 142859 2839
rect 154117 2839 154175 2845
rect 154117 2836 154129 2839
rect 142847 2808 154129 2836
rect 142847 2805 142859 2808
rect 142801 2799 142859 2805
rect 154117 2805 154129 2808
rect 154163 2805 154175 2839
rect 154117 2799 154175 2805
rect 154209 2839 154267 2845
rect 154209 2805 154221 2839
rect 154255 2836 154267 2839
rect 157245 2839 157303 2845
rect 157245 2836 157257 2839
rect 154255 2808 157257 2836
rect 154255 2805 154267 2808
rect 154209 2799 154267 2805
rect 157245 2805 157257 2808
rect 157291 2805 157303 2839
rect 157245 2799 157303 2805
rect 157337 2839 157395 2845
rect 157337 2805 157349 2839
rect 157383 2836 157395 2839
rect 166905 2839 166963 2845
rect 166905 2836 166917 2839
rect 157383 2808 166917 2836
rect 157383 2805 157395 2808
rect 157337 2799 157395 2805
rect 166905 2805 166917 2808
rect 166951 2805 166963 2839
rect 166905 2799 166963 2805
rect 201497 2839 201555 2845
rect 201497 2805 201509 2839
rect 201543 2836 201555 2839
rect 211065 2839 211123 2845
rect 211065 2836 211077 2839
rect 201543 2808 211077 2836
rect 201543 2805 201555 2808
rect 201497 2799 201555 2805
rect 211065 2805 211077 2808
rect 211111 2805 211123 2839
rect 211065 2799 211123 2805
rect 358814 2796 358820 2848
rect 358872 2836 358878 2848
rect 358872 2808 359780 2836
rect 358872 2796 358878 2808
rect 359752 2780 359780 2808
rect 384666 2796 384672 2848
rect 384724 2836 384730 2848
rect 384942 2836 384948 2848
rect 384724 2808 384948 2836
rect 384724 2796 384730 2808
rect 384942 2796 384948 2808
rect 385000 2796 385006 2848
rect 481082 2796 481088 2848
rect 481140 2836 481146 2848
rect 490561 2839 490619 2845
rect 490561 2836 490573 2839
rect 481140 2808 490573 2836
rect 481140 2796 481146 2808
rect 490561 2805 490573 2808
rect 490607 2805 490619 2839
rect 490561 2799 490619 2805
rect 490653 2839 490711 2845
rect 490653 2805 490665 2839
rect 490699 2836 490711 2839
rect 494977 2839 495035 2845
rect 494977 2836 494989 2839
rect 490699 2808 494989 2836
rect 490699 2805 490711 2808
rect 490653 2799 490711 2805
rect 494977 2805 494989 2808
rect 495023 2805 495035 2839
rect 494977 2799 495035 2805
rect 496725 2839 496783 2845
rect 496725 2805 496737 2839
rect 496771 2836 496783 2839
rect 499485 2839 499543 2845
rect 499485 2836 499497 2839
rect 496771 2808 499497 2836
rect 496771 2805 496783 2808
rect 496725 2799 496783 2805
rect 499485 2805 499497 2808
rect 499531 2805 499543 2839
rect 508222 2836 508228 2848
rect 499485 2799 499543 2805
rect 500328 2808 508228 2836
rect 85574 2728 85580 2780
rect 85632 2768 85638 2780
rect 95142 2768 95148 2780
rect 85632 2740 95148 2768
rect 85632 2728 85638 2740
rect 95142 2728 95148 2740
rect 95200 2728 95206 2780
rect 96890 2728 96896 2780
rect 96948 2768 96954 2780
rect 109037 2771 109095 2777
rect 109037 2768 109049 2771
rect 96948 2740 109049 2768
rect 96948 2728 96954 2740
rect 109037 2737 109049 2740
rect 109083 2737 109095 2771
rect 109037 2731 109095 2737
rect 122837 2771 122895 2777
rect 122837 2737 122849 2771
rect 122883 2768 122895 2771
rect 132405 2771 132463 2777
rect 132405 2768 132417 2771
rect 122883 2740 132417 2768
rect 122883 2737 122895 2740
rect 122837 2731 122895 2737
rect 132405 2737 132417 2740
rect 132451 2737 132463 2771
rect 132405 2731 132463 2737
rect 161382 2728 161388 2780
rect 161440 2768 161446 2780
rect 162302 2768 162308 2780
rect 161440 2740 162308 2768
rect 161440 2728 161446 2740
rect 162302 2728 162308 2740
rect 162360 2728 162366 2780
rect 359734 2728 359740 2780
rect 359792 2728 359798 2780
rect 499577 2771 499635 2777
rect 499577 2737 499589 2771
rect 499623 2768 499635 2771
rect 500328 2768 500356 2808
rect 508222 2796 508228 2808
rect 508280 2796 508286 2848
rect 499623 2740 500356 2768
rect 499623 2737 499635 2740
rect 499577 2731 499635 2737
rect 563054 2728 563060 2780
rect 563112 2768 563118 2780
rect 564342 2768 564348 2780
rect 563112 2740 564348 2768
rect 563112 2728 563118 2740
rect 564342 2728 564348 2740
rect 564400 2728 564406 2780
rect 304994 1232 305000 1284
rect 305052 1272 305058 1284
rect 306190 1272 306196 1284
rect 305052 1244 306196 1272
rect 305052 1232 305058 1244
rect 306190 1232 306196 1244
rect 306248 1232 306254 1284
rect 80238 552 80244 604
rect 80296 592 80302 604
rect 80330 592 80336 604
rect 80296 564 80336 592
rect 80296 552 80302 564
rect 80330 552 80336 564
rect 80388 552 80394 604
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92382 592 92388 604
rect 92164 564 92388 592
rect 92164 552 92170 564
rect 92382 552 92388 564
rect 92440 552 92446 604
rect 100478 592 100484 604
rect 100439 564 100484 592
rect 100478 552 100484 564
rect 100536 552 100542 604
rect 111150 592 111156 604
rect 111111 564 111156 592
rect 111150 552 111156 564
rect 111208 552 111214 604
rect 134886 592 134892 604
rect 134847 564 134892 592
rect 134886 552 134892 564
rect 134944 552 134950 604
rect 186038 592 186044 604
rect 185999 564 186044 592
rect 186038 552 186044 564
rect 186096 552 186102 604
rect 190362 552 190368 604
rect 190420 592 190426 604
rect 190822 592 190828 604
rect 190420 564 190828 592
rect 190420 552 190426 564
rect 190822 552 190828 564
rect 190880 552 190886 604
rect 205634 552 205640 604
rect 205692 592 205698 604
rect 206278 592 206284 604
rect 205692 564 206284 592
rect 205692 552 205698 564
rect 206278 552 206284 564
rect 206336 552 206342 604
rect 212534 552 212540 604
rect 212592 592 212598 604
rect 213454 592 213460 604
rect 212592 564 213460 592
rect 212592 552 212598 564
rect 213454 552 213460 564
rect 213512 552 213518 604
rect 247954 552 247960 604
rect 248012 592 248018 604
rect 248322 592 248328 604
rect 248012 564 248328 592
rect 248012 552 248018 564
rect 248322 552 248328 564
rect 248380 552 248386 604
rect 258626 592 258632 604
rect 258587 564 258632 592
rect 258626 552 258632 564
rect 258684 552 258690 604
rect 289538 552 289544 604
rect 289596 592 289602 604
rect 289906 592 289912 604
rect 289596 564 289912 592
rect 289596 552 289602 564
rect 289906 552 289912 564
rect 289964 552 289970 604
rect 370406 592 370412 604
rect 370367 564 370412 592
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 371602 592 371608 604
rect 371563 564 371608 592
rect 371602 552 371608 564
rect 371660 552 371666 604
rect 372798 592 372804 604
rect 372759 564 372804 592
rect 372798 552 372804 564
rect 372856 552 372862 604
rect 377582 592 377588 604
rect 377543 564 377588 592
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 378778 592 378784 604
rect 378739 564 378784 592
rect 378778 552 378784 564
rect 378836 552 378842 604
rect 396074 552 396080 604
rect 396132 592 396138 604
rect 396626 592 396632 604
rect 396132 564 396632 592
rect 396132 552 396138 564
rect 396626 552 396632 564
rect 396684 552 396690 604
rect 412634 552 412640 604
rect 412692 592 412698 604
rect 413278 592 413284 604
rect 412692 564 413284 592
rect 412692 552 412698 564
rect 413278 552 413284 564
rect 413336 552 413342 604
rect 428734 592 428740 604
rect 428695 564 428740 592
rect 428734 552 428740 564
rect 428792 552 428798 604
rect 437014 592 437020 604
rect 436975 564 437020 592
rect 437014 552 437020 564
rect 437072 552 437078 604
rect 437474 552 437480 604
rect 437532 592 437538 604
rect 438210 592 438216 604
rect 437532 564 438216 592
rect 437532 552 437538 564
rect 438210 552 438216 564
rect 438268 552 438274 604
rect 444466 552 444472 604
rect 444524 592 444530 604
rect 445386 592 445392 604
rect 444524 564 445392 592
rect 444524 552 444530 564
rect 445386 552 445392 564
rect 445444 552 445450 604
rect 445754 552 445760 604
rect 445812 592 445818 604
rect 446582 592 446588 604
rect 445812 564 446588 592
rect 445812 552 445818 564
rect 446582 552 446588 564
rect 446640 552 446646 604
rect 448514 552 448520 604
rect 448572 592 448578 604
rect 448974 592 448980 604
rect 448572 564 448980 592
rect 448572 552 448578 564
rect 448974 552 448980 564
rect 449032 552 449038 604
rect 453666 552 453672 604
rect 453724 592 453730 604
rect 453942 592 453948 604
rect 453724 564 453948 592
rect 453724 552 453730 564
rect 453942 552 453948 564
rect 454000 552 454006 604
rect 454034 552 454040 604
rect 454092 592 454098 604
rect 454862 592 454868 604
rect 454092 564 454868 592
rect 454092 552 454098 564
rect 454862 552 454868 564
rect 454920 552 454926 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
rect 492674 552 492680 604
rect 492732 592 492738 604
rect 492950 592 492956 604
rect 492732 564 492956 592
rect 492732 552 492738 564
rect 492950 552 492956 564
rect 493008 552 493014 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 506658 552 506664 604
rect 506716 592 506722 604
rect 507210 592 507216 604
rect 506716 564 507216 592
rect 506716 552 506722 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 512086 552 512092 604
rect 512144 592 512150 604
rect 513190 592 513196 604
rect 512144 564 513196 592
rect 512144 552 512150 564
rect 513190 552 513196 564
rect 513248 552 513254 604
rect 513374 552 513380 604
rect 513432 592 513438 604
rect 514386 592 514392 604
rect 513432 564 514392 592
rect 513432 552 513438 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 514754 552 514760 604
rect 514812 592 514818 604
rect 515582 592 515588 604
rect 514812 564 515588 592
rect 514812 552 514818 564
rect 515582 552 515588 564
rect 515640 552 515646 604
rect 576854 552 576860 604
rect 576912 592 576918 604
rect 577406 592 577412 604
rect 576912 564 577412 592
rect 576912 552 576918 564
rect 577406 552 577412 564
rect 577464 552 577470 604
rect 579614 552 579620 604
rect 579672 592 579678 604
rect 579798 592 579804 604
rect 579672 564 579804 592
rect 579672 552 579678 564
rect 579798 552 579804 564
rect 579856 552 579862 604
<< via1 >>
rect 335268 700816 335320 700868
rect 429844 700816 429896 700868
rect 283840 700748 283892 700800
rect 343640 700748 343692 700800
rect 364984 700748 365036 700800
rect 508136 700748 508188 700800
rect 78220 700680 78272 700732
rect 235172 700680 235224 700732
rect 269028 700680 269080 700732
rect 300124 700680 300176 700732
rect 332508 700680 332560 700732
rect 501604 700680 501656 700732
rect 137836 700612 137888 700664
rect 386420 700612 386472 700664
rect 397460 700612 397512 700664
rect 502524 700612 502576 700664
rect 81900 700544 81952 700596
rect 170312 700544 170364 700596
rect 202788 700544 202840 700596
rect 501788 700544 501840 700596
rect 40500 700476 40552 700528
rect 402980 700476 403032 700528
rect 81440 700408 81492 700460
rect 462320 700408 462372 700460
rect 494796 700408 494848 700460
rect 508412 700408 508464 700460
rect 79968 700340 80020 700392
rect 478512 700340 478564 700392
rect 504456 700340 504508 700392
rect 543464 700340 543516 700392
rect 8116 700272 8168 700324
rect 19984 700272 20036 700324
rect 72976 700272 73028 700324
rect 77944 700272 77996 700324
rect 78588 700272 78640 700324
rect 105452 700272 105504 700324
rect 142068 700272 142120 700324
rect 559656 700272 559708 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 412824 692724 412876 692776
rect 508780 685856 508832 685908
rect 580172 685856 580224 685908
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 412640 683068 412692 683120
rect 3516 681708 3568 681760
rect 9312 681708 9364 681760
rect 81532 673480 81584 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 502616 667904 502668 667956
rect 413100 666544 413152 666596
rect 3056 652740 3108 652792
rect 15936 652740 15988 652792
rect 190368 650020 190420 650072
rect 580172 650020 580224 650072
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 507124 638936 507176 638988
rect 580172 638936 580224 638988
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 82084 626560 82136 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 14464 623772 14516 623824
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 3424 609968 3476 610020
rect 8852 609968 8904 610020
rect 412824 608583 412876 608592
rect 412824 608549 412833 608583
rect 412833 608549 412867 608583
rect 412867 608549 412876 608583
rect 412824 608540 412876 608549
rect 83556 603100 83608 603152
rect 580172 603100 580224 603152
rect 413008 601672 413060 601724
rect 413008 598884 413060 598936
rect 3240 594804 3292 594856
rect 31116 594804 31168 594856
rect 89352 593308 89404 593360
rect 89444 593308 89496 593360
rect 507216 592016 507268 592068
rect 580172 592016 580224 592068
rect 83556 590724 83608 590776
rect 83740 590724 83792 590776
rect 412916 589339 412968 589348
rect 412916 589305 412925 589339
rect 412925 589305 412959 589339
rect 412959 589305 412968 589339
rect 412916 589296 412968 589305
rect 78496 586508 78548 586560
rect 236920 586508 236972 586560
rect 83556 586440 83608 586492
rect 83648 586372 83700 586424
rect 46204 585080 46256 585132
rect 163136 585080 163188 585132
rect 189264 585080 189316 585132
rect 190368 585080 190420 585132
rect 197084 585080 197136 585132
rect 477592 585080 477644 585132
rect 487160 585080 487212 585132
rect 509884 585080 509936 585132
rect 90916 585012 90968 585064
rect 432328 585012 432380 585064
rect 439504 585012 439556 585064
rect 511356 585012 511408 585064
rect 71044 584944 71096 584996
rect 468024 584944 468076 584996
rect 475200 584944 475252 584996
rect 508044 584944 508096 584996
rect 57244 584876 57296 584928
rect 470416 584876 470468 584928
rect 479984 584876 480036 584928
rect 511264 584876 511316 584928
rect 92112 584808 92164 584860
rect 167920 584808 167972 584860
rect 182272 584808 182324 584860
rect 191748 584808 191800 584860
rect 446680 584808 446732 584860
rect 506480 584808 506532 584860
rect 105360 584740 105412 584792
rect 215576 584740 215628 584792
rect 226340 584740 226392 584792
rect 294144 584740 294196 584792
rect 437112 584740 437164 584792
rect 506572 584740 506624 584792
rect 77024 584672 77076 584724
rect 103520 584672 103572 584724
rect 117872 584672 117924 584724
rect 233240 584672 233292 584724
rect 238760 584672 238812 584724
rect 244096 584672 244148 584724
rect 456064 584672 456116 584724
rect 507952 584672 508004 584724
rect 61384 584604 61436 584656
rect 217968 584604 218020 584656
rect 227812 584604 227864 584656
rect 234528 584604 234580 584656
rect 249708 584604 249760 584656
rect 372712 584604 372764 584656
rect 377496 584604 377548 584656
rect 494704 584604 494756 584656
rect 508320 584604 508372 584656
rect 60004 584536 60056 584588
rect 248880 584536 248932 584588
rect 348976 584536 349028 584588
rect 485780 584536 485832 584588
rect 491944 584536 491996 584588
rect 511172 584536 511224 584588
rect 64144 584468 64196 584520
rect 270408 584468 270460 584520
rect 382280 584468 382332 584520
rect 524420 584468 524472 584520
rect 50344 584400 50396 584452
rect 272800 584400 272852 584452
rect 444288 584400 444340 584452
rect 505284 584400 505336 584452
rect 53104 584332 53156 584384
rect 322664 584332 322716 584384
rect 367928 584332 367980 584384
rect 510804 584332 510856 584384
rect 31024 584264 31076 584316
rect 310888 584264 310940 584316
rect 341800 584264 341852 584316
rect 501512 584264 501564 584316
rect 76932 584196 76984 584248
rect 210792 584196 210844 584248
rect 339408 584196 339460 584248
rect 456800 584196 456852 584248
rect 458456 584196 458508 584248
rect 505376 584196 505428 584248
rect 51724 584128 51776 584180
rect 356152 584128 356204 584180
rect 370320 584128 370372 584180
rect 556160 584128 556212 584180
rect 75184 584060 75236 584112
rect 77208 583992 77260 584044
rect 96344 583992 96396 584044
rect 131948 584060 132000 584112
rect 449072 584060 449124 584112
rect 453856 584060 453908 584112
rect 534080 584060 534132 584112
rect 136824 583992 136876 584044
rect 141608 583992 141660 584044
rect 142068 583992 142120 584044
rect 170312 583992 170364 584044
rect 490380 583992 490432 584044
rect 494336 583992 494388 584044
rect 511540 583992 511592 584044
rect 73804 583924 73856 583976
rect 127440 583924 127492 583976
rect 268016 583924 268068 583976
rect 269028 583924 269080 583976
rect 289360 583924 289412 583976
rect 455328 583924 455380 583976
rect 484768 583924 484820 583976
rect 509792 583924 509844 583976
rect 42064 583856 42116 583908
rect 413192 583856 413244 583908
rect 422760 583856 422812 583908
rect 509424 583856 509476 583908
rect 78312 583788 78364 583840
rect 105912 583788 105964 583840
rect 107660 583788 107712 583840
rect 125048 583788 125100 583840
rect 415584 583788 415636 583840
rect 502340 583788 502392 583840
rect 78404 583720 78456 583772
rect 113088 583720 113140 583772
rect 308496 583720 308548 583772
rect 314660 583720 314712 583772
rect 408592 583720 408644 583772
rect 424968 583720 425020 583772
rect 429936 583720 429988 583772
rect 501328 583720 501380 583772
rect 505836 583720 505888 583772
rect 35808 583448 35860 583500
rect 441896 583448 441948 583500
rect 485780 583448 485832 583500
rect 502984 583448 503036 583500
rect 75828 583380 75880 583432
rect 131948 583380 132000 583432
rect 456800 583380 456852 583432
rect 509516 583380 509568 583432
rect 77116 583312 77168 583364
rect 197084 583312 197136 583364
rect 455328 583312 455380 583364
rect 510988 583312 511040 583364
rect 75276 583244 75328 583296
rect 279792 583244 279844 583296
rect 410800 583244 410852 583296
rect 503352 583244 503404 583296
rect 10416 583176 10468 583228
rect 256056 583176 256108 583228
rect 379888 583176 379940 583228
rect 503076 583176 503128 583228
rect 9496 583108 9548 583160
rect 265624 583108 265676 583160
rect 337016 583108 337068 583160
rect 509700 583108 509752 583160
rect 10600 583040 10652 583092
rect 284576 583040 284628 583092
rect 327448 583040 327500 583092
rect 507676 583040 507728 583092
rect 77760 582972 77812 583024
rect 353760 582972 353812 583024
rect 360936 582972 360988 583024
rect 510068 582972 510120 583024
rect 80704 582904 80756 582956
rect 198832 582904 198884 582956
rect 229744 582904 229796 582956
rect 510896 582904 510948 582956
rect 184480 582836 184532 582888
rect 503260 582836 503312 582888
rect 15844 582768 15896 582820
rect 110696 582768 110748 582820
rect 177488 582768 177540 582820
rect 501972 582768 502024 582820
rect 8944 582700 8996 582752
rect 146392 582700 146444 582752
rect 220360 582700 220412 582752
rect 560944 582700 560996 582752
rect 10692 582632 10744 582684
rect 129832 582632 129884 582684
rect 132224 582632 132276 582684
rect 503168 582632 503220 582684
rect 86316 582564 86368 582616
rect 96528 582564 96580 582616
rect 96620 582564 96672 582616
rect 101312 582564 101364 582616
rect 115848 582564 115900 582616
rect 425152 582564 425204 582616
rect 514024 582564 514076 582616
rect 64788 582496 64840 582548
rect 499120 582496 499172 582548
rect 9588 582428 9640 582480
rect 463240 582428 463292 582480
rect 482376 582428 482428 582480
rect 507492 582428 507544 582480
rect 6184 582360 6236 582412
rect 489552 582360 489604 582412
rect 490196 582360 490248 582412
rect 497556 582360 497608 582412
rect 90456 582292 90508 582344
rect 99840 582292 99892 582344
rect 111064 582292 111116 582344
rect 460848 582292 460900 582344
rect 510712 582292 510764 582344
rect 10508 582224 10560 582276
rect 93952 582224 94004 582276
rect 100024 582224 100076 582276
rect 105360 582224 105412 582276
rect 118700 582224 118752 582276
rect 123760 582224 123812 582276
rect 150992 582224 151044 582276
rect 157156 582224 157208 582276
rect 157248 582224 157300 582276
rect 162492 582224 162544 582276
rect 494704 582224 494756 582276
rect 511080 582224 511132 582276
rect 93216 582156 93268 582208
rect 122656 582156 122708 582208
rect 128360 582156 128412 582208
rect 137928 582156 137980 582208
rect 146944 582156 146996 582208
rect 160468 582156 160520 582208
rect 167092 582156 167144 582208
rect 176568 582156 176620 582208
rect 401416 582156 401468 582208
rect 502064 582156 502116 582208
rect 73068 582088 73120 582140
rect 226340 582088 226392 582140
rect 406200 582088 406252 582140
rect 509332 582088 509384 582140
rect 89720 582020 89772 582072
rect 91928 582020 91980 582072
rect 92664 582020 92716 582072
rect 286692 582020 286744 582072
rect 394608 582020 394660 582072
rect 509608 582020 509660 582072
rect 85212 581952 85264 582004
rect 320180 581952 320232 582004
rect 321560 581952 321612 582004
rect 326436 581952 326488 582004
rect 363696 581952 363748 582004
rect 501880 581952 501932 582004
rect 48228 581884 48280 581936
rect 372620 581884 372672 581936
rect 399392 581884 399444 581936
rect 543740 581884 543792 581936
rect 3424 581816 3476 581868
rect 262956 581816 263008 581868
rect 296720 581816 296772 581868
rect 510620 581816 510672 581868
rect 85488 581748 85540 581800
rect 172520 581748 172572 581800
rect 186320 581748 186372 581800
rect 192208 581748 192260 581800
rect 246856 581748 246908 581800
rect 508228 581748 508280 581800
rect 52368 581680 52420 581732
rect 249708 581680 249760 581732
rect 251640 581680 251692 581732
rect 554872 581680 554924 581732
rect 9128 581612 9180 581664
rect 120080 581612 120132 581664
rect 134340 581655 134392 581664
rect 134340 581621 134349 581655
rect 134349 581621 134383 581655
rect 134383 581621 134392 581655
rect 134340 581612 134392 581621
rect 144368 581655 144420 581664
rect 144368 581621 144377 581655
rect 144377 581621 144411 581655
rect 144411 581621 144420 581655
rect 144368 581612 144420 581621
rect 157064 581612 157116 581664
rect 157524 581612 157576 581664
rect 198004 581612 198056 581664
rect 200856 581612 200908 581664
rect 227720 581612 227772 581664
rect 532700 581612 532752 581664
rect 4804 581544 4856 581596
rect 313188 581544 313240 581596
rect 375288 581544 375340 581596
rect 569960 581544 570012 581596
rect 10324 581476 10376 581528
rect 165252 581476 165304 581528
rect 176568 581476 176620 581528
rect 176752 581476 176804 581528
rect 194416 581476 194468 581528
rect 505100 581476 505152 581528
rect 67548 581408 67600 581460
rect 420092 581408 420144 581460
rect 435088 581408 435140 581460
rect 580540 581408 580592 581460
rect 9220 581340 9272 581392
rect 98460 581340 98512 581392
rect 99472 581340 99524 581392
rect 103428 581340 103480 581392
rect 108672 581340 108724 581392
rect 491852 581340 491904 581392
rect 494612 581340 494664 581392
rect 504364 581340 504416 581392
rect 82636 581272 82688 581324
rect 580356 581272 580408 581324
rect 9036 581204 9088 581256
rect 580448 581204 580500 581256
rect 501696 581068 501748 581120
rect 501880 581068 501932 581120
rect 502064 581000 502116 581052
rect 501880 580932 501932 580984
rect 507308 579640 507360 579692
rect 580172 579640 580224 579692
rect 48964 572704 49016 572756
rect 78680 572704 78732 572756
rect 532700 568556 532752 568608
rect 532884 568556 532936 568608
rect 524420 568531 524472 568540
rect 524420 568497 524429 568531
rect 524429 568497 524463 568531
rect 524463 568497 524472 568531
rect 524420 568488 524472 568497
rect 3516 567196 3568 567248
rect 33784 567196 33836 567248
rect 503812 565836 503864 565888
rect 511724 565836 511776 565888
rect 503812 563048 503864 563100
rect 574100 563048 574152 563100
rect 70308 558900 70360 558952
rect 78680 558900 78732 558952
rect 532424 558900 532476 558952
rect 532516 558900 532568 558952
rect 504916 556248 504968 556300
rect 536840 556248 536892 556300
rect 529204 556180 529256 556232
rect 580172 556180 580224 556232
rect 532516 553256 532568 553308
rect 532884 553256 532936 553308
rect 3148 552032 3200 552084
rect 42156 552032 42208 552084
rect 504824 552032 504876 552084
rect 507400 552032 507452 552084
rect 524604 550604 524656 550656
rect 505008 549312 505060 549364
rect 508596 549312 508648 549364
rect 529940 545164 529992 545216
rect 531964 545164 532016 545216
rect 524420 543736 524472 543788
rect 524604 543736 524656 543788
rect 532700 540948 532752 541000
rect 532976 540948 533028 541000
rect 3516 538228 3568 538280
rect 9404 538228 9456 538280
rect 503352 534012 503404 534064
rect 580172 534012 580224 534064
rect 82820 529907 82872 529916
rect 82820 529873 82829 529907
rect 82829 529873 82863 529907
rect 82863 529873 82872 529907
rect 82820 529864 82872 529873
rect 505008 527144 505060 527196
rect 510160 527144 510212 527196
rect 532700 521636 532752 521688
rect 532884 521636 532936 521688
rect 82912 520276 82964 520328
rect 503720 514700 503772 514752
rect 503904 514700 503956 514752
rect 504456 510552 504508 510604
rect 580172 510552 580224 510604
rect 2872 509260 2924 509312
rect 17224 509260 17276 509312
rect 503720 505112 503772 505164
rect 503904 505112 503956 505164
rect 532700 502324 532752 502376
rect 532884 502324 532936 502376
rect 82820 501032 82872 501084
rect 82912 500964 82964 501016
rect 82820 500939 82872 500948
rect 82820 500905 82829 500939
rect 82829 500905 82863 500939
rect 82863 500905 82872 500939
rect 82820 500896 82872 500905
rect 501972 499468 502024 499520
rect 579988 499468 580040 499520
rect 3516 496748 3568 496800
rect 80704 496748 80756 496800
rect 505008 492668 505060 492720
rect 510252 492668 510304 492720
rect 532700 492600 532752 492652
rect 532884 492600 532936 492652
rect 82820 491351 82872 491360
rect 82820 491317 82829 491351
rect 82829 491317 82863 491351
rect 82863 491317 82872 491351
rect 82820 491308 82872 491317
rect 504456 485800 504508 485852
rect 519544 485800 519596 485852
rect 580172 485800 580224 485852
rect 511632 485732 511684 485784
rect 3332 481516 3384 481568
rect 8760 481516 8812 481568
rect 505008 478864 505060 478916
rect 513380 478864 513432 478916
rect 8852 478796 8904 478848
rect 77576 478796 77628 478848
rect 503720 475736 503772 475788
rect 504088 475736 504140 475788
rect 82636 474036 82688 474088
rect 82912 474036 82964 474088
rect 524420 471971 524472 471980
rect 524420 471937 524429 471971
rect 524429 471937 524463 471971
rect 524463 471937 524472 471971
rect 524420 471928 524472 471937
rect 503536 470568 503588 470620
rect 531964 470568 532016 470620
rect 524420 462451 524472 462460
rect 524420 462417 524429 462451
rect 524429 462417 524463 462451
rect 524463 462417 524472 462451
rect 524420 462408 524472 462417
rect 505744 462340 505796 462392
rect 580172 462340 580224 462392
rect 503720 461388 503772 461440
rect 504088 461388 504140 461440
rect 503720 456424 503772 456476
rect 504088 456424 504140 456476
rect 504548 454044 504600 454096
rect 510344 454044 510396 454096
rect 524420 452591 524472 452600
rect 524420 452557 524429 452591
rect 524429 452557 524463 452591
rect 524463 452557 524472 452591
rect 524420 452548 524472 452557
rect 82636 450168 82688 450220
rect 82912 450168 82964 450220
rect 83004 447788 83056 447840
rect 503720 447108 503772 447160
rect 504088 447108 504140 447160
rect 524420 443003 524472 443012
rect 524420 442969 524429 443003
rect 524429 442969 524463 443003
rect 524463 442969 524472 443003
rect 524420 442960 524472 442969
rect 82820 442892 82872 442944
rect 82820 442144 82872 442196
rect 83004 442144 83056 442196
rect 503260 440172 503312 440224
rect 579988 440172 580040 440224
rect 82912 439492 82964 439544
rect 82820 438132 82872 438184
rect 503720 437384 503772 437436
rect 504272 437384 504324 437436
rect 12348 436092 12400 436144
rect 75092 436092 75144 436144
rect 524420 433279 524472 433288
rect 524420 433245 524429 433279
rect 524429 433245 524463 433279
rect 524463 433245 524472 433279
rect 524420 433236 524472 433245
rect 38568 427796 38620 427848
rect 77576 427796 77628 427848
rect 503720 427796 503772 427848
rect 504272 427796 504324 427848
rect 2964 424192 3016 424244
rect 9588 424192 9640 424244
rect 524420 423691 524472 423700
rect 524420 423657 524429 423691
rect 524429 423657 524463 423691
rect 524463 423657 524472 423691
rect 524420 423648 524472 423657
rect 82820 423623 82872 423632
rect 82820 423589 82829 423623
rect 82829 423589 82863 423623
rect 82863 423589 82872 423623
rect 82820 423580 82872 423589
rect 82912 423011 82964 423020
rect 82912 422977 82921 423011
rect 82921 422977 82955 423011
rect 82955 422977 82964 423011
rect 82912 422968 82964 422977
rect 82912 418999 82964 419008
rect 82912 418965 82921 418999
rect 82921 418965 82955 418999
rect 82955 418965 82964 418999
rect 82912 418956 82964 418965
rect 503260 418208 503312 418260
rect 505468 418208 505520 418260
rect 503720 418072 503772 418124
rect 504272 418072 504324 418124
rect 514024 416712 514076 416764
rect 580172 416712 580224 416764
rect 82820 414035 82872 414044
rect 82820 414001 82829 414035
rect 82829 414001 82863 414035
rect 82863 414001 82872 414035
rect 82820 413992 82872 414001
rect 524420 413967 524472 413976
rect 524420 413933 524429 413967
rect 524429 413933 524463 413967
rect 524463 413933 524472 413967
rect 524420 413924 524472 413933
rect 503720 408484 503772 408536
rect 504272 408484 504324 408536
rect 4896 407124 4948 407176
rect 77668 407124 77720 407176
rect 82912 406283 82964 406292
rect 82912 406249 82921 406283
rect 82921 406249 82955 406283
rect 82955 406249 82964 406283
rect 82912 406240 82964 406249
rect 524420 404379 524472 404388
rect 524420 404345 524429 404379
rect 524429 404345 524463 404379
rect 524463 404345 524472 404379
rect 524420 404336 524472 404345
rect 505008 402772 505060 402824
rect 505928 402772 505980 402824
rect 83004 400664 83056 400716
rect 83004 400324 83056 400376
rect 77852 400188 77904 400240
rect 78772 400188 78824 400240
rect 83004 400188 83056 400240
rect 83004 399508 83056 399560
rect 3332 394680 3384 394732
rect 9588 394680 9640 394732
rect 524420 394655 524472 394664
rect 524420 394621 524429 394655
rect 524429 394621 524463 394655
rect 524463 394621 524472 394655
rect 524420 394612 524472 394621
rect 69664 393320 69716 393372
rect 78772 393320 78824 393372
rect 503168 393252 503220 393304
rect 579712 393252 579764 393304
rect 504548 390532 504600 390584
rect 508688 390532 508740 390584
rect 82084 387948 82136 388000
rect 82268 387948 82320 388000
rect 83004 387880 83056 387932
rect 524420 385067 524472 385076
rect 524420 385033 524429 385067
rect 524429 385033 524463 385067
rect 524463 385033 524472 385067
rect 524420 385024 524472 385033
rect 82820 384999 82872 385008
rect 82820 384965 82829 384999
rect 82829 384965 82863 384999
rect 82863 384965 82872 384999
rect 82820 384956 82872 384965
rect 3056 379516 3108 379568
rect 21364 379516 21416 379568
rect 49608 379516 49660 379568
rect 77576 379516 77628 379568
rect 504180 376728 504232 376780
rect 507768 376728 507820 376780
rect 82820 375479 82872 375488
rect 82820 375445 82829 375479
rect 82829 375445 82863 375479
rect 82863 375445 82872 375479
rect 82820 375436 82872 375445
rect 82268 375300 82320 375352
rect 82820 375300 82872 375352
rect 524420 375343 524472 375352
rect 524420 375309 524429 375343
rect 524429 375309 524463 375343
rect 524463 375309 524472 375343
rect 524420 375300 524472 375309
rect 10968 372580 11020 372632
rect 77576 372580 77628 372632
rect 83004 372716 83056 372768
rect 83004 372580 83056 372632
rect 504180 372580 504232 372632
rect 540244 372580 540296 372632
rect 83004 372444 83056 372496
rect 82268 370855 82320 370864
rect 82268 370821 82277 370855
rect 82277 370821 82311 370855
rect 82311 370821 82320 370855
rect 82268 370812 82320 370821
rect 504548 369860 504600 369912
rect 511816 369860 511868 369912
rect 83004 369316 83056 369368
rect 507584 368500 507636 368552
rect 580172 368500 580224 368552
rect 82544 366800 82596 366852
rect 82912 366800 82964 366852
rect 3608 365712 3660 365764
rect 42248 365712 42300 365764
rect 524420 365755 524472 365764
rect 524420 365721 524429 365755
rect 524429 365721 524463 365755
rect 524463 365721 524472 365755
rect 524420 365712 524472 365721
rect 82544 365236 82596 365288
rect 21364 362856 21416 362908
rect 77576 362856 77628 362908
rect 504548 362788 504600 362840
rect 508780 362788 508832 362840
rect 505928 358028 505980 358080
rect 506112 358028 506164 358080
rect 33876 357416 33928 357468
rect 74172 357416 74224 357468
rect 524420 356031 524472 356040
rect 524420 355997 524429 356031
rect 524429 355997 524463 356031
rect 524463 355997 524472 356031
rect 524420 355988 524472 355997
rect 504180 351908 504232 351960
rect 508780 351908 508832 351960
rect 524420 346443 524472 346452
rect 524420 346409 524429 346443
rect 524429 346409 524463 346443
rect 524463 346409 524472 346443
rect 524420 346400 524472 346409
rect 507676 346332 507728 346384
rect 580172 346332 580224 346384
rect 82820 344972 82872 345024
rect 82912 344972 82964 345024
rect 63408 343612 63460 343664
rect 77576 343612 77628 343664
rect 15936 342184 15988 342236
rect 73620 342184 73672 342236
rect 503444 340892 503496 340944
rect 511908 340892 511960 340944
rect 505928 339668 505980 339720
rect 506204 339668 506256 339720
rect 2964 336744 3016 336796
rect 8852 336744 8904 336796
rect 524420 336719 524472 336728
rect 524420 336685 524429 336719
rect 524429 336685 524463 336719
rect 524463 336685 524472 336719
rect 524420 336676 524472 336685
rect 17224 333888 17276 333940
rect 76472 333888 76524 333940
rect 17224 329808 17276 329860
rect 77576 329808 77628 329860
rect 504456 329808 504508 329860
rect 538864 329808 538916 329860
rect 82912 328516 82964 328568
rect 82820 328448 82872 328500
rect 79600 327972 79652 328024
rect 79968 327972 80020 328024
rect 524420 327131 524472 327140
rect 524420 327097 524429 327131
rect 524429 327097 524463 327131
rect 524463 327097 524472 327131
rect 524420 327088 524472 327097
rect 83004 326952 83056 327004
rect 3332 324232 3384 324284
rect 75276 324232 75328 324284
rect 504456 324232 504508 324284
rect 529204 324232 529256 324284
rect 505836 322872 505888 322924
rect 580172 322872 580224 322924
rect 79600 319107 79652 319116
rect 79600 319073 79609 319107
rect 79609 319073 79643 319107
rect 79643 319073 79652 319107
rect 79600 319064 79652 319073
rect 506020 318792 506072 318844
rect 506296 318792 506348 318844
rect 83004 317432 83056 317484
rect 524420 317407 524472 317416
rect 524420 317373 524429 317407
rect 524429 317373 524463 317407
rect 524463 317373 524472 317407
rect 524420 317364 524472 317373
rect 82728 316072 82780 316124
rect 82912 316072 82964 316124
rect 82636 315936 82688 315988
rect 82912 315936 82964 315988
rect 82820 313284 82872 313336
rect 82912 311312 82964 311364
rect 83004 310836 83056 310888
rect 82636 310700 82688 310752
rect 83004 310700 83056 310752
rect 83004 310564 83056 310616
rect 70216 309136 70268 309188
rect 77576 309136 77628 309188
rect 504456 309136 504508 309188
rect 506756 309136 506808 309188
rect 3332 309068 3384 309120
rect 17224 309068 17276 309120
rect 82820 309068 82872 309120
rect 524420 307819 524472 307828
rect 524420 307785 524429 307819
rect 524429 307785 524463 307819
rect 524463 307785 524472 307819
rect 524420 307776 524472 307785
rect 507032 307096 507084 307148
rect 507676 307096 507728 307148
rect 504456 306348 504508 306400
rect 564440 306348 564492 306400
rect 82820 303288 82872 303340
rect 82912 303288 82964 303340
rect 82912 303059 82964 303068
rect 82912 303025 82921 303059
rect 82921 303025 82955 303059
rect 82955 303025 82964 303059
rect 82912 303016 82964 303025
rect 82820 302880 82872 302932
rect 82912 302880 82964 302932
rect 82636 300500 82688 300552
rect 82912 300500 82964 300552
rect 511724 299412 511776 299464
rect 580172 299412 580224 299464
rect 82728 298256 82780 298308
rect 82820 298052 82872 298104
rect 524420 298095 524472 298104
rect 524420 298061 524429 298095
rect 524429 298061 524463 298095
rect 524463 298061 524472 298095
rect 524420 298052 524472 298061
rect 504456 296624 504508 296676
rect 519544 296624 519596 296676
rect 79324 296080 79376 296132
rect 3240 294720 3292 294772
rect 9496 294720 9548 294772
rect 82912 293360 82964 293412
rect 82820 291864 82872 291916
rect 82912 291771 82964 291780
rect 82912 291737 82921 291771
rect 82921 291737 82955 291771
rect 82955 291737 82964 291771
rect 82912 291728 82964 291737
rect 501972 290275 502024 290284
rect 501972 290241 501981 290275
rect 501981 290241 502015 290275
rect 502015 290241 502024 290275
rect 501972 290232 502024 290241
rect 82912 288804 82964 288856
rect 524420 288439 524472 288448
rect 524420 288405 524429 288439
rect 524429 288405 524463 288439
rect 524463 288405 524472 288439
rect 524420 288396 524472 288405
rect 82912 287759 82964 287768
rect 82912 287725 82921 287759
rect 82921 287725 82955 287759
rect 82955 287725 82964 287759
rect 82912 287716 82964 287725
rect 79324 287351 79376 287360
rect 79324 287317 79333 287351
rect 79333 287317 79367 287351
rect 79367 287317 79376 287351
rect 79324 287308 79376 287317
rect 79784 287351 79836 287360
rect 79784 287317 79793 287351
rect 79793 287317 79827 287351
rect 79827 287317 79836 287351
rect 79784 287308 79836 287317
rect 82820 286356 82872 286408
rect 82728 286220 82780 286272
rect 82912 286220 82964 286272
rect 77576 284588 77628 284640
rect 82636 284588 82688 284640
rect 82912 282251 82964 282260
rect 82912 282217 82921 282251
rect 82921 282217 82955 282251
rect 82955 282217 82964 282251
rect 82912 282208 82964 282217
rect 501972 282208 502024 282260
rect 79600 280780 79652 280832
rect 79784 280823 79836 280832
rect 79784 280789 79793 280823
rect 79793 280789 79827 280823
rect 79827 280789 79836 280823
rect 79784 280780 79836 280789
rect 57888 280168 57940 280220
rect 75644 280168 75696 280220
rect 14464 278672 14516 278724
rect 75460 278672 75512 278724
rect 501972 278400 502024 278452
rect 501972 278264 502024 278316
rect 502248 278264 502300 278316
rect 506112 277856 506164 277908
rect 502248 277788 502300 277840
rect 509056 277788 509108 277840
rect 502248 277584 502300 277636
rect 504180 277584 504232 277636
rect 82912 277423 82964 277432
rect 82912 277389 82921 277423
rect 82921 277389 82955 277423
rect 82955 277389 82964 277423
rect 82912 277380 82964 277389
rect 560944 275952 560996 276004
rect 580172 275952 580224 276004
rect 504180 274660 504232 274712
rect 545120 274660 545172 274712
rect 504180 274524 504232 274576
rect 504732 274524 504784 274576
rect 82912 273819 82964 273828
rect 82912 273785 82921 273819
rect 82921 273785 82955 273819
rect 82955 273785 82964 273819
rect 82912 273776 82964 273785
rect 501972 272756 502024 272808
rect 501972 272620 502024 272672
rect 501972 272527 502024 272536
rect 501972 272493 501981 272527
rect 501981 272493 502015 272527
rect 502015 272493 502024 272527
rect 501972 272484 502024 272493
rect 501972 272348 502024 272400
rect 79600 272144 79652 272196
rect 79968 272144 80020 272196
rect 501972 270852 502024 270904
rect 501972 270376 502024 270428
rect 82912 269764 82964 269816
rect 82912 269560 82964 269612
rect 82912 269424 82964 269476
rect 524420 269084 524472 269136
rect 524604 269084 524656 269136
rect 501972 267112 502024 267164
rect 503628 267112 503680 267164
rect 501972 266976 502024 267028
rect 82636 265888 82688 265940
rect 83004 265888 83056 265940
rect 82912 265820 82964 265872
rect 82912 265412 82964 265464
rect 2964 264936 3016 264988
rect 77300 264936 77352 264988
rect 506296 264800 506348 264852
rect 79416 264596 79468 264648
rect 80060 264596 80112 264648
rect 82912 263508 82964 263560
rect 82912 263143 82964 263152
rect 82912 263109 82921 263143
rect 82921 263109 82955 263143
rect 82955 263109 82964 263143
rect 82912 263100 82964 263109
rect 79600 260448 79652 260500
rect 79968 260448 80020 260500
rect 505836 254847 505888 254856
rect 505836 254813 505845 254847
rect 505845 254813 505879 254847
rect 505879 254813 505888 254847
rect 505836 254804 505888 254813
rect 503352 254600 503404 254652
rect 503444 253172 503496 253224
rect 503444 252968 503496 253020
rect 79600 252560 79652 252612
rect 79968 252560 80020 252612
rect 506204 251268 506256 251320
rect 3332 251200 3384 251252
rect 14464 251200 14516 251252
rect 506112 251200 506164 251252
rect 580172 251200 580224 251252
rect 505928 249772 505980 249824
rect 506296 249772 506348 249824
rect 524420 249772 524472 249824
rect 524604 249772 524656 249824
rect 41328 248412 41380 248464
rect 76012 248412 76064 248464
rect 82912 248455 82964 248464
rect 82912 248421 82921 248455
rect 82921 248421 82955 248455
rect 82955 248421 82964 248455
rect 82912 248412 82964 248421
rect 504640 246415 504692 246424
rect 504640 246381 504649 246415
rect 504649 246381 504683 246415
rect 504683 246381 504692 246415
rect 504640 246372 504692 246381
rect 82912 246304 82964 246356
rect 82820 246168 82872 246220
rect 82912 245896 82964 245948
rect 503444 245284 503496 245336
rect 503444 245148 503496 245200
rect 82912 245055 82964 245064
rect 82912 245021 82921 245055
rect 82921 245021 82955 245055
rect 82955 245021 82964 245055
rect 82912 245012 82964 245021
rect 82820 244944 82872 244996
rect 82728 243788 82780 243840
rect 82912 243788 82964 243840
rect 82912 243652 82964 243704
rect 82912 243516 82964 243568
rect 503352 242088 503404 242140
rect 503444 241884 503496 241936
rect 503628 241587 503680 241596
rect 503628 241553 503637 241587
rect 503637 241553 503671 241587
rect 503671 241553 503680 241587
rect 503628 241544 503680 241553
rect 503444 238824 503496 238876
rect 539508 238960 539560 239012
rect 549260 238960 549312 239012
rect 529940 238824 529992 238876
rect 82820 238756 82872 238808
rect 82912 238731 82964 238740
rect 82912 238697 82921 238731
rect 82921 238697 82955 238731
rect 82955 238697 82964 238731
rect 82912 238688 82964 238697
rect 82820 238620 82872 238672
rect 82452 238076 82504 238128
rect 79416 237464 79468 237516
rect 79968 237464 80020 237516
rect 3240 237328 3292 237380
rect 77760 237328 77812 237380
rect 504640 235968 504692 236020
rect 508872 235968 508924 236020
rect 503628 235220 503680 235272
rect 504640 235220 504692 235272
rect 82452 235016 82504 235068
rect 82728 235016 82780 235068
rect 81440 233699 81492 233708
rect 81440 233665 81449 233699
rect 81449 233665 81483 233699
rect 81483 233665 81492 233699
rect 81440 233656 81492 233665
rect 503536 233588 503588 233640
rect 83188 233044 83240 233096
rect 82912 232976 82964 233028
rect 82728 232840 82780 232892
rect 82912 232840 82964 232892
rect 82636 232611 82688 232620
rect 82636 232577 82645 232611
rect 82645 232577 82679 232611
rect 82679 232577 82688 232611
rect 82636 232568 82688 232577
rect 81440 230639 81492 230648
rect 81440 230605 81449 230639
rect 81449 230605 81483 230639
rect 81483 230605 81492 230639
rect 81440 230596 81492 230605
rect 524420 230460 524472 230512
rect 524604 230460 524656 230512
rect 81440 229236 81492 229288
rect 507492 229032 507544 229084
rect 580172 229032 580224 229084
rect 82728 228964 82780 229016
rect 82912 228964 82964 229016
rect 82912 228828 82964 228880
rect 81440 227876 81492 227928
rect 503628 227443 503680 227452
rect 503628 227409 503637 227443
rect 503637 227409 503671 227443
rect 503671 227409 503680 227443
rect 503628 227400 503680 227409
rect 82912 226559 82964 226568
rect 82912 226525 82921 226559
rect 82921 226525 82955 226559
rect 82955 226525 82964 226559
rect 82912 226516 82964 226525
rect 79416 225632 79468 225684
rect 79600 225632 79652 225684
rect 82912 225632 82964 225684
rect 503444 225496 503496 225548
rect 503444 224952 503496 225004
rect 519544 224952 519596 225004
rect 505836 224612 505888 224664
rect 506296 224612 506348 224664
rect 505928 224068 505980 224120
rect 506388 224068 506440 224120
rect 3332 223524 3384 223576
rect 10692 223524 10744 223576
rect 503444 221824 503496 221876
rect 508964 221824 509016 221876
rect 503628 221527 503680 221536
rect 503628 221493 503637 221527
rect 503637 221493 503671 221527
rect 503671 221493 503680 221527
rect 503628 221484 503680 221493
rect 503628 221255 503680 221264
rect 503628 221221 503637 221255
rect 503637 221221 503671 221255
rect 503671 221221 503680 221255
rect 503628 221212 503680 221221
rect 82912 220847 82964 220856
rect 82912 220813 82921 220847
rect 82921 220813 82955 220847
rect 82955 220813 82964 220847
rect 82912 220804 82964 220813
rect 503628 220192 503680 220244
rect 503536 219988 503588 220040
rect 503536 219691 503588 219700
rect 503536 219657 503545 219691
rect 503545 219657 503579 219691
rect 503579 219657 503588 219691
rect 503536 219648 503588 219657
rect 82912 219487 82964 219496
rect 82912 219453 82921 219487
rect 82921 219453 82955 219487
rect 82955 219453 82964 219487
rect 82912 219444 82964 219453
rect 506204 217991 506256 218000
rect 506204 217957 506213 217991
rect 506213 217957 506247 217991
rect 506247 217957 506256 217991
rect 506204 217948 506256 217957
rect 509056 217948 509108 218000
rect 580172 217948 580224 218000
rect 77760 216656 77812 216708
rect 80336 216656 80388 216708
rect 79600 215228 79652 215280
rect 79968 215228 80020 215280
rect 505928 214344 505980 214396
rect 506388 214344 506440 214396
rect 81532 213392 81584 213444
rect 82728 213392 82780 213444
rect 505836 212304 505888 212356
rect 506296 212304 506348 212356
rect 506296 212168 506348 212220
rect 82912 211148 82964 211200
rect 83004 211148 83056 211200
rect 503628 210740 503680 210792
rect 82636 209491 82688 209500
rect 82636 209457 82645 209491
rect 82645 209457 82679 209491
rect 82679 209457 82688 209491
rect 82636 209448 82688 209457
rect 502156 209355 502208 209364
rect 502156 209321 502165 209355
rect 502165 209321 502199 209355
rect 502199 209321 502208 209355
rect 502156 209312 502208 209321
rect 3148 208292 3200 208344
rect 10600 208292 10652 208344
rect 504824 207816 504876 207868
rect 503628 207000 503680 207052
rect 572720 207000 572772 207052
rect 79600 205640 79652 205692
rect 79968 205640 80020 205692
rect 503536 204867 503588 204876
rect 503536 204833 503545 204867
rect 503545 204833 503579 204867
rect 503579 204833 503588 204867
rect 503536 204824 503588 204833
rect 506204 204280 506256 204332
rect 580172 204280 580224 204332
rect 505836 203940 505888 203992
rect 506388 203940 506440 203992
rect 81532 202487 81584 202496
rect 81532 202453 81541 202487
rect 81541 202453 81575 202487
rect 81575 202453 81584 202487
rect 81532 202444 81584 202453
rect 79140 202104 79192 202156
rect 80336 202104 80388 202156
rect 81532 201764 81584 201816
rect 524420 201424 524472 201476
rect 524604 201424 524656 201476
rect 81532 201220 81584 201272
rect 76472 200744 76524 200796
rect 76932 200744 76984 200796
rect 81532 200268 81584 200320
rect 80336 200200 80388 200252
rect 81440 200200 81492 200252
rect 81532 200175 81584 200184
rect 81532 200141 81541 200175
rect 81541 200141 81575 200175
rect 81575 200141 81584 200175
rect 81532 200132 81584 200141
rect 505928 199631 505980 199640
rect 505928 199597 505937 199631
rect 505937 199597 505971 199631
rect 505971 199597 505980 199631
rect 505928 199588 505980 199597
rect 76932 199520 76984 199572
rect 77116 199520 77168 199572
rect 503628 199495 503680 199504
rect 503628 199461 503637 199495
rect 503637 199461 503671 199495
rect 503671 199461 503680 199495
rect 503628 199452 503680 199461
rect 503628 199316 503680 199368
rect 502156 197727 502208 197736
rect 502156 197693 502165 197727
rect 502165 197693 502199 197727
rect 502199 197693 502208 197727
rect 502156 197684 502208 197693
rect 79600 196800 79652 196852
rect 79968 196800 80020 196852
rect 503536 196188 503588 196240
rect 504824 195984 504876 196036
rect 509148 195984 509200 196036
rect 82912 195304 82964 195356
rect 82728 195279 82780 195288
rect 82728 195245 82737 195279
rect 82737 195245 82771 195279
rect 82771 195245 82780 195279
rect 82728 195236 82780 195245
rect 82912 195211 82964 195220
rect 82912 195177 82921 195211
rect 82921 195177 82955 195211
rect 82955 195177 82964 195211
rect 82912 195168 82964 195177
rect 82728 195100 82780 195152
rect 82636 195032 82688 195084
rect 82636 194896 82688 194948
rect 82912 194896 82964 194948
rect 82636 194760 82688 194812
rect 82912 194803 82964 194812
rect 82912 194769 82921 194803
rect 82921 194769 82955 194803
rect 82955 194769 82964 194803
rect 82912 194760 82964 194769
rect 503536 194352 503588 194404
rect 503076 192584 503128 192636
rect 510528 192584 510580 192636
rect 81532 192423 81584 192432
rect 81532 192389 81541 192423
rect 81541 192389 81575 192423
rect 81575 192389 81584 192423
rect 81532 192380 81584 192389
rect 81532 192176 81584 192228
rect 82912 192176 82964 192228
rect 81532 191768 81584 191820
rect 82636 191224 82688 191276
rect 76932 191088 76984 191140
rect 77116 191088 77168 191140
rect 80244 191088 80296 191140
rect 82636 191131 82688 191140
rect 82636 191097 82645 191131
rect 82645 191097 82679 191131
rect 82679 191097 82688 191131
rect 82636 191088 82688 191097
rect 76472 190952 76524 191004
rect 76932 190952 76984 191004
rect 82636 190952 82688 191004
rect 82544 190859 82596 190868
rect 82544 190825 82553 190859
rect 82553 190825 82587 190859
rect 82587 190825 82596 190859
rect 82544 190816 82596 190825
rect 82636 190748 82688 190800
rect 505928 190791 505980 190800
rect 505928 190757 505937 190791
rect 505937 190757 505971 190791
rect 505971 190757 505980 190791
rect 505928 190748 505980 190757
rect 81532 190680 81584 190732
rect 82544 190680 82596 190732
rect 82544 190476 82596 190528
rect 503076 189703 503128 189712
rect 503076 189669 503085 189703
rect 503085 189669 503119 189703
rect 503119 189669 503128 189703
rect 503076 189660 503128 189669
rect 82636 188572 82688 188624
rect 78772 188368 78824 188420
rect 82636 187212 82688 187264
rect 82636 186940 82688 186992
rect 82912 186983 82964 186992
rect 82912 186949 82921 186983
rect 82921 186949 82955 186983
rect 82955 186949 82964 186983
rect 82912 186940 82964 186949
rect 503628 186983 503680 186992
rect 503628 186949 503637 186983
rect 503637 186949 503671 186983
rect 503671 186949 503680 186983
rect 503628 186940 503680 186949
rect 82728 186668 82780 186720
rect 82912 186668 82964 186720
rect 79600 185648 79652 185700
rect 79968 185648 80020 185700
rect 82728 185691 82780 185700
rect 82728 185657 82737 185691
rect 82737 185657 82771 185691
rect 82771 185657 82780 185691
rect 82728 185648 82780 185657
rect 14464 183472 14516 183524
rect 78772 183472 78824 183524
rect 82636 182427 82688 182436
rect 82636 182393 82645 182427
rect 82645 182393 82679 182427
rect 82679 182393 82688 182427
rect 82636 182384 82688 182393
rect 504824 182180 504876 182232
rect 571984 182180 572036 182232
rect 524420 182112 524472 182164
rect 524604 182112 524656 182164
rect 503076 181772 503128 181824
rect 504824 181772 504876 181824
rect 514668 181092 514720 181144
rect 521568 181092 521620 181144
rect 533988 180956 534040 181008
rect 535460 180956 535512 181008
rect 3240 180752 3292 180804
rect 10508 180752 10560 180804
rect 503812 180140 503864 180192
rect 82636 178755 82688 178764
rect 82636 178721 82645 178755
rect 82645 178721 82679 178755
rect 82679 178721 82688 178755
rect 82636 178712 82688 178721
rect 82636 178576 82688 178628
rect 505836 178168 505888 178220
rect 82912 177216 82964 177268
rect 82912 177080 82964 177132
rect 82912 176987 82964 176996
rect 82912 176953 82921 176987
rect 82921 176953 82955 176987
rect 82955 176953 82964 176987
rect 82912 176944 82964 176953
rect 19984 176604 20036 176656
rect 79968 176604 80020 176656
rect 82912 176647 82964 176656
rect 82912 176613 82921 176647
rect 82921 176613 82955 176647
rect 82955 176613 82964 176647
rect 82912 176604 82964 176613
rect 79600 176579 79652 176588
rect 79600 176545 79609 176579
rect 79609 176545 79643 176579
rect 79643 176545 79652 176579
rect 79600 176536 79652 176545
rect 79968 175516 80020 175568
rect 82912 173136 82964 173188
rect 503076 172932 503128 172984
rect 505008 172932 505060 172984
rect 77392 171096 77444 171148
rect 78680 171096 78732 171148
rect 510068 171028 510120 171080
rect 580172 171028 580224 171080
rect 82636 170348 82688 170400
rect 82636 170255 82688 170264
rect 82636 170221 82645 170255
rect 82645 170221 82679 170255
rect 82679 170221 82688 170255
rect 82636 170212 82688 170221
rect 82636 170076 82688 170128
rect 505836 170008 505888 170060
rect 506388 170008 506440 170060
rect 503628 169235 503680 169244
rect 503628 169201 503637 169235
rect 503637 169201 503671 169235
rect 503671 169201 503680 169235
rect 503628 169192 503680 169201
rect 6828 168376 6880 168428
rect 78680 168376 78732 168428
rect 83004 168376 83056 168428
rect 83004 167220 83056 167272
rect 83004 167084 83056 167136
rect 79600 167016 79652 167068
rect 79968 167016 80020 167068
rect 83004 166676 83056 166728
rect 502984 166676 503036 166728
rect 506388 166676 506440 166728
rect 502984 166336 503036 166388
rect 83004 165996 83056 166048
rect 502984 165588 503036 165640
rect 3424 165520 3476 165572
rect 10416 165520 10468 165572
rect 503904 165520 503956 165572
rect 527180 165520 527232 165572
rect 502984 164951 503036 164960
rect 502984 164917 502993 164951
rect 502993 164917 503027 164951
rect 503027 164917 503036 164951
rect 502984 164908 503036 164917
rect 13728 164228 13780 164280
rect 78680 164228 78732 164280
rect 502984 163752 503036 163804
rect 505836 162979 505888 162988
rect 505836 162945 505845 162979
rect 505845 162945 505879 162979
rect 505879 162945 505888 162979
rect 505836 162936 505888 162945
rect 78772 162800 78824 162852
rect 502984 162800 503036 162852
rect 524420 162843 524472 162852
rect 524420 162809 524429 162843
rect 524429 162809 524463 162843
rect 524463 162809 524472 162843
rect 524420 162800 524472 162809
rect 532700 162843 532752 162852
rect 532700 162809 532709 162843
rect 532709 162809 532743 162843
rect 532743 162809 532752 162843
rect 532700 162800 532752 162809
rect 502984 162392 503036 162444
rect 81532 162120 81584 162172
rect 502984 162120 503036 162172
rect 503628 160692 503680 160744
rect 503904 160692 503956 160744
rect 501696 159103 501748 159112
rect 501696 159069 501705 159103
rect 501705 159069 501739 159103
rect 501739 159069 501748 159103
rect 501696 159060 501748 159069
rect 501880 158788 501932 158840
rect 503628 158788 503680 158840
rect 501880 158652 501932 158704
rect 507768 158652 507820 158704
rect 580172 158652 580224 158704
rect 82912 157564 82964 157616
rect 501604 157564 501656 157616
rect 507492 157564 507544 157616
rect 83004 157496 83056 157548
rect 81532 157471 81584 157480
rect 81532 157437 81541 157471
rect 81541 157437 81575 157471
rect 81575 157437 81584 157471
rect 81532 157428 81584 157437
rect 501604 157428 501656 157480
rect 78772 157292 78824 157344
rect 79600 157292 79652 157344
rect 81532 157292 81584 157344
rect 81532 157199 81584 157208
rect 81532 157165 81541 157199
rect 81541 157165 81575 157199
rect 81575 157165 81584 157199
rect 81532 157156 81584 157165
rect 83004 157020 83056 157072
rect 82912 156952 82964 157004
rect 82912 156816 82964 156868
rect 83004 156748 83056 156800
rect 82636 156340 82688 156392
rect 82912 156340 82964 156392
rect 82636 156247 82688 156256
rect 82636 156213 82645 156247
rect 82645 156213 82679 156247
rect 82679 156213 82688 156247
rect 82636 156204 82688 156213
rect 501880 155524 501932 155576
rect 501880 155388 501932 155440
rect 506296 155320 506348 155372
rect 502340 155184 502392 155236
rect 501880 155116 501932 155168
rect 506388 155116 506440 155168
rect 502340 155048 502392 155100
rect 501604 154844 501656 154896
rect 501696 154708 501748 154760
rect 501696 154572 501748 154624
rect 524420 153255 524472 153264
rect 524420 153221 524429 153255
rect 524429 153221 524463 153255
rect 524463 153221 524472 153255
rect 524420 153212 524472 153221
rect 532700 153255 532752 153264
rect 532700 153221 532709 153255
rect 532709 153221 532743 153255
rect 532743 153221 532752 153255
rect 532700 153212 532752 153221
rect 505836 152532 505888 152584
rect 82912 152507 82964 152516
rect 82912 152473 82921 152507
rect 82921 152473 82955 152507
rect 82955 152473 82964 152507
rect 82912 152464 82964 152473
rect 82912 152328 82964 152380
rect 82912 152124 82964 152176
rect 505836 152056 505888 152108
rect 501512 151920 501564 151972
rect 501512 151827 501564 151836
rect 501512 151793 501521 151827
rect 501521 151793 501555 151827
rect 501555 151793 501564 151827
rect 501512 151784 501564 151793
rect 3148 151716 3200 151768
rect 10324 151716 10376 151768
rect 501512 151648 501564 151700
rect 505836 151852 505888 151904
rect 505836 151283 505888 151292
rect 505836 151249 505845 151283
rect 505845 151249 505879 151283
rect 505879 151249 505888 151283
rect 505836 151240 505888 151249
rect 78772 151011 78824 151020
rect 78772 150977 78781 151011
rect 78781 150977 78815 151011
rect 78815 150977 78824 151011
rect 78772 150968 78824 150977
rect 56508 150424 56560 150476
rect 78772 150424 78824 150476
rect 78772 150331 78824 150340
rect 78772 150297 78781 150331
rect 78781 150297 78815 150331
rect 78815 150297 78824 150331
rect 78772 150288 78824 150297
rect 504548 148996 504600 149048
rect 502340 148928 502392 148980
rect 502340 148792 502392 148844
rect 504364 148724 504416 148776
rect 504548 148724 504600 148776
rect 504088 148588 504140 148640
rect 504364 148588 504416 148640
rect 503720 148019 503772 148028
rect 503720 147985 503729 148019
rect 503729 147985 503763 148019
rect 503763 147985 503772 148019
rect 503720 147976 503772 147985
rect 78772 147636 78824 147688
rect 79600 147636 79652 147688
rect 503720 147636 503772 147688
rect 563060 147636 563112 147688
rect 502340 147475 502392 147484
rect 502340 147441 502349 147475
rect 502349 147441 502383 147475
rect 502383 147441 502392 147475
rect 502340 147432 502392 147441
rect 504548 147364 504600 147416
rect 502340 147228 502392 147280
rect 503720 146999 503772 147008
rect 503720 146965 503729 146999
rect 503729 146965 503763 146999
rect 503763 146965 503772 146999
rect 503720 146956 503772 146965
rect 504088 146140 504140 146192
rect 504088 145979 504140 145988
rect 504088 145945 504097 145979
rect 504097 145945 504131 145979
rect 504131 145945 504140 145979
rect 504088 145936 504140 145945
rect 82912 145868 82964 145920
rect 82912 145775 82964 145784
rect 82912 145741 82921 145775
rect 82921 145741 82955 145775
rect 82955 145741 82964 145775
rect 82912 145732 82964 145741
rect 82912 145460 82964 145512
rect 504088 144440 504140 144492
rect 80244 144032 80296 144084
rect 504548 143624 504600 143676
rect 505836 143667 505888 143676
rect 505836 143633 505845 143667
rect 505845 143633 505879 143667
rect 505879 143633 505888 143667
rect 505836 143624 505888 143633
rect 524420 143531 524472 143540
rect 524420 143497 524429 143531
rect 524429 143497 524463 143531
rect 524463 143497 524472 143531
rect 524420 143488 524472 143497
rect 532700 143531 532752 143540
rect 532700 143497 532709 143531
rect 532709 143497 532743 143531
rect 532743 143497 532752 143531
rect 532700 143488 532752 143497
rect 504548 143352 504600 143404
rect 502156 141788 502208 141840
rect 501880 141652 501932 141704
rect 502156 141652 502208 141704
rect 506296 140632 506348 140684
rect 507768 140632 507820 140684
rect 501880 140496 501932 140548
rect 80152 140403 80204 140412
rect 80152 140369 80161 140403
rect 80161 140369 80195 140403
rect 80195 140369 80204 140403
rect 80152 140360 80204 140369
rect 501880 140360 501932 140412
rect 501880 140224 501932 140276
rect 501880 140088 501932 140140
rect 501880 139952 501932 140004
rect 82912 138703 82964 138712
rect 82912 138669 82921 138703
rect 82921 138669 82955 138703
rect 82955 138669 82964 138703
rect 82912 138660 82964 138669
rect 82912 138456 82964 138508
rect 502340 138252 502392 138304
rect 501880 138048 501932 138100
rect 501880 137776 501932 137828
rect 502340 137436 502392 137488
rect 82912 137300 82964 137352
rect 80428 137207 80480 137216
rect 80428 137173 80437 137207
rect 80437 137173 80471 137207
rect 80471 137173 80480 137207
rect 80428 137164 80480 137173
rect 82912 137164 82964 137216
rect 80428 137028 80480 137080
rect 82912 137071 82964 137080
rect 82912 137037 82921 137071
rect 82921 137037 82955 137071
rect 82955 137037 82964 137071
rect 82912 137028 82964 137037
rect 501880 137028 501932 137080
rect 82912 136892 82964 136944
rect 501880 136892 501932 136944
rect 80980 136867 81032 136876
rect 80980 136833 80989 136867
rect 80989 136833 81023 136867
rect 81023 136833 81032 136867
rect 80980 136824 81032 136833
rect 80980 136620 81032 136672
rect 82912 136620 82964 136672
rect 80980 136527 81032 136536
rect 80980 136493 80989 136527
rect 80989 136493 81023 136527
rect 81023 136493 81032 136527
rect 80980 136484 81032 136493
rect 503720 136280 503772 136332
rect 501696 136144 501748 136196
rect 78772 135668 78824 135720
rect 79600 135668 79652 135720
rect 501880 135507 501932 135516
rect 501880 135473 501889 135507
rect 501889 135473 501923 135507
rect 501923 135473 501932 135507
rect 501880 135464 501932 135473
rect 503720 133943 503772 133952
rect 503720 133909 503729 133943
rect 503729 133909 503763 133943
rect 503763 133909 503772 133943
rect 503720 133900 503772 133909
rect 524420 133943 524472 133952
rect 524420 133909 524429 133943
rect 524429 133909 524463 133943
rect 524463 133909 524472 133943
rect 524420 133900 524472 133909
rect 532700 133943 532752 133952
rect 532700 133909 532709 133943
rect 532709 133909 532743 133943
rect 532743 133909 532752 133943
rect 532700 133900 532752 133909
rect 78772 133288 78824 133340
rect 501696 133288 501748 133340
rect 83004 133152 83056 133204
rect 501696 133195 501748 133204
rect 501696 133161 501705 133195
rect 501705 133161 501739 133195
rect 501739 133161 501748 133195
rect 501696 133152 501748 133161
rect 82912 133016 82964 133068
rect 503628 132472 503680 132524
rect 82912 132268 82964 132320
rect 505836 131835 505888 131844
rect 505836 131801 505845 131835
rect 505845 131801 505879 131835
rect 505879 131801 505888 131835
rect 505836 131792 505888 131801
rect 506388 131835 506440 131844
rect 506388 131801 506397 131835
rect 506397 131801 506431 131835
rect 506431 131801 506440 131835
rect 506388 131792 506440 131801
rect 503720 131087 503772 131096
rect 503720 131053 503729 131087
rect 503729 131053 503763 131087
rect 503763 131053 503772 131087
rect 503720 131044 503772 131053
rect 503720 130568 503772 130620
rect 503720 129956 503772 130008
rect 82636 129072 82688 129124
rect 82728 128868 82780 128920
rect 79876 127848 79928 127900
rect 80428 127848 80480 127900
rect 503628 127780 503680 127832
rect 503628 127687 503680 127696
rect 503628 127653 503637 127687
rect 503637 127653 503671 127687
rect 503671 127653 503680 127687
rect 503628 127644 503680 127653
rect 501604 127347 501656 127356
rect 501604 127313 501613 127347
rect 501613 127313 501647 127347
rect 501647 127313 501656 127347
rect 501604 127304 501656 127313
rect 501880 127347 501932 127356
rect 501880 127313 501889 127347
rect 501889 127313 501923 127347
rect 501923 127313 501932 127347
rect 501880 127304 501932 127313
rect 502156 127347 502208 127356
rect 502156 127313 502165 127347
rect 502165 127313 502199 127347
rect 502199 127313 502208 127347
rect 502156 127304 502208 127313
rect 501880 127168 501932 127220
rect 502156 127100 502208 127152
rect 505836 126420 505888 126472
rect 506296 126420 506348 126472
rect 82360 125536 82412 125588
rect 82452 125332 82504 125384
rect 503628 124788 503680 124840
rect 501512 124763 501564 124772
rect 501512 124729 501521 124763
rect 501521 124729 501555 124763
rect 501555 124729 501564 124763
rect 501512 124720 501564 124729
rect 502616 124763 502668 124772
rect 502616 124729 502625 124763
rect 502625 124729 502659 124763
rect 502659 124729 502668 124763
rect 502616 124720 502668 124729
rect 501512 124584 501564 124636
rect 501788 124584 501840 124636
rect 507400 124108 507452 124160
rect 580172 124108 580224 124160
rect 524420 124083 524472 124092
rect 524420 124049 524429 124083
rect 524429 124049 524463 124083
rect 524463 124049 524472 124083
rect 524420 124040 524472 124049
rect 532700 124083 532752 124092
rect 532700 124049 532709 124083
rect 532709 124049 532743 124083
rect 532743 124049 532752 124083
rect 532700 124040 532752 124049
rect 501788 123836 501840 123888
rect 502156 123743 502208 123752
rect 502156 123709 502165 123743
rect 502165 123709 502199 123743
rect 502199 123709 502208 123743
rect 502156 123700 502208 123709
rect 82084 123675 82136 123684
rect 82084 123641 82093 123675
rect 82093 123641 82127 123675
rect 82127 123641 82136 123675
rect 82084 123632 82136 123641
rect 82912 123632 82964 123684
rect 82452 123607 82504 123616
rect 82452 123573 82461 123607
rect 82461 123573 82495 123607
rect 82495 123573 82504 123607
rect 82452 123564 82504 123573
rect 81992 123496 82044 123548
rect 82084 123428 82136 123480
rect 81992 123360 82044 123412
rect 82268 123360 82320 123412
rect 501604 123428 501656 123480
rect 501604 123335 501656 123344
rect 501604 123301 501613 123335
rect 501613 123301 501647 123335
rect 501647 123301 501656 123335
rect 501604 123292 501656 123301
rect 82452 123156 82504 123208
rect 82176 123088 82228 123140
rect 82544 123088 82596 123140
rect 76932 122748 76984 122800
rect 510160 122748 510212 122800
rect 83464 122680 83516 122732
rect 120540 122680 120592 122732
rect 124312 122680 124364 122732
rect 133788 122680 133840 122732
rect 286968 122680 287020 122732
rect 504364 122680 504416 122732
rect 81164 122612 81216 122664
rect 128360 122612 128412 122664
rect 143632 122612 143684 122664
rect 153108 122612 153160 122664
rect 249892 122612 249944 122664
rect 259368 122612 259420 122664
rect 284208 122612 284260 122664
rect 507032 122612 507084 122664
rect 81348 122544 81400 122596
rect 253848 122544 253900 122596
rect 503812 122544 503864 122596
rect 82360 122476 82412 122528
rect 365628 122476 365680 122528
rect 505284 122476 505336 122528
rect 83556 122408 83608 122460
rect 167000 122408 167052 122460
rect 172612 122408 172664 122460
rect 182088 122408 182140 122460
rect 241428 122408 241480 122460
rect 506756 122408 506808 122460
rect 212540 122340 212592 122392
rect 229008 122340 229060 122392
rect 80796 122272 80848 122324
rect 223580 122272 223632 122324
rect 227628 122272 227680 122324
rect 509056 122272 509108 122324
rect 80704 122204 80756 122256
rect 205640 122204 205692 122256
rect 212448 122204 212500 122256
rect 508780 122204 508832 122256
rect 82820 122136 82872 122188
rect 196072 122136 196124 122188
rect 198648 122136 198700 122188
rect 506940 122136 506992 122188
rect 78772 122068 78824 122120
rect 400128 122068 400180 122120
rect 509884 122068 509936 122120
rect 80888 122000 80940 122052
rect 99380 122000 99432 122052
rect 103520 122043 103572 122052
rect 103520 122009 103529 122043
rect 103529 122009 103563 122043
rect 103563 122009 103572 122043
rect 103520 122000 103572 122009
rect 124312 122000 124364 122052
rect 133788 122000 133840 122052
rect 143632 122000 143684 122052
rect 153108 122000 153160 122052
rect 162952 122000 163004 122052
rect 172428 122000 172480 122052
rect 172520 122000 172572 122052
rect 172796 122000 172848 122052
rect 182364 122000 182416 122052
rect 191748 122000 191800 122052
rect 240324 122000 240376 122052
rect 241520 122000 241572 122052
rect 326988 122043 327040 122052
rect 326988 122009 326997 122043
rect 326997 122009 327031 122043
rect 327031 122009 327040 122043
rect 326988 122000 327040 122009
rect 367008 122000 367060 122052
rect 503168 122000 503220 122052
rect 86868 121932 86920 121984
rect 95148 121932 95200 121984
rect 95332 121932 95384 121984
rect 101036 121932 101088 121984
rect 376852 121932 376904 121984
rect 386144 121932 386196 121984
rect 393964 121975 394016 121984
rect 393964 121941 393973 121975
rect 393973 121941 394007 121975
rect 394007 121941 394016 121975
rect 393964 121932 394016 121941
rect 404452 121932 404504 121984
rect 413928 121932 413980 121984
rect 415768 121932 415820 121984
rect 424968 121932 425020 121984
rect 440148 121932 440200 121984
rect 511540 121932 511592 121984
rect 95240 121864 95292 121916
rect 105360 121864 105412 121916
rect 469128 121864 469180 121916
rect 503444 121864 503496 121916
rect 79692 121796 79744 121848
rect 84936 121796 84988 121848
rect 90640 121796 90692 121848
rect 129740 121796 129792 121848
rect 338120 121796 338172 121848
rect 342996 121796 343048 121848
rect 484308 121796 484360 121848
rect 505376 121796 505428 121848
rect 78864 121728 78916 121780
rect 92296 121728 92348 121780
rect 123024 121728 123076 121780
rect 330944 121728 330996 121780
rect 336648 121728 336700 121780
rect 480168 121728 480220 121780
rect 78220 121660 78272 121712
rect 111064 121660 111116 121712
rect 338120 121703 338172 121712
rect 338120 121669 338129 121703
rect 338129 121669 338163 121703
rect 338163 121669 338172 121703
rect 338120 121660 338172 121669
rect 491300 121660 491352 121712
rect 492312 121660 492364 121712
rect 493324 121660 493376 121712
rect 498476 121660 498528 121712
rect 499304 121660 499356 121712
rect 507308 121660 507360 121712
rect 9588 121592 9640 121644
rect 175280 121592 175332 121644
rect 399392 121592 399444 121644
rect 506848 121592 506900 121644
rect 3516 121524 3568 121576
rect 277768 121524 277820 121576
rect 377864 121524 377916 121576
rect 507216 121524 507268 121576
rect 79692 121456 79744 121508
rect 445852 121456 445904 121508
rect 496084 121456 496136 121508
rect 507308 121456 507360 121508
rect 510528 121456 510580 121508
rect 9312 121388 9364 121440
rect 494520 121388 494572 121440
rect 499396 121388 499448 121440
rect 509884 121388 509936 121440
rect 511632 121388 511684 121440
rect 8852 121320 8904 121372
rect 454040 121320 454092 121372
rect 456708 121320 456760 121372
rect 502892 121320 502944 121372
rect 42248 121252 42300 121304
rect 466000 121252 466052 121304
rect 488448 121252 488500 121304
rect 499764 121252 499816 121304
rect 24768 121184 24820 121236
rect 427912 121184 427964 121236
rect 431868 121184 431920 121236
rect 502800 121252 502852 121304
rect 499948 121184 500000 121236
rect 501788 121184 501840 121236
rect 3700 121116 3752 121168
rect 173072 121116 173124 121168
rect 189632 121116 189684 121168
rect 580632 121116 580684 121168
rect 85028 121048 85080 121100
rect 392216 121048 392268 121100
rect 500040 121048 500092 121100
rect 511816 121048 511868 121100
rect 33784 120980 33836 121032
rect 127808 120980 127860 121032
rect 144368 120980 144420 121032
rect 506112 120980 506164 121032
rect 3424 120912 3476 120964
rect 146760 120912 146812 120964
rect 165896 120912 165948 120964
rect 505744 120912 505796 120964
rect 9404 120844 9456 120896
rect 337384 120844 337436 120896
rect 349068 120844 349120 120896
rect 511908 120844 511960 120896
rect 42156 120776 42208 120828
rect 163504 120776 163556 120828
rect 239680 120776 239732 120828
rect 506204 120776 506256 120828
rect 77300 120708 77352 120760
rect 313464 120708 313516 120760
rect 318248 120708 318300 120760
rect 580448 120708 580500 120760
rect 79048 120640 79100 120692
rect 150624 120640 150676 120692
rect 274548 120640 274600 120692
rect 84016 120572 84068 120624
rect 118424 120572 118476 120624
rect 284944 120572 284996 120624
rect 498936 120640 498988 120692
rect 507124 120640 507176 120692
rect 506664 120572 506716 120624
rect 80980 120504 81032 120556
rect 304908 120504 304960 120556
rect 509700 120504 509752 120556
rect 106464 120436 106516 120488
rect 329748 120436 329800 120488
rect 393228 120368 393280 120420
rect 510436 120368 510488 120420
rect 31116 120300 31168 120352
rect 401600 120300 401652 120352
rect 508504 120300 508556 120352
rect 15108 120028 15160 120080
rect 137192 120028 137244 120080
rect 149152 120028 149204 120080
rect 150348 120028 150400 120080
rect 199200 120028 199252 120080
rect 200028 120028 200080 120080
rect 201592 120028 201644 120080
rect 225052 120028 225104 120080
rect 244464 120028 244516 120080
rect 245568 120028 245620 120080
rect 251088 120028 251140 120080
rect 496912 120028 496964 120080
rect 84752 119960 84804 120012
rect 242900 119960 242952 120012
rect 261208 119960 261260 120012
rect 262128 119960 262180 120012
rect 265808 119960 265860 120012
rect 22008 119892 22060 119944
rect 156328 119892 156380 119944
rect 179328 119892 179380 119944
rect 430304 119892 430356 119944
rect 437480 119892 437532 119944
rect 438768 119892 438820 119944
rect 461216 119892 461268 119944
rect 508136 119892 508188 119944
rect 17224 119824 17276 119876
rect 270592 119824 270644 119876
rect 275376 119824 275428 119876
rect 522304 119824 522356 119876
rect 71688 119756 71740 119808
rect 234896 119756 234948 119808
rect 242072 119756 242124 119808
rect 495440 119756 495492 119808
rect 51816 119688 51868 119740
rect 306472 119688 306524 119740
rect 311072 119688 311124 119740
rect 349160 119688 349212 119740
rect 352564 119688 352616 119740
rect 356336 119688 356388 119740
rect 363512 119688 363564 119740
rect 519636 119688 519688 119740
rect 59268 119620 59320 119672
rect 227720 119620 227772 119672
rect 230112 119620 230164 119672
rect 489920 119620 489972 119672
rect 491208 119620 491260 119672
rect 80612 119552 80664 119604
rect 103888 119552 103940 119604
rect 104808 119552 104860 119604
rect 106280 119552 106332 119604
rect 107476 119552 107528 119604
rect 382648 119552 382700 119604
rect 391848 119552 391900 119604
rect 473176 119552 473228 119604
rect 479524 119552 479576 119604
rect 509976 119552 510028 119604
rect 28908 119484 28960 119536
rect 194416 119484 194468 119536
rect 211160 119484 211212 119536
rect 212356 119484 212408 119536
rect 509148 119484 509200 119536
rect 46296 119416 46348 119468
rect 82728 119459 82780 119468
rect 20628 119348 20680 119400
rect 82728 119425 82737 119459
rect 82737 119425 82771 119459
rect 82771 119425 82780 119459
rect 82728 119416 82780 119425
rect 425520 119416 425572 119468
rect 463608 119416 463660 119468
rect 471244 119416 471296 119468
rect 476764 119416 476816 119468
rect 510344 119416 510396 119468
rect 91928 119348 91980 119400
rect 94320 119348 94372 119400
rect 473360 119348 473412 119400
rect 492680 119348 492732 119400
rect 571340 119348 571392 119400
rect 38476 119280 38528 119332
rect 151544 119280 151596 119332
rect 365904 119280 365956 119332
rect 373080 119280 373132 119332
rect 373908 119280 373960 119332
rect 380256 119280 380308 119332
rect 441712 119280 441764 119332
rect 467748 119280 467800 119332
rect 480352 119280 480404 119332
rect 487068 119280 487120 119332
rect 501512 119280 501564 119332
rect 83648 119212 83700 119264
rect 87328 119212 87380 119264
rect 102048 119212 102100 119264
rect 113456 119212 113508 119264
rect 114468 119212 114520 119264
rect 232504 119212 232556 119264
rect 240048 119212 240100 119264
rect 449256 119212 449308 119264
rect 487528 119212 487580 119264
rect 92388 119144 92440 119196
rect 208768 119144 208820 119196
rect 211068 119144 211120 119196
rect 218336 119144 218388 119196
rect 219348 119144 219400 119196
rect 222936 119144 222988 119196
rect 416780 119144 416832 119196
rect 500868 119144 500920 119196
rect 91008 119076 91060 119128
rect 196808 119076 196860 119128
rect 206376 119076 206428 119128
rect 396080 119076 396132 119128
rect 402244 119076 402296 119128
rect 451648 119076 451700 119128
rect 78588 119008 78640 119060
rect 161112 119008 161164 119060
rect 180064 119008 180116 119060
rect 360200 119008 360252 119060
rect 384948 119008 385000 119060
rect 447048 119008 447100 119060
rect 106188 118940 106240 118992
rect 203984 118940 204036 118992
rect 233148 118940 233200 118992
rect 301688 118940 301740 118992
rect 313924 118940 313976 118992
rect 332600 118940 332652 118992
rect 355968 118940 356020 118992
rect 509608 118940 509660 118992
rect 72976 118872 73028 118924
rect 125416 118872 125468 118924
rect 246948 118872 247000 118924
rect 375472 118872 375524 118924
rect 407028 118872 407080 118924
rect 423128 118872 423180 118924
rect 113088 118804 113140 118856
rect 120632 118804 120684 118856
rect 169760 118804 169812 118856
rect 222108 118804 222160 118856
rect 237196 118804 237248 118856
rect 304080 118804 304132 118856
rect 433340 118804 433392 118856
rect 435088 118804 435140 118856
rect 436008 118804 436060 118856
rect 107568 118736 107620 118788
rect 132408 118736 132460 118788
rect 201408 118736 201460 118788
rect 268200 118736 268252 118788
rect 280160 118736 280212 118788
rect 310520 118736 310572 118788
rect 344560 118736 344612 118788
rect 419540 118736 419592 118788
rect 225328 118668 225380 118720
rect 226248 118668 226300 118720
rect 156052 118643 156104 118652
rect 156052 118609 156061 118643
rect 156061 118609 156095 118643
rect 156095 118609 156104 118643
rect 156052 118600 156104 118609
rect 263600 118668 263652 118720
rect 307024 118668 307076 118720
rect 315856 118668 315908 118720
rect 349344 118668 349396 118720
rect 368296 118668 368348 118720
rect 369952 118668 370004 118720
rect 81624 118532 81676 118584
rect 258172 118532 258224 118584
rect 502064 118575 502116 118584
rect 502064 118541 502073 118575
rect 502073 118541 502107 118575
rect 502107 118541 502116 118575
rect 502064 118532 502116 118541
rect 83280 118464 83332 118516
rect 267740 118464 267792 118516
rect 81808 118396 81860 118448
rect 269120 118396 269172 118448
rect 83096 118328 83148 118380
rect 287060 118328 287112 118380
rect 500224 118328 500276 118380
rect 504548 118328 504600 118380
rect 80520 118260 80572 118312
rect 305000 118260 305052 118312
rect 413560 118260 413612 118312
rect 413928 118260 413980 118312
rect 422208 118260 422260 118312
rect 503536 118260 503588 118312
rect 78956 118192 79008 118244
rect 320180 118192 320232 118244
rect 398748 118192 398800 118244
rect 503260 118192 503312 118244
rect 82544 118124 82596 118176
rect 84844 118124 84896 118176
rect 82176 118056 82228 118108
rect 244372 118124 244424 118176
rect 249708 118124 249760 118176
rect 503352 118124 503404 118176
rect 132592 118056 132644 118108
rect 220728 118056 220780 118108
rect 504272 118056 504324 118108
rect 81992 117988 82044 118040
rect 514760 117988 514812 118040
rect 82084 117920 82136 117972
rect 536932 117920 536984 117972
rect 500132 117784 500184 117836
rect 492312 117308 492364 117360
rect 496728 117308 496780 117360
rect 490564 117104 490616 117156
rect 493508 117104 493560 117156
rect 82452 116764 82504 116816
rect 161480 116764 161532 116816
rect 322756 116764 322808 116816
rect 511172 116764 511224 116816
rect 83832 116696 83884 116748
rect 372528 116696 372580 116748
rect 401508 116696 401560 116748
rect 502984 116696 503036 116748
rect 136548 116628 136600 116680
rect 505008 116628 505060 116680
rect 79140 116560 79192 116612
rect 451280 116560 451332 116612
rect 415492 116084 415544 116136
rect 415952 116084 416004 116136
rect 161296 116059 161348 116068
rect 161296 116025 161305 116059
rect 161305 116025 161339 116059
rect 161339 116025 161348 116059
rect 161296 116016 161348 116025
rect 153016 115948 153068 116000
rect 153108 115948 153160 116000
rect 509608 115948 509660 116000
rect 511448 115948 511500 116000
rect 131212 115923 131264 115932
rect 131212 115889 131221 115923
rect 131221 115889 131255 115923
rect 131255 115889 131264 115923
rect 131212 115880 131264 115889
rect 155868 115880 155920 115932
rect 156144 115880 156196 115932
rect 161296 115923 161348 115932
rect 161296 115889 161305 115923
rect 161305 115889 161339 115923
rect 161339 115889 161348 115923
rect 161296 115880 161348 115889
rect 179328 115923 179380 115932
rect 179328 115889 179337 115923
rect 179337 115889 179371 115923
rect 179371 115889 179380 115923
rect 179328 115880 179380 115889
rect 244280 115923 244332 115932
rect 244280 115889 244289 115923
rect 244289 115889 244323 115923
rect 244323 115889 244332 115923
rect 244280 115880 244332 115889
rect 258080 115923 258132 115932
rect 258080 115889 258089 115923
rect 258089 115889 258123 115923
rect 258123 115889 258132 115923
rect 258080 115880 258132 115889
rect 445852 115923 445904 115932
rect 445852 115889 445861 115923
rect 445861 115889 445895 115923
rect 445895 115889 445904 115923
rect 445852 115880 445904 115889
rect 153016 115855 153068 115864
rect 153016 115821 153025 115855
rect 153025 115821 153059 115855
rect 153059 115821 153068 115855
rect 153016 115812 153068 115821
rect 511632 115855 511684 115864
rect 511632 115821 511641 115855
rect 511641 115821 511675 115855
rect 511675 115821 511684 115855
rect 511632 115812 511684 115821
rect 278688 115404 278740 115456
rect 502708 115404 502760 115456
rect 504916 115336 504968 115388
rect 183468 115268 183520 115320
rect 504640 115268 504692 115320
rect 80336 115200 80388 115252
rect 552020 115200 552072 115252
rect 393320 115132 393372 115184
rect 394608 115132 394660 115184
rect 500316 114656 500368 114708
rect 507308 114656 507360 114708
rect 110420 114563 110472 114572
rect 110420 114529 110429 114563
rect 110429 114529 110463 114563
rect 110463 114529 110472 114563
rect 110420 114520 110472 114529
rect 186228 114563 186280 114572
rect 186228 114529 186237 114563
rect 186237 114529 186271 114563
rect 186271 114529 186280 114563
rect 186228 114520 186280 114529
rect 272984 114520 273036 114572
rect 273076 114520 273128 114572
rect 524420 114563 524472 114572
rect 524420 114529 524429 114563
rect 524429 114529 524463 114563
rect 524463 114529 524472 114563
rect 524420 114520 524472 114529
rect 532700 114563 532752 114572
rect 532700 114529 532709 114563
rect 532709 114529 532743 114563
rect 532743 114529 532752 114563
rect 532700 114520 532752 114529
rect 155868 114495 155920 114504
rect 155868 114461 155877 114495
rect 155877 114461 155911 114495
rect 155911 114461 155920 114495
rect 155868 114452 155920 114461
rect 511632 114452 511684 114504
rect 110420 114427 110472 114436
rect 110420 114393 110429 114427
rect 110429 114393 110463 114427
rect 110463 114393 110472 114427
rect 110420 114384 110472 114393
rect 487528 114112 487580 114164
rect 492312 114112 492364 114164
rect 348976 113840 349028 113892
rect 502340 113840 502392 113892
rect 79232 113772 79284 113824
rect 454040 113772 454092 113824
rect 82728 113203 82780 113212
rect 82728 113169 82737 113203
rect 82737 113169 82771 113203
rect 82771 113169 82780 113203
rect 82728 113160 82780 113169
rect 505836 113160 505888 113212
rect 506296 113160 506348 113212
rect 89536 113092 89588 113144
rect 89628 113024 89680 113076
rect 110328 112412 110380 112464
rect 505928 112412 505980 112464
rect 481732 111800 481784 111852
rect 487528 111800 487580 111852
rect 506940 111800 506992 111852
rect 509608 111800 509660 111852
rect 80060 111775 80112 111784
rect 80060 111741 80069 111775
rect 80069 111741 80103 111775
rect 80103 111741 80112 111775
rect 80060 111732 80112 111741
rect 82636 111732 82688 111784
rect 82728 111732 82780 111784
rect 83372 111732 83424 111784
rect 83740 111732 83792 111784
rect 83832 111732 83884 111784
rect 83464 111664 83516 111716
rect 508136 111392 508188 111444
rect 509884 111392 509936 111444
rect 304908 111299 304960 111308
rect 304908 111265 304917 111299
rect 304917 111265 304951 111299
rect 304951 111265 304960 111299
rect 304908 111256 304960 111265
rect 440148 111256 440200 111308
rect 295340 111188 295392 111240
rect 304816 111188 304868 111240
rect 372712 111188 372764 111240
rect 382096 111188 382148 111240
rect 411260 111188 411312 111240
rect 420736 111188 420788 111240
rect 81072 111120 81124 111172
rect 263600 111120 263652 111172
rect 276020 111120 276072 111172
rect 285496 111120 285548 111172
rect 314660 111120 314712 111172
rect 323584 111120 323636 111172
rect 353300 111120 353352 111172
rect 362776 111120 362828 111172
rect 430580 111120 430632 111172
rect 440056 111120 440108 111172
rect 79324 111052 79376 111104
rect 440148 111052 440200 111104
rect 378140 111027 378192 111036
rect 378140 110993 378149 111027
rect 378149 110993 378183 111027
rect 378183 110993 378192 111027
rect 378140 110984 378192 110993
rect 117688 110372 117740 110424
rect 505836 109828 505888 109880
rect 506112 109828 506164 109880
rect 481364 109760 481416 109812
rect 481732 109760 481784 109812
rect 85488 109692 85540 109744
rect 505652 109692 505704 109744
rect 272984 109148 273036 109200
rect 3240 108944 3292 108996
rect 508964 108944 509016 108996
rect 121368 108876 121420 108928
rect 121552 108876 121604 108928
rect 153016 108919 153068 108928
rect 153016 108885 153025 108919
rect 153025 108885 153059 108919
rect 153059 108885 153068 108919
rect 153016 108876 153068 108885
rect 161296 108919 161348 108928
rect 161296 108885 161305 108919
rect 161305 108885 161339 108919
rect 161339 108885 161348 108919
rect 161296 108876 161348 108885
rect 272892 108919 272944 108928
rect 272892 108885 272901 108919
rect 272901 108885 272935 108919
rect 272935 108885 272944 108919
rect 272892 108876 272944 108885
rect 479616 107448 479668 107500
rect 481364 107448 481416 107500
rect 179328 106403 179380 106412
rect 179328 106369 179337 106403
rect 179337 106369 179371 106403
rect 179371 106369 179380 106403
rect 179328 106360 179380 106369
rect 131212 106335 131264 106344
rect 131212 106301 131221 106335
rect 131221 106301 131255 106335
rect 131255 106301 131264 106335
rect 131212 106292 131264 106301
rect 244280 106335 244332 106344
rect 244280 106301 244289 106335
rect 244289 106301 244323 106335
rect 244323 106301 244332 106335
rect 244280 106292 244332 106301
rect 445852 106335 445904 106344
rect 445852 106301 445861 106335
rect 445861 106301 445895 106335
rect 445895 106301 445904 106335
rect 445852 106292 445904 106301
rect 505744 106292 505796 106344
rect 508136 106292 508188 106344
rect 304908 105519 304960 105528
rect 304908 105485 304917 105519
rect 304917 105485 304951 105519
rect 304951 105485 304960 105519
rect 304908 105476 304960 105485
rect 351736 104932 351788 104984
rect 351920 104932 351972 104984
rect 110420 104907 110472 104916
rect 110420 104873 110429 104907
rect 110429 104873 110463 104907
rect 110463 104873 110472 104907
rect 110420 104864 110472 104873
rect 156052 104864 156104 104916
rect 511540 104907 511592 104916
rect 511540 104873 511549 104907
rect 511549 104873 511583 104907
rect 511583 104873 511592 104907
rect 511540 104864 511592 104873
rect 179328 104839 179380 104848
rect 179328 104805 179337 104839
rect 179337 104805 179371 104839
rect 179371 104805 179380 104839
rect 179328 104796 179380 104805
rect 186228 104839 186280 104848
rect 186228 104805 186237 104839
rect 186237 104805 186271 104839
rect 186271 104805 186280 104839
rect 186228 104796 186280 104805
rect 220728 104839 220780 104848
rect 220728 104805 220737 104839
rect 220737 104805 220771 104839
rect 220771 104805 220780 104839
rect 220728 104796 220780 104805
rect 223580 104839 223632 104848
rect 223580 104805 223589 104839
rect 223589 104805 223623 104839
rect 223623 104805 223632 104839
rect 223580 104796 223632 104805
rect 351736 104839 351788 104848
rect 351736 104805 351745 104839
rect 351745 104805 351779 104839
rect 351779 104805 351788 104839
rect 351736 104796 351788 104805
rect 524420 104839 524472 104848
rect 524420 104805 524429 104839
rect 524429 104805 524463 104839
rect 524463 104805 524472 104839
rect 524420 104796 524472 104805
rect 532700 104839 532752 104848
rect 532700 104805 532709 104839
rect 532709 104805 532743 104839
rect 532743 104805 532752 104839
rect 532700 104796 532752 104805
rect 156144 104728 156196 104780
rect 511632 104728 511684 104780
rect 489184 103096 489236 103148
rect 490564 103096 490616 103148
rect 258080 102935 258132 102944
rect 258080 102901 258089 102935
rect 258089 102901 258123 102935
rect 258123 102901 258132 102935
rect 258080 102892 258132 102901
rect 80060 102187 80112 102196
rect 80060 102153 80069 102187
rect 80069 102153 80103 102187
rect 80103 102153 80112 102187
rect 80060 102144 80112 102153
rect 266084 102144 266136 102196
rect 266268 102144 266320 102196
rect 501236 102076 501288 102128
rect 506940 102144 506992 102196
rect 117504 100827 117556 100836
rect 117504 100793 117513 100827
rect 117513 100793 117547 100827
rect 117547 100793 117556 100827
rect 117504 100784 117556 100793
rect 117504 100648 117556 100700
rect 117780 100648 117832 100700
rect 497464 99832 497516 99884
rect 500316 99832 500368 99884
rect 299296 99424 299348 99476
rect 121460 99356 121512 99408
rect 121644 99356 121696 99408
rect 161204 99356 161256 99408
rect 161388 99356 161440 99408
rect 79692 99288 79744 99340
rect 79968 99288 80020 99340
rect 117780 99288 117832 99340
rect 299296 99288 299348 99340
rect 272616 99220 272668 99272
rect 272984 99220 273036 99272
rect 475384 98404 475436 98456
rect 479616 98404 479668 98456
rect 500316 97996 500368 98048
rect 501236 97996 501288 98048
rect 436100 96747 436152 96756
rect 436100 96713 436109 96747
rect 436109 96713 436143 96747
rect 436143 96713 436152 96747
rect 436100 96704 436152 96713
rect 131212 96611 131264 96620
rect 131212 96577 131221 96611
rect 131221 96577 131255 96611
rect 131255 96577 131264 96611
rect 131212 96568 131264 96577
rect 161204 96568 161256 96620
rect 161296 96568 161348 96620
rect 244280 96611 244332 96620
rect 244280 96577 244289 96611
rect 244289 96577 244323 96611
rect 244323 96577 244332 96611
rect 244280 96568 244332 96577
rect 258080 96611 258132 96620
rect 258080 96577 258089 96611
rect 258089 96577 258123 96611
rect 258123 96577 258132 96611
rect 258080 96568 258132 96577
rect 272984 96611 273036 96620
rect 272984 96577 272993 96611
rect 272993 96577 273027 96611
rect 273027 96577 273036 96611
rect 272984 96568 273036 96577
rect 289544 96568 289596 96620
rect 289728 96568 289780 96620
rect 299296 96611 299348 96620
rect 299296 96577 299305 96611
rect 299305 96577 299339 96611
rect 299339 96577 299348 96611
rect 299296 96568 299348 96577
rect 436100 96568 436152 96620
rect 436284 96568 436336 96620
rect 445852 96611 445904 96620
rect 445852 96577 445861 96611
rect 445861 96577 445895 96611
rect 445895 96577 445904 96611
rect 445852 96568 445904 96577
rect 511724 96543 511776 96552
rect 511724 96509 511733 96543
rect 511733 96509 511767 96543
rect 511767 96509 511776 96543
rect 511724 96500 511776 96509
rect 120264 95276 120316 95328
rect 120356 95276 120408 95328
rect 152924 95208 152976 95260
rect 153108 95208 153160 95260
rect 156236 95251 156288 95260
rect 156236 95217 156245 95251
rect 156245 95217 156279 95251
rect 156279 95217 156288 95251
rect 156236 95208 156288 95217
rect 186228 95251 186280 95260
rect 186228 95217 186237 95251
rect 186237 95217 186271 95251
rect 186271 95217 186280 95251
rect 186228 95208 186280 95217
rect 220728 95251 220780 95260
rect 220728 95217 220737 95251
rect 220737 95217 220771 95251
rect 220771 95217 220780 95251
rect 220728 95208 220780 95217
rect 223580 95251 223632 95260
rect 223580 95217 223589 95251
rect 223589 95217 223623 95251
rect 223623 95217 223632 95251
rect 223580 95208 223632 95217
rect 378140 95251 378192 95260
rect 378140 95217 378149 95251
rect 378149 95217 378183 95251
rect 378183 95217 378192 95251
rect 378140 95208 378192 95217
rect 524420 95251 524472 95260
rect 524420 95217 524429 95251
rect 524429 95217 524463 95251
rect 524463 95217 524472 95251
rect 524420 95208 524472 95217
rect 532700 95251 532752 95260
rect 532700 95217 532709 95251
rect 532709 95217 532743 95251
rect 532743 95217 532752 95251
rect 532700 95208 532752 95217
rect 110420 95183 110472 95192
rect 110420 95149 110429 95183
rect 110429 95149 110463 95183
rect 110463 95149 110472 95183
rect 110420 95140 110472 95149
rect 220544 95183 220596 95192
rect 220544 95149 220553 95183
rect 220553 95149 220587 95183
rect 220587 95149 220596 95183
rect 220544 95140 220596 95149
rect 500224 93891 500276 93900
rect 500224 93857 500233 93891
rect 500233 93857 500267 93891
rect 500267 93857 500276 93891
rect 500224 93848 500276 93857
rect 3424 93780 3476 93832
rect 33876 93780 33928 93832
rect 120264 92420 120316 92472
rect 120356 92420 120408 92472
rect 474004 91060 474056 91112
rect 475384 91060 475436 91112
rect 79324 90992 79376 91044
rect 79968 90992 80020 91044
rect 117504 89743 117556 89752
rect 117504 89709 117513 89743
rect 117513 89709 117547 89743
rect 117547 89709 117556 89743
rect 117504 89700 117556 89709
rect 121460 89700 121512 89752
rect 121644 89700 121696 89752
rect 351736 89675 351788 89684
rect 351736 89641 351745 89675
rect 351745 89641 351779 89675
rect 351779 89641 351788 89675
rect 351736 89632 351788 89641
rect 179328 87091 179380 87100
rect 179328 87057 179337 87091
rect 179337 87057 179371 87091
rect 179371 87057 179380 87091
rect 179328 87048 179380 87057
rect 131212 87023 131264 87032
rect 131212 86989 131221 87023
rect 131221 86989 131255 87023
rect 131255 86989 131264 87023
rect 131212 86980 131264 86989
rect 244280 87023 244332 87032
rect 244280 86989 244289 87023
rect 244289 86989 244323 87023
rect 244323 86989 244332 87023
rect 244280 86980 244332 86989
rect 258080 87023 258132 87032
rect 258080 86989 258089 87023
rect 258089 86989 258123 87023
rect 258123 86989 258132 87023
rect 258080 86980 258132 86989
rect 272984 87023 273036 87032
rect 272984 86989 272993 87023
rect 272993 86989 273027 87023
rect 273027 86989 273036 87023
rect 272984 86980 273036 86989
rect 299296 87023 299348 87032
rect 299296 86989 299305 87023
rect 299305 86989 299339 87023
rect 299339 86989 299348 87023
rect 299296 86980 299348 86989
rect 445852 87023 445904 87032
rect 445852 86989 445861 87023
rect 445861 86989 445895 87023
rect 445895 86989 445904 87023
rect 445852 86980 445904 86989
rect 511632 86980 511684 87032
rect 511724 86980 511776 87032
rect 436100 86955 436152 86964
rect 436100 86921 436109 86955
rect 436109 86921 436143 86955
rect 436143 86921 436152 86955
rect 436100 86912 436152 86921
rect 487160 86708 487212 86760
rect 489184 86708 489236 86760
rect 135076 86232 135128 86284
rect 504456 86232 504508 86284
rect 110420 85663 110472 85672
rect 110420 85629 110429 85663
rect 110429 85629 110463 85663
rect 110463 85629 110472 85663
rect 110420 85620 110472 85629
rect 161020 85552 161072 85604
rect 161296 85552 161348 85604
rect 220544 85595 220596 85604
rect 220544 85561 220553 85595
rect 220553 85561 220587 85595
rect 220587 85561 220596 85595
rect 220544 85552 220596 85561
rect 110420 85484 110472 85536
rect 110512 85484 110564 85536
rect 179328 85527 179380 85536
rect 179328 85493 179337 85527
rect 179337 85493 179371 85527
rect 179371 85493 179380 85527
rect 179328 85484 179380 85493
rect 186228 85527 186280 85536
rect 186228 85493 186237 85527
rect 186237 85493 186271 85527
rect 186271 85493 186280 85527
rect 186228 85484 186280 85493
rect 220728 85484 220780 85536
rect 223580 85527 223632 85536
rect 223580 85493 223589 85527
rect 223589 85493 223623 85527
rect 223623 85493 223632 85527
rect 223580 85484 223632 85493
rect 378140 85527 378192 85536
rect 378140 85493 378149 85527
rect 378149 85493 378183 85527
rect 378183 85493 378192 85527
rect 378140 85484 378192 85493
rect 511540 85527 511592 85536
rect 511540 85493 511549 85527
rect 511549 85493 511583 85527
rect 511583 85493 511592 85527
rect 511540 85484 511592 85493
rect 524420 85527 524472 85536
rect 524420 85493 524429 85527
rect 524429 85493 524463 85527
rect 524463 85493 524472 85527
rect 524420 85484 524472 85493
rect 532700 85527 532752 85536
rect 532700 85493 532709 85527
rect 532709 85493 532743 85527
rect 532743 85493 532752 85527
rect 532700 85484 532752 85493
rect 497556 84464 497608 84516
rect 500316 84464 500368 84516
rect 80244 83444 80296 83496
rect 444472 83444 444524 83496
rect 120356 82875 120408 82884
rect 120356 82841 120365 82875
rect 120365 82841 120399 82875
rect 120399 82841 120408 82875
rect 120356 82832 120408 82841
rect 80060 82807 80112 82816
rect 80060 82773 80069 82807
rect 80069 82773 80103 82807
rect 80103 82773 80112 82807
rect 80060 82764 80112 82773
rect 210976 82084 211028 82136
rect 504732 82084 504784 82136
rect 79324 81880 79376 81932
rect 79968 81880 80020 81932
rect 117504 81404 117556 81456
rect 117596 81404 117648 81456
rect 120356 81447 120408 81456
rect 120356 81413 120365 81447
rect 120365 81413 120399 81447
rect 120399 81413 120408 81447
rect 120356 81404 120408 81413
rect 472348 81404 472400 81456
rect 474004 81404 474056 81456
rect 486148 81404 486200 81456
rect 487160 81404 487212 81456
rect 117596 80112 117648 80164
rect 120356 80112 120408 80164
rect 220544 80112 220596 80164
rect 272984 80112 273036 80164
rect 299296 80112 299348 80164
rect 351736 80112 351788 80164
rect 506020 80112 506072 80164
rect 117504 79976 117556 80028
rect 120264 79976 120316 80028
rect 220544 79976 220596 80028
rect 272984 79976 273036 80028
rect 299296 79976 299348 80028
rect 351736 79976 351788 80028
rect 506020 79976 506072 80028
rect 503720 79636 503772 79688
rect 505744 79636 505796 79688
rect 485044 79160 485096 79212
rect 486148 79160 486200 79212
rect 495992 78684 496044 78736
rect 497464 78684 497516 78736
rect 505928 78004 505980 78056
rect 506112 78004 506164 78056
rect 289728 77528 289780 77580
rect 289728 77256 289780 77308
rect 436100 77299 436152 77308
rect 436100 77265 436109 77299
rect 436109 77265 436143 77299
rect 436143 77265 436152 77299
rect 436100 77256 436152 77265
rect 500224 77299 500276 77308
rect 500224 77265 500233 77299
rect 500233 77265 500267 77299
rect 500267 77265 500276 77299
rect 500224 77256 500276 77265
rect 76564 77188 76616 77240
rect 580172 77188 580224 77240
rect 244280 77163 244332 77172
rect 244280 77129 244289 77163
rect 244289 77129 244323 77163
rect 244323 77129 244332 77163
rect 244280 77120 244332 77129
rect 258080 77163 258132 77172
rect 258080 77129 258089 77163
rect 258089 77129 258123 77163
rect 258123 77129 258132 77163
rect 258080 77120 258132 77129
rect 445852 77163 445904 77172
rect 445852 77129 445861 77163
rect 445861 77129 445895 77163
rect 445895 77129 445904 77163
rect 445852 77120 445904 77129
rect 470692 77120 470744 77172
rect 472348 77120 472400 77172
rect 494060 76576 494112 76628
rect 495992 76576 496044 76628
rect 155960 75964 156012 76016
rect 156144 75964 156196 76016
rect 161020 75896 161072 75948
rect 161204 75896 161256 75948
rect 179328 75939 179380 75948
rect 179328 75905 179337 75939
rect 179337 75905 179371 75939
rect 179371 75905 179380 75939
rect 179328 75896 179380 75905
rect 186228 75939 186280 75948
rect 186228 75905 186237 75939
rect 186237 75905 186271 75939
rect 186271 75905 186280 75939
rect 186228 75896 186280 75905
rect 220728 75896 220780 75948
rect 223580 75939 223632 75948
rect 223580 75905 223589 75939
rect 223589 75905 223623 75939
rect 223623 75905 223632 75939
rect 223580 75896 223632 75905
rect 378140 75939 378192 75948
rect 378140 75905 378149 75939
rect 378149 75905 378183 75939
rect 378183 75905 378192 75939
rect 378140 75896 378192 75905
rect 511540 75939 511592 75948
rect 511540 75905 511549 75939
rect 511549 75905 511583 75939
rect 511583 75905 511592 75939
rect 511540 75896 511592 75905
rect 524420 75939 524472 75948
rect 524420 75905 524429 75939
rect 524429 75905 524463 75939
rect 524463 75905 524472 75939
rect 524420 75896 524472 75905
rect 532700 75939 532752 75948
rect 532700 75905 532709 75939
rect 532709 75905 532743 75939
rect 532743 75905 532752 75939
rect 532700 75896 532752 75905
rect 110420 75871 110472 75880
rect 110420 75837 110429 75871
rect 110429 75837 110463 75871
rect 110463 75837 110472 75871
rect 110420 75828 110472 75837
rect 494704 74468 494756 74520
rect 497556 74536 497608 74588
rect 80152 73176 80204 73228
rect 492772 73176 492824 73228
rect 494060 73176 494112 73228
rect 496728 73108 496780 73160
rect 503628 73176 503680 73228
rect 499948 73108 500000 73160
rect 500040 73108 500092 73160
rect 500684 73108 500736 73160
rect 500776 73108 500828 73160
rect 482560 71748 482612 71800
rect 485044 71748 485096 71800
rect 155960 70388 156012 70440
rect 156144 70252 156196 70304
rect 79692 69776 79744 69828
rect 79968 69776 80020 69828
rect 467104 68892 467156 68944
rect 470692 69028 470744 69080
rect 491024 68960 491076 69012
rect 492772 69028 492824 69080
rect 244280 67643 244332 67652
rect 244280 67609 244289 67643
rect 244289 67609 244323 67643
rect 244323 67609 244332 67643
rect 244280 67600 244332 67609
rect 258080 67643 258132 67652
rect 258080 67609 258089 67643
rect 258089 67609 258123 67643
rect 258123 67609 258132 67643
rect 258080 67600 258132 67609
rect 445852 67643 445904 67652
rect 445852 67609 445861 67643
rect 445861 67609 445895 67643
rect 445895 67609 445904 67643
rect 445852 67600 445904 67609
rect 436100 67575 436152 67584
rect 436100 67541 436109 67575
rect 436109 67541 436143 67575
rect 436143 67541 436152 67575
rect 436100 67532 436152 67541
rect 494244 66920 494296 66972
rect 496728 66920 496780 66972
rect 80060 66240 80112 66292
rect 80152 66240 80204 66292
rect 110420 66283 110472 66292
rect 110420 66249 110429 66283
rect 110429 66249 110463 66283
rect 110463 66249 110472 66283
rect 110420 66240 110472 66249
rect 152832 66172 152884 66224
rect 152924 66172 152976 66224
rect 156144 66172 156196 66224
rect 179328 66215 179380 66224
rect 179328 66181 179337 66215
rect 179337 66181 179371 66215
rect 179371 66181 179380 66215
rect 179328 66172 179380 66181
rect 186228 66215 186280 66224
rect 186228 66181 186237 66215
rect 186237 66181 186271 66215
rect 186271 66181 186280 66215
rect 186228 66172 186280 66181
rect 220728 66215 220780 66224
rect 220728 66181 220737 66215
rect 220737 66181 220771 66215
rect 220771 66181 220780 66215
rect 220728 66172 220780 66181
rect 223580 66215 223632 66224
rect 223580 66181 223589 66215
rect 223589 66181 223623 66215
rect 223623 66181 223632 66215
rect 223580 66172 223632 66181
rect 378140 66215 378192 66224
rect 378140 66181 378149 66215
rect 378149 66181 378183 66215
rect 378183 66181 378192 66215
rect 378140 66172 378192 66181
rect 511540 66215 511592 66224
rect 511540 66181 511549 66215
rect 511549 66181 511583 66215
rect 511583 66181 511592 66215
rect 511540 66172 511592 66181
rect 524420 66215 524472 66224
rect 524420 66181 524429 66215
rect 524429 66181 524463 66215
rect 524463 66181 524472 66215
rect 524420 66172 524472 66181
rect 532700 66215 532752 66224
rect 532700 66181 532709 66215
rect 532709 66181 532743 66215
rect 532743 66181 532752 66215
rect 532700 66172 532752 66181
rect 161020 64855 161072 64864
rect 161020 64821 161029 64855
rect 161029 64821 161063 64855
rect 161063 64821 161072 64855
rect 161020 64812 161072 64821
rect 478880 64812 478932 64864
rect 482560 64880 482612 64932
rect 487160 64880 487212 64932
rect 491024 64880 491076 64932
rect 519544 64812 519596 64864
rect 580172 64812 580224 64864
rect 2780 64540 2832 64592
rect 4896 64540 4948 64592
rect 505836 63520 505888 63572
rect 505928 63520 505980 63572
rect 117320 62092 117372 62144
rect 117596 62092 117648 62144
rect 120080 62092 120132 62144
rect 120356 62092 120408 62144
rect 476028 62024 476080 62076
rect 478880 62092 478932 62144
rect 482284 62092 482336 62144
rect 487160 62092 487212 62144
rect 491944 62092 491996 62144
rect 494244 62092 494296 62144
rect 117596 60800 117648 60852
rect 120356 60800 120408 60852
rect 505836 60732 505888 60784
rect 117504 60664 117556 60716
rect 120264 60664 120316 60716
rect 505928 60596 505980 60648
rect 436100 57987 436152 57996
rect 436100 57953 436109 57987
rect 436109 57953 436143 57987
rect 436143 57953 436152 57987
rect 436100 57944 436152 57953
rect 244280 57919 244332 57928
rect 244280 57885 244289 57919
rect 244289 57885 244323 57919
rect 244323 57885 244332 57919
rect 244280 57876 244332 57885
rect 258080 57919 258132 57928
rect 258080 57885 258089 57919
rect 258089 57885 258123 57919
rect 258123 57885 258132 57919
rect 258080 57876 258132 57885
rect 289544 57876 289596 57928
rect 289728 57876 289780 57928
rect 445852 57919 445904 57928
rect 445852 57885 445861 57919
rect 445861 57885 445895 57919
rect 445895 57885 445904 57919
rect 445852 57876 445904 57885
rect 471980 57876 472032 57928
rect 476028 57944 476080 57996
rect 436100 57851 436152 57860
rect 436100 57817 436109 57851
rect 436109 57817 436143 57851
rect 436143 57817 436152 57851
rect 436100 57808 436152 57817
rect 465724 57604 465776 57656
rect 467104 57604 467156 57656
rect 493600 57468 493652 57520
rect 494704 57468 494756 57520
rect 110420 56720 110472 56772
rect 79600 56584 79652 56636
rect 79692 56584 79744 56636
rect 110420 56584 110472 56636
rect 155960 56627 156012 56636
rect 155960 56593 155969 56627
rect 155969 56593 156003 56627
rect 156003 56593 156012 56627
rect 155960 56584 156012 56593
rect 179328 56627 179380 56636
rect 179328 56593 179337 56627
rect 179337 56593 179371 56627
rect 179371 56593 179380 56627
rect 179328 56584 179380 56593
rect 186228 56627 186280 56636
rect 186228 56593 186237 56627
rect 186237 56593 186271 56627
rect 186271 56593 186280 56627
rect 186228 56584 186280 56593
rect 220728 56627 220780 56636
rect 220728 56593 220737 56627
rect 220737 56593 220771 56627
rect 220771 56593 220780 56627
rect 220728 56584 220780 56593
rect 223580 56627 223632 56636
rect 223580 56593 223589 56627
rect 223589 56593 223623 56627
rect 223623 56593 223632 56627
rect 223580 56584 223632 56593
rect 378140 56627 378192 56636
rect 378140 56593 378149 56627
rect 378149 56593 378183 56627
rect 378183 56593 378192 56627
rect 378140 56584 378192 56593
rect 511540 56627 511592 56636
rect 511540 56593 511549 56627
rect 511549 56593 511583 56627
rect 511583 56593 511592 56627
rect 511540 56584 511592 56593
rect 524420 56627 524472 56636
rect 524420 56593 524429 56627
rect 524429 56593 524463 56627
rect 524463 56593 524472 56627
rect 524420 56584 524472 56593
rect 532700 56627 532752 56636
rect 532700 56593 532709 56627
rect 532709 56593 532743 56627
rect 532743 56593 532752 56627
rect 532700 56584 532752 56593
rect 110420 56491 110472 56500
rect 110420 56457 110429 56491
rect 110429 56457 110463 56491
rect 110463 56457 110472 56491
rect 110420 56448 110472 56457
rect 161388 55224 161440 55276
rect 289544 53864 289596 53916
rect 289728 53864 289780 53916
rect 490288 53864 490340 53916
rect 491944 53864 491996 53916
rect 467104 53660 467156 53712
rect 471980 53796 472032 53848
rect 481272 53796 481324 53848
rect 482284 53796 482336 53848
rect 488540 53728 488592 53780
rect 490288 53728 490340 53780
rect 79600 53388 79652 53440
rect 79968 53388 80020 53440
rect 220544 51076 220596 51128
rect 3424 51008 3476 51060
rect 15844 51008 15896 51060
rect 220360 51008 220412 51060
rect 272892 51008 272944 51060
rect 273076 51008 273128 51060
rect 299204 51008 299256 51060
rect 299388 51008 299440 51060
rect 351644 51008 351696 51060
rect 351828 51008 351880 51060
rect 155960 50872 156012 50924
rect 156144 50872 156196 50924
rect 491484 49784 491536 49836
rect 493600 49784 493652 49836
rect 289636 48424 289688 48476
rect 161112 48288 161164 48340
rect 161388 48288 161440 48340
rect 244280 48331 244332 48340
rect 244280 48297 244289 48331
rect 244289 48297 244323 48331
rect 244323 48297 244332 48331
rect 244280 48288 244332 48297
rect 258080 48331 258132 48340
rect 258080 48297 258089 48331
rect 258089 48297 258123 48331
rect 258123 48297 258132 48331
rect 258080 48288 258132 48297
rect 436100 48331 436152 48340
rect 436100 48297 436109 48331
rect 436109 48297 436143 48331
rect 436143 48297 436152 48331
rect 436100 48288 436152 48297
rect 445852 48331 445904 48340
rect 445852 48297 445861 48331
rect 445861 48297 445895 48331
rect 445895 48297 445904 48331
rect 445852 48288 445904 48297
rect 273076 48220 273128 48272
rect 289636 48220 289688 48272
rect 299388 48263 299440 48272
rect 299388 48229 299397 48263
rect 299397 48229 299431 48263
rect 299431 48229 299440 48263
rect 299388 48220 299440 48229
rect 351828 48220 351880 48272
rect 487896 47336 487948 47388
rect 488540 47336 488592 47388
rect 488540 46996 488592 47048
rect 491484 46996 491536 47048
rect 110420 46971 110472 46980
rect 110420 46937 110429 46971
rect 110429 46937 110463 46971
rect 110463 46937 110472 46971
rect 110420 46928 110472 46937
rect 479616 46928 479668 46980
rect 481272 46928 481324 46980
rect 156144 46860 156196 46912
rect 161112 46903 161164 46912
rect 161112 46869 161121 46903
rect 161121 46869 161155 46903
rect 161155 46869 161164 46903
rect 161112 46860 161164 46869
rect 179328 46860 179380 46912
rect 186228 46903 186280 46912
rect 186228 46869 186237 46903
rect 186237 46869 186271 46903
rect 186271 46869 186280 46903
rect 186228 46860 186280 46869
rect 220728 46860 220780 46912
rect 223580 46903 223632 46912
rect 223580 46869 223589 46903
rect 223589 46869 223623 46903
rect 223623 46869 223632 46903
rect 223580 46860 223632 46869
rect 289728 46903 289780 46912
rect 289728 46869 289737 46903
rect 289737 46869 289771 46903
rect 289771 46869 289780 46903
rect 289728 46860 289780 46869
rect 378140 46903 378192 46912
rect 378140 46869 378149 46903
rect 378149 46869 378183 46903
rect 378183 46869 378192 46903
rect 378140 46860 378192 46869
rect 505928 46860 505980 46912
rect 511540 46903 511592 46912
rect 511540 46869 511549 46903
rect 511549 46869 511583 46903
rect 511583 46869 511592 46903
rect 511540 46860 511592 46869
rect 524420 46903 524472 46912
rect 524420 46869 524429 46903
rect 524429 46869 524463 46903
rect 524463 46869 524472 46903
rect 524420 46860 524472 46869
rect 532700 46903 532752 46912
rect 532700 46869 532709 46903
rect 532709 46869 532743 46903
rect 532743 46869 532752 46903
rect 532700 46860 532752 46869
rect 82636 45611 82688 45620
rect 82636 45577 82645 45611
rect 82645 45577 82679 45611
rect 82679 45577 82688 45611
rect 82636 45568 82688 45577
rect 121552 45568 121604 45620
rect 121644 45568 121696 45620
rect 79968 44820 80020 44872
rect 335360 44820 335412 44872
rect 82636 44183 82688 44192
rect 82636 44149 82645 44183
rect 82645 44149 82679 44183
rect 82679 44149 82688 44183
rect 82636 44140 82688 44149
rect 83372 44140 83424 44192
rect 83464 44140 83516 44192
rect 500684 44140 500736 44192
rect 500776 44140 500828 44192
rect 156052 41395 156104 41404
rect 156052 41361 156061 41395
rect 156061 41361 156095 41395
rect 156095 41361 156104 41395
rect 156052 41352 156104 41361
rect 540244 41352 540296 41404
rect 580172 41352 580224 41404
rect 505928 41216 505980 41268
rect 486148 40128 486200 40180
rect 487896 40128 487948 40180
rect 487804 39992 487856 40044
rect 488540 39992 488592 40044
rect 117688 39312 117740 39364
rect 120448 39312 120500 39364
rect 459560 39312 459612 39364
rect 465724 39312 465776 39364
rect 272984 38675 273036 38684
rect 272984 38641 272993 38675
rect 272993 38641 273027 38675
rect 273027 38641 273036 38675
rect 272984 38632 273036 38641
rect 299296 38632 299348 38684
rect 351736 38675 351788 38684
rect 351736 38641 351745 38675
rect 351745 38641 351779 38675
rect 351779 38641 351788 38675
rect 351736 38632 351788 38641
rect 244280 38607 244332 38616
rect 244280 38573 244289 38607
rect 244289 38573 244323 38607
rect 244323 38573 244332 38607
rect 244280 38564 244332 38573
rect 258080 38607 258132 38616
rect 258080 38573 258089 38607
rect 258089 38573 258123 38607
rect 258123 38573 258132 38607
rect 258080 38564 258132 38573
rect 436100 38607 436152 38616
rect 436100 38573 436109 38607
rect 436109 38573 436143 38607
rect 436143 38573 436152 38607
rect 436100 38564 436152 38573
rect 445852 38607 445904 38616
rect 445852 38573 445861 38607
rect 445861 38573 445895 38607
rect 445895 38573 445904 38607
rect 445852 38564 445904 38573
rect 476856 38564 476908 38616
rect 479616 38564 479668 38616
rect 505836 38564 505888 38616
rect 505928 38564 505980 38616
rect 88248 37884 88300 37936
rect 505560 37884 505612 37936
rect 110420 37408 110472 37460
rect 110420 37272 110472 37324
rect 161204 37272 161256 37324
rect 179236 37315 179288 37324
rect 179236 37281 179245 37315
rect 179245 37281 179279 37315
rect 179279 37281 179288 37315
rect 179236 37272 179288 37281
rect 186228 37315 186280 37324
rect 186228 37281 186237 37315
rect 186237 37281 186271 37315
rect 186271 37281 186280 37315
rect 186228 37272 186280 37281
rect 220728 37272 220780 37324
rect 223580 37315 223632 37324
rect 223580 37281 223589 37315
rect 223589 37281 223623 37315
rect 223623 37281 223632 37315
rect 223580 37272 223632 37281
rect 289728 37315 289780 37324
rect 289728 37281 289737 37315
rect 289737 37281 289771 37315
rect 289771 37281 289780 37315
rect 289728 37272 289780 37281
rect 361488 37272 361540 37324
rect 362960 37272 363012 37324
rect 378140 37315 378192 37324
rect 378140 37281 378149 37315
rect 378149 37281 378183 37315
rect 378183 37281 378192 37315
rect 378140 37272 378192 37281
rect 524420 37315 524472 37324
rect 524420 37281 524429 37315
rect 524429 37281 524463 37315
rect 524463 37281 524472 37315
rect 524420 37272 524472 37281
rect 532700 37315 532752 37324
rect 532700 37281 532709 37315
rect 532709 37281 532743 37315
rect 532743 37281 532752 37315
rect 532700 37272 532752 37281
rect 220452 37247 220504 37256
rect 220452 37213 220461 37247
rect 220461 37213 220495 37247
rect 220495 37213 220504 37247
rect 220452 37204 220504 37213
rect 110420 37179 110472 37188
rect 110420 37145 110429 37179
rect 110429 37145 110463 37179
rect 110463 37145 110472 37179
rect 110420 37136 110472 37145
rect 484216 36864 484268 36916
rect 486148 36864 486200 36916
rect 457444 36320 457496 36372
rect 459560 36320 459612 36372
rect 3148 35844 3200 35896
rect 6184 35844 6236 35896
rect 83740 35844 83792 35896
rect 83832 35844 83884 35896
rect 161204 32487 161256 32496
rect 161204 32453 161213 32487
rect 161213 32453 161247 32487
rect 161247 32453 161256 32487
rect 161204 32444 161256 32453
rect 351736 31832 351788 31884
rect 153108 31764 153160 31816
rect 156052 31696 156104 31748
rect 156236 31696 156288 31748
rect 351736 31696 351788 31748
rect 505836 29656 505888 29708
rect 436100 29087 436152 29096
rect 436100 29053 436109 29087
rect 436109 29053 436143 29087
rect 436143 29053 436152 29087
rect 436100 29044 436152 29053
rect 511540 29087 511592 29096
rect 511540 29053 511549 29087
rect 511549 29053 511583 29087
rect 511583 29053 511592 29087
rect 511540 29044 511592 29053
rect 152924 29019 152976 29028
rect 152924 28985 152933 29019
rect 152933 28985 152967 29019
rect 152967 28985 152976 29019
rect 152924 28976 152976 28985
rect 244280 29019 244332 29028
rect 244280 28985 244289 29019
rect 244289 28985 244323 29019
rect 244323 28985 244332 29019
rect 244280 28976 244332 28985
rect 258080 29019 258132 29028
rect 258080 28985 258089 29019
rect 258089 28985 258123 29019
rect 258123 28985 258132 29019
rect 258080 28976 258132 28985
rect 425612 28976 425664 29028
rect 427820 28976 427872 29028
rect 445852 29019 445904 29028
rect 445852 28985 445861 29019
rect 445861 28985 445895 29019
rect 445895 28985 445904 29019
rect 445852 28976 445904 28985
rect 156236 28908 156288 28960
rect 161480 28951 161532 28960
rect 161480 28917 161489 28951
rect 161489 28917 161523 28951
rect 161523 28917 161532 28951
rect 161480 28908 161532 28917
rect 436100 28908 436152 28960
rect 436192 28908 436244 28960
rect 480260 28908 480312 28960
rect 484216 28976 484268 29028
rect 110420 27659 110472 27668
rect 110420 27625 110429 27659
rect 110429 27625 110463 27659
rect 110463 27625 110472 27659
rect 110420 27616 110472 27625
rect 117596 27616 117648 27668
rect 120356 27616 120408 27668
rect 161204 27659 161256 27668
rect 161204 27625 161213 27659
rect 161213 27625 161247 27659
rect 161247 27625 161256 27659
rect 161204 27616 161256 27625
rect 220544 27616 220596 27668
rect 152924 27591 152976 27600
rect 152924 27557 152933 27591
rect 152933 27557 152967 27591
rect 152967 27557 152976 27591
rect 152924 27548 152976 27557
rect 179328 27548 179380 27600
rect 186228 27548 186280 27600
rect 220728 27591 220780 27600
rect 220728 27557 220737 27591
rect 220737 27557 220771 27591
rect 220771 27557 220780 27591
rect 220728 27548 220780 27557
rect 223580 27591 223632 27600
rect 223580 27557 223589 27591
rect 223589 27557 223623 27591
rect 223623 27557 223632 27591
rect 223580 27548 223632 27557
rect 289728 27591 289780 27600
rect 289728 27557 289737 27591
rect 289737 27557 289771 27591
rect 289771 27557 289780 27591
rect 289728 27548 289780 27557
rect 299112 27591 299164 27600
rect 299112 27557 299121 27591
rect 299121 27557 299155 27591
rect 299155 27557 299164 27591
rect 299112 27548 299164 27557
rect 362960 27548 363012 27600
rect 363236 27548 363288 27600
rect 378140 27591 378192 27600
rect 378140 27557 378149 27591
rect 378149 27557 378183 27591
rect 378183 27557 378192 27591
rect 378140 27548 378192 27557
rect 454684 27548 454736 27600
rect 457444 27548 457496 27600
rect 511540 27591 511592 27600
rect 511540 27557 511549 27591
rect 511549 27557 511583 27591
rect 511583 27557 511592 27591
rect 511540 27548 511592 27557
rect 524420 27591 524472 27600
rect 524420 27557 524429 27591
rect 524429 27557 524463 27591
rect 524463 27557 524472 27591
rect 524420 27548 524472 27557
rect 532700 27591 532752 27600
rect 532700 27557 532709 27591
rect 532709 27557 532743 27591
rect 532743 27557 532752 27591
rect 532700 27548 532752 27557
rect 478880 24828 478932 24880
rect 480260 24828 480312 24880
rect 117504 22108 117556 22160
rect 272892 22040 272944 22092
rect 273076 22040 273128 22092
rect 161112 20544 161164 20596
rect 161296 20544 161348 20596
rect 156144 19363 156196 19372
rect 156144 19329 156153 19363
rect 156153 19329 156187 19363
rect 156187 19329 156196 19363
rect 156144 19320 156196 19329
rect 131212 19295 131264 19304
rect 131212 19261 131221 19295
rect 131221 19261 131255 19295
rect 131255 19261 131264 19295
rect 131212 19252 131264 19261
rect 244280 19295 244332 19304
rect 244280 19261 244289 19295
rect 244289 19261 244323 19295
rect 244323 19261 244332 19295
rect 244280 19252 244332 19261
rect 258080 19252 258132 19304
rect 258264 19252 258316 19304
rect 351828 19252 351880 19304
rect 427636 19252 427688 19304
rect 427820 19252 427872 19304
rect 436100 19295 436152 19304
rect 436100 19261 436109 19295
rect 436109 19261 436143 19295
rect 436143 19261 436152 19295
rect 436100 19252 436152 19261
rect 445852 19295 445904 19304
rect 445852 19261 445861 19295
rect 445861 19261 445895 19295
rect 445895 19261 445904 19295
rect 445852 19252 445904 19261
rect 474832 19252 474884 19304
rect 478880 19388 478932 19440
rect 463700 19184 463752 19236
rect 467104 19184 467156 19236
rect 505744 19227 505796 19236
rect 505744 19193 505753 19227
rect 505753 19193 505787 19227
rect 505787 19193 505796 19227
rect 505744 19184 505796 19193
rect 475016 18300 475068 18352
rect 476856 18300 476908 18352
rect 110420 18096 110472 18148
rect 110420 17960 110472 18012
rect 153016 17960 153068 18012
rect 161572 17960 161624 18012
rect 220728 18003 220780 18012
rect 220728 17969 220737 18003
rect 220737 17969 220771 18003
rect 220771 17969 220780 18003
rect 220728 17960 220780 17969
rect 223580 18003 223632 18012
rect 223580 17969 223589 18003
rect 223589 17969 223623 18003
rect 223623 17969 223632 18003
rect 223580 17960 223632 17969
rect 299204 17960 299256 18012
rect 378140 18003 378192 18012
rect 378140 17969 378149 18003
rect 378149 17969 378183 18003
rect 378183 17969 378192 18003
rect 378140 17960 378192 17969
rect 511540 18003 511592 18012
rect 511540 17969 511549 18003
rect 511549 17969 511583 18003
rect 511583 17969 511592 18003
rect 511540 17960 511592 17969
rect 524420 18003 524472 18012
rect 524420 17969 524429 18003
rect 524429 17969 524463 18003
rect 524463 17969 524472 18003
rect 524420 17960 524472 17969
rect 340788 17484 340840 17536
rect 505192 17484 505244 17536
rect 119528 17416 119580 17468
rect 504180 17416 504232 17468
rect 99196 17348 99248 17400
rect 504824 17348 504876 17400
rect 96528 17280 96580 17332
rect 503904 17280 503956 17332
rect 56416 17212 56468 17264
rect 506020 17212 506072 17264
rect 452660 17144 452712 17196
rect 454684 17144 454736 17196
rect 471336 16600 471388 16652
rect 474832 16600 474884 16652
rect 259368 15988 259420 16040
rect 401600 15988 401652 16040
rect 293868 15920 293920 15972
rect 505468 15920 505520 15972
rect 158628 15852 158680 15904
rect 504088 15852 504140 15904
rect 117412 15215 117464 15224
rect 117412 15181 117421 15215
rect 117421 15181 117455 15215
rect 117455 15181 117464 15215
rect 117412 15172 117464 15181
rect 120080 15172 120132 15224
rect 120172 15172 120224 15224
rect 461860 15172 461912 15224
rect 463700 15172 463752 15224
rect 295248 14832 295300 14884
rect 302240 14832 302292 14884
rect 256608 14764 256660 14816
rect 313280 14764 313332 14816
rect 272892 14696 272944 14748
rect 333980 14696 334032 14748
rect 474740 14696 474792 14748
rect 226248 14628 226300 14680
rect 365720 14628 365772 14680
rect 156144 14603 156196 14612
rect 156144 14569 156153 14603
rect 156153 14569 156187 14603
rect 156187 14569 156196 14603
rect 156144 14560 156196 14569
rect 200028 14560 200080 14612
rect 351920 14560 351972 14612
rect 81256 14492 81308 14544
rect 367100 14492 367152 14544
rect 375196 14492 375248 14544
rect 405740 14492 405792 14544
rect 79416 14424 79468 14476
rect 412640 14424 412692 14476
rect 332508 13608 332560 13660
rect 501972 13608 502024 13660
rect 335268 13540 335320 13592
rect 193128 13472 193180 13524
rect 386420 13472 386472 13524
rect 498200 13404 498252 13456
rect 78680 13336 78732 13388
rect 358820 13336 358872 13388
rect 371148 13336 371200 13388
rect 184848 13268 184900 13320
rect 470600 13268 470652 13320
rect 220452 13200 220504 13252
rect 284300 13200 284352 13252
rect 289636 13200 289688 13252
rect 576860 13200 576912 13252
rect 79876 13132 79928 13184
rect 377680 13132 377732 13184
rect 109960 13064 110012 13116
rect 110328 13064 110380 13116
rect 219348 13064 219400 13116
rect 565820 13064 565872 13116
rect 220728 12520 220780 12572
rect 393228 12520 393280 12572
rect 119528 12452 119580 12504
rect 135076 12452 135128 12504
rect 153016 12452 153068 12504
rect 222108 12452 222160 12504
rect 289728 12495 289780 12504
rect 289728 12461 289737 12495
rect 289737 12461 289771 12495
rect 289771 12461 289780 12495
rect 289728 12452 289780 12461
rect 369952 12452 370004 12504
rect 371240 12452 371292 12504
rect 372620 12452 372672 12504
rect 378140 12452 378192 12504
rect 99012 12384 99064 12436
rect 99196 12384 99248 12436
rect 106464 12384 106516 12436
rect 107384 12384 107436 12436
rect 119436 12384 119488 12436
rect 128360 12384 128412 12436
rect 129004 12384 129056 12436
rect 134892 12384 134944 12436
rect 152740 12384 152792 12436
rect 196072 12384 196124 12436
rect 196808 12384 196860 12436
rect 349160 12384 349212 12436
rect 350264 12384 350316 12436
rect 351920 12384 351972 12436
rect 352472 12384 352524 12436
rect 360200 12384 360252 12436
rect 360936 12384 360988 12436
rect 367100 12384 367152 12436
rect 368020 12384 368072 12436
rect 370412 12316 370464 12368
rect 371608 12316 371660 12368
rect 372804 12316 372856 12368
rect 426440 12384 426492 12436
rect 427544 12384 427596 12436
rect 458272 12384 458324 12436
rect 461860 12452 461912 12504
rect 482836 12452 482888 12504
rect 487804 12452 487856 12504
rect 511540 12452 511592 12504
rect 524420 12452 524472 12504
rect 511448 12384 511500 12436
rect 523040 12384 523092 12436
rect 523868 12384 523920 12436
rect 378784 12316 378836 12368
rect 529940 12384 529992 12436
rect 531044 12384 531096 12436
rect 534080 12384 534132 12436
rect 534540 12384 534592 12436
rect 538220 12384 538272 12436
rect 539324 12384 539376 12436
rect 542360 12384 542412 12436
rect 542912 12384 542964 12436
rect 525064 12316 525116 12368
rect 527456 12359 527508 12368
rect 527456 12325 527465 12359
rect 527465 12325 527499 12359
rect 527499 12325 527508 12359
rect 527456 12316 527508 12325
rect 181352 12112 181404 12164
rect 245660 12112 245712 12164
rect 138480 12044 138532 12096
rect 251180 12044 251232 12096
rect 325608 12044 325660 12096
rect 429936 12044 429988 12096
rect 154488 11976 154540 12028
rect 230480 11976 230532 12028
rect 249616 11976 249668 12028
rect 462044 11976 462096 12028
rect 216496 11908 216548 11960
rect 506020 11908 506072 11960
rect 76564 11840 76616 11892
rect 76840 11840 76892 11892
rect 155132 11840 155184 11892
rect 477500 11840 477552 11892
rect 104808 11772 104860 11824
rect 495348 11772 495400 11824
rect 84016 11704 84068 11756
rect 509608 11704 509660 11756
rect 245476 11543 245528 11552
rect 245476 11509 245485 11543
rect 245485 11509 245519 11543
rect 245519 11509 245528 11543
rect 245476 11500 245528 11509
rect 471612 10956 471664 11008
rect 475016 11024 475068 11076
rect 445760 10888 445812 10940
rect 452660 10888 452712 10940
rect 84108 10548 84160 10600
rect 309140 10548 309192 10600
rect 354588 10548 354640 10600
rect 546592 10548 546644 10600
rect 115848 10480 115900 10532
rect 137284 10480 137336 10532
rect 173808 10480 173860 10532
rect 191840 10480 191892 10532
rect 194416 10480 194468 10532
rect 467840 10480 467892 10532
rect 79784 10412 79836 10464
rect 383568 10412 383620 10464
rect 491208 10412 491260 10464
rect 571432 10412 571484 10464
rect 79508 10344 79560 10396
rect 404912 10344 404964 10396
rect 438768 10344 438820 10396
rect 581092 10344 581144 10396
rect 135168 10276 135220 10328
rect 491392 10276 491444 10328
rect 186044 9775 186096 9784
rect 186044 9741 186053 9775
rect 186053 9741 186087 9775
rect 186087 9741 186096 9775
rect 186044 9732 186096 9741
rect 351736 9775 351788 9784
rect 351736 9741 351745 9775
rect 351745 9741 351779 9775
rect 351779 9741 351788 9775
rect 351736 9732 351788 9741
rect 436100 9775 436152 9784
rect 436100 9741 436109 9775
rect 436109 9741 436143 9775
rect 436143 9741 436152 9775
rect 436100 9732 436152 9741
rect 131212 9707 131264 9716
rect 131212 9673 131221 9707
rect 131221 9673 131255 9707
rect 131255 9673 131264 9707
rect 131212 9664 131264 9673
rect 156236 9664 156288 9716
rect 161480 9664 161532 9716
rect 161572 9664 161624 9716
rect 178960 9707 179012 9716
rect 178960 9673 178969 9707
rect 178969 9673 179003 9707
rect 179003 9673 179012 9707
rect 178960 9664 179012 9673
rect 220544 9707 220596 9716
rect 220544 9673 220553 9707
rect 220553 9673 220587 9707
rect 220587 9673 220596 9707
rect 220544 9664 220596 9673
rect 221740 9707 221792 9716
rect 221740 9673 221749 9707
rect 221749 9673 221783 9707
rect 221783 9673 221792 9707
rect 221740 9664 221792 9673
rect 244280 9707 244332 9716
rect 244280 9673 244289 9707
rect 244289 9673 244323 9707
rect 244323 9673 244332 9707
rect 244280 9664 244332 9673
rect 341892 9707 341944 9716
rect 341892 9673 341901 9707
rect 341901 9673 341935 9707
rect 341935 9673 341944 9707
rect 341892 9664 341944 9673
rect 393044 9707 393096 9716
rect 393044 9673 393053 9707
rect 393053 9673 393087 9707
rect 393087 9673 393096 9707
rect 393044 9664 393096 9673
rect 445852 9707 445904 9716
rect 445852 9673 445861 9707
rect 445861 9673 445895 9707
rect 445895 9673 445904 9707
rect 445852 9664 445904 9673
rect 533436 9664 533488 9716
rect 541716 9707 541768 9716
rect 541716 9673 541725 9707
rect 541725 9673 541759 9707
rect 541759 9673 541768 9707
rect 541716 9664 541768 9673
rect 99472 9596 99524 9648
rect 134892 9639 134944 9648
rect 134892 9605 134901 9639
rect 134901 9605 134935 9639
rect 134935 9605 134944 9639
rect 134892 9596 134944 9605
rect 186044 9639 186096 9648
rect 186044 9605 186053 9639
rect 186053 9605 186087 9639
rect 186087 9605 186096 9639
rect 186044 9596 186096 9605
rect 195612 9596 195664 9648
rect 245476 9596 245528 9648
rect 245660 9596 245712 9648
rect 258080 9596 258132 9648
rect 351736 9639 351788 9648
rect 351736 9605 351745 9639
rect 351745 9605 351779 9639
rect 351779 9605 351788 9639
rect 351736 9596 351788 9605
rect 370412 9639 370464 9648
rect 370412 9605 370421 9639
rect 370421 9605 370455 9639
rect 370455 9605 370464 9639
rect 370412 9596 370464 9605
rect 371608 9639 371660 9648
rect 371608 9605 371617 9639
rect 371617 9605 371651 9639
rect 371651 9605 371660 9639
rect 371608 9596 371660 9605
rect 372804 9639 372856 9648
rect 372804 9605 372813 9639
rect 372813 9605 372847 9639
rect 372847 9605 372856 9639
rect 372804 9596 372856 9605
rect 377588 9639 377640 9648
rect 377588 9605 377597 9639
rect 377597 9605 377631 9639
rect 377631 9605 377640 9639
rect 377588 9596 377640 9605
rect 378784 9639 378836 9648
rect 378784 9605 378793 9639
rect 378793 9605 378827 9639
rect 378827 9605 378836 9639
rect 378784 9596 378836 9605
rect 427820 9596 427872 9648
rect 436100 9596 436152 9648
rect 525064 9596 525116 9648
rect 527456 9596 527508 9648
rect 195612 9460 195664 9512
rect 525064 9460 525116 9512
rect 527456 9460 527508 9512
rect 83832 9392 83884 9444
rect 171784 9392 171836 9444
rect 81716 9324 81768 9376
rect 222936 9324 222988 9376
rect 126612 9256 126664 9308
rect 287152 9256 287204 9308
rect 83464 9188 83516 9240
rect 308588 9188 308640 9240
rect 413928 9188 413980 9240
rect 501236 9188 501288 9240
rect 81440 9120 81492 9172
rect 358544 9120 358596 9172
rect 436008 9120 436060 9172
rect 526260 9120 526312 9172
rect 150348 9052 150400 9104
rect 540520 9052 540572 9104
rect 89536 8984 89588 9036
rect 519084 8984 519136 9036
rect 108948 8916 109000 8968
rect 551192 8916 551244 8968
rect 3424 8236 3476 8288
rect 508688 8236 508740 8288
rect 117136 8168 117188 8220
rect 253940 8168 253992 8220
rect 262128 8168 262180 8220
rect 400220 8168 400272 8220
rect 113548 8100 113600 8152
rect 327080 8100 327132 8152
rect 171048 8032 171100 8084
rect 457260 8032 457312 8084
rect 102784 7964 102836 8016
rect 408500 7964 408552 8016
rect 33876 7896 33928 7948
rect 340880 7896 340932 7948
rect 18328 7828 18380 7880
rect 329840 7828 329892 7880
rect 124220 7760 124272 7812
rect 438860 7760 438912 7812
rect 21916 7692 21968 7744
rect 346400 7692 346452 7744
rect 357348 7692 357400 7744
rect 402980 7692 403032 7744
rect 44548 7624 44600 7676
rect 396172 7624 396224 7676
rect 401600 7624 401652 7676
rect 402520 7624 402572 7676
rect 419540 7624 419592 7676
rect 420368 7624 420420 7676
rect 433340 7624 433392 7676
rect 434628 7624 434680 7676
rect 459468 7624 459520 7676
rect 529848 7624 529900 7676
rect 50528 7556 50580 7608
rect 484400 7556 484452 7608
rect 520280 7556 520332 7608
rect 521476 7556 521528 7608
rect 536840 7556 536892 7608
rect 538128 7556 538180 7608
rect 81532 7488 81584 7540
rect 183744 7488 183796 7540
rect 287060 7488 287112 7540
rect 288348 7488 288400 7540
rect 365720 7488 365772 7540
rect 366916 7488 366968 7540
rect 478052 7352 478104 7404
rect 482836 7352 482888 7404
rect 500040 7216 500092 7268
rect 500684 7216 500736 7268
rect 469312 7148 469364 7200
rect 471612 7148 471664 7200
rect 76564 6876 76616 6928
rect 76932 6876 76984 6928
rect 82636 6876 82688 6928
rect 120172 6876 120224 6928
rect 120264 6876 120316 6928
rect 82544 6672 82596 6724
rect 110420 6808 110472 6860
rect 117412 6808 117464 6860
rect 118240 6808 118292 6860
rect 395436 6808 395488 6860
rect 510896 6808 510948 6860
rect 382372 6740 382424 6792
rect 511080 6740 511132 6792
rect 376392 6672 376444 6724
rect 507768 6672 507820 6724
rect 77024 6604 77076 6656
rect 159916 6604 159968 6656
rect 345480 6604 345532 6656
rect 509516 6604 509568 6656
rect 78312 6536 78364 6588
rect 261024 6536 261076 6588
rect 346676 6536 346728 6588
rect 510988 6536 511040 6588
rect 78496 6468 78548 6520
rect 281264 6468 281316 6520
rect 299204 6468 299256 6520
rect 520280 6468 520332 6520
rect 99288 6400 99340 6452
rect 409696 6400 409748 6452
rect 410892 6400 410944 6452
rect 502432 6400 502484 6452
rect 78404 6332 78456 6384
rect 417976 6332 418028 6384
rect 423956 6332 424008 6384
rect 509424 6332 509476 6384
rect 74356 6264 74408 6316
rect 472716 6264 472768 6316
rect 497740 6264 497792 6316
rect 510804 6264 510856 6316
rect 77760 6196 77812 6248
rect 502432 6196 502484 6248
rect 74448 6128 74500 6180
rect 516784 6128 516836 6180
rect 432328 6060 432380 6112
rect 505744 6060 505796 6112
rect 451372 5992 451424 6044
rect 508320 5992 508372 6044
rect 471244 5652 471296 5704
rect 478052 5652 478104 5704
rect 469220 5516 469272 5568
rect 471336 5516 471388 5568
rect 499948 5516 500000 5568
rect 500132 5516 500184 5568
rect 256240 5448 256292 5500
rect 296720 5448 296772 5500
rect 297824 5448 297876 5500
rect 418160 5448 418212 5500
rect 442908 5448 442960 5500
rect 467932 5448 467984 5500
rect 213828 5380 213880 5432
rect 294328 5380 294380 5432
rect 300308 5380 300360 5432
rect 445760 5380 445812 5432
rect 245568 5312 245620 5364
rect 394240 5312 394292 5364
rect 415676 5312 415728 5364
rect 491300 5312 491352 5364
rect 176568 5244 176620 5296
rect 183560 5244 183612 5296
rect 201592 5244 201644 5296
rect 357440 5244 357492 5296
rect 373908 5244 373960 5296
rect 476304 5244 476356 5296
rect 127808 5176 127860 5228
rect 281540 5176 281592 5228
rect 291936 5176 291988 5228
rect 458272 5176 458324 5228
rect 107476 5108 107528 5160
rect 312176 5108 312228 5160
rect 337108 5108 337160 5160
rect 481640 5108 481692 5160
rect 114468 5040 114520 5092
rect 187240 5040 187292 5092
rect 262220 5040 262272 5092
rect 469220 5040 469272 5092
rect 118608 4972 118660 5024
rect 205088 4972 205140 5024
rect 212356 4972 212408 5024
rect 233700 4972 233752 5024
rect 251456 4972 251508 5024
rect 469312 4972 469364 5024
rect 84844 4904 84896 4956
rect 140872 4904 140924 4956
rect 144460 4904 144512 4956
rect 387800 4904 387852 4956
rect 471244 4904 471296 4956
rect 101956 4836 102008 4888
rect 426348 4836 426400 4888
rect 433248 4836 433300 4888
rect 475108 4836 475160 4888
rect 81900 4768 81952 4820
rect 522672 4768 522724 4820
rect 333612 4700 333664 4752
rect 444380 4700 444432 4752
rect 362132 4632 362184 4684
rect 385040 4632 385092 4684
rect 408500 4632 408552 4684
rect 455420 4632 455472 4684
rect 379980 4564 380032 4616
rect 419632 4564 419684 4616
rect 500132 4292 500184 4344
rect 494704 4224 494756 4276
rect 495624 4224 495676 4276
rect 572 4088 624 4140
rect 9036 4088 9088 4140
rect 32680 4088 32732 4140
rect 51724 4088 51776 4140
rect 76656 4088 76708 4140
rect 77116 4088 77168 4140
rect 84936 4088 84988 4140
rect 85488 4088 85540 4140
rect 87328 4088 87380 4140
rect 88248 4088 88300 4140
rect 95700 4088 95752 4140
rect 96528 4088 96580 4140
rect 162952 4156 163004 4208
rect 164700 4156 164752 4208
rect 405648 4156 405700 4208
rect 413836 4156 413888 4208
rect 414020 4156 414072 4208
rect 424968 4156 425020 4208
rect 495072 4156 495124 4208
rect 495532 4156 495584 4208
rect 98092 4088 98144 4140
rect 99104 4088 99156 4140
rect 352564 4088 352616 4140
rect 354956 4088 355008 4140
rect 355968 4088 356020 4140
rect 364524 4088 364576 4140
rect 365628 4088 365680 4140
rect 365720 4088 365772 4140
rect 367008 4088 367060 4140
rect 374000 4088 374052 4140
rect 375196 4088 375248 4140
rect 381176 4088 381228 4140
rect 500132 4088 500184 4140
rect 500868 4088 500920 4140
rect 501604 4088 501656 4140
rect 502524 4088 502576 4140
rect 503628 4088 503680 4140
rect 507676 4088 507728 4140
rect 508412 4088 508464 4140
rect 511264 4088 511316 4140
rect 512000 4088 512052 4140
rect 42156 4020 42208 4072
rect 64144 4020 64196 4072
rect 76748 4020 76800 4072
rect 340696 4020 340748 4072
rect 347872 4020 347924 4072
rect 348976 4020 349028 4072
rect 509332 4020 509384 4072
rect 43352 3952 43404 4004
rect 506572 3952 506624 4004
rect 30288 3884 30340 3936
rect 51816 3884 51868 3936
rect 52828 3884 52880 3936
rect 57244 3884 57296 3936
rect 76840 3884 76892 3936
rect 351368 3884 351420 3936
rect 385868 3884 385920 3936
rect 506480 3884 506532 3936
rect 26700 3816 26752 3868
rect 50344 3816 50396 3868
rect 80428 3816 80480 3868
rect 208676 3816 208728 3868
rect 209688 3816 209740 3868
rect 209872 3816 209924 3868
rect 210976 3816 211028 3868
rect 215852 3816 215904 3868
rect 216588 3816 216640 3868
rect 217048 3816 217100 3868
rect 217968 3816 218020 3868
rect 226524 3816 226576 3868
rect 227628 3816 227680 3868
rect 227720 3816 227772 3868
rect 498936 3816 498988 3868
rect 501696 3816 501748 3868
rect 25504 3748 25556 3800
rect 31024 3748 31076 3800
rect 39764 3748 39816 3800
rect 313924 3748 313976 3800
rect 315764 3748 315816 3800
rect 502248 3748 502300 3800
rect 538864 3748 538916 3800
rect 548892 3748 548944 3800
rect 31484 3680 31536 3732
rect 60004 3680 60056 3732
rect 73804 3680 73856 3732
rect 89720 3680 89772 3732
rect 91008 3680 91060 3732
rect 93308 3680 93360 3732
rect 101588 3680 101640 3732
rect 102048 3680 102100 3732
rect 103520 3680 103572 3732
rect 103980 3680 104032 3732
rect 105176 3680 105228 3732
rect 106188 3680 106240 3732
rect 106372 3680 106424 3732
rect 107568 3680 107620 3732
rect 112352 3680 112404 3732
rect 113088 3680 113140 3732
rect 115756 3680 115808 3732
rect 116860 3680 116912 3732
rect 393320 3680 393372 3732
rect 393872 3680 393924 3732
rect 567844 3680 567896 3732
rect 29092 3612 29144 3664
rect 42064 3612 42116 3664
rect 45744 3612 45796 3664
rect 397828 3612 397880 3664
rect 398748 3612 398800 3664
rect 399024 3612 399076 3664
rect 400128 3612 400180 3664
rect 406108 3612 406160 3664
rect 407028 3612 407080 3664
rect 412088 3612 412140 3664
rect 415492 3612 415544 3664
rect 431132 3612 431184 3664
rect 431868 3612 431920 3664
rect 439412 3612 439464 3664
rect 440148 3612 440200 3664
rect 444196 3612 444248 3664
rect 519636 3612 519688 3664
rect 528652 3612 528704 3664
rect 531964 3612 532016 3664
rect 17316 3544 17368 3596
rect 46296 3544 46348 3596
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 12348 3476 12400 3528
rect 8852 3408 8904 3460
rect 17224 3476 17276 3528
rect 19524 3476 19576 3528
rect 20628 3476 20680 3528
rect 23112 3476 23164 3528
rect 53104 3544 53156 3596
rect 55220 3544 55272 3596
rect 56416 3544 56468 3596
rect 60004 3544 60056 3596
rect 71044 3544 71096 3596
rect 77668 3544 77720 3596
rect 504824 3544 504876 3596
rect 522304 3544 522356 3596
rect 532240 3544 532292 3596
rect 540336 3612 540388 3664
rect 582196 3612 582248 3664
rect 46940 3476 46992 3528
rect 48964 3476 49016 3528
rect 51632 3476 51684 3528
rect 52368 3476 52420 3528
rect 58808 3476 58860 3528
rect 59268 3476 59320 3528
rect 24308 3408 24360 3460
rect 61384 3476 61436 3528
rect 62396 3476 62448 3528
rect 63408 3476 63460 3528
rect 63592 3476 63644 3528
rect 64696 3476 64748 3528
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 34980 3340 35032 3392
rect 35808 3340 35860 3392
rect 37372 3340 37424 3392
rect 38476 3340 38528 3392
rect 1676 3272 1728 3324
rect 7656 3272 7708 3324
rect 9128 3272 9180 3324
rect 36176 3272 36228 3324
rect 46204 3340 46256 3392
rect 61200 3340 61252 3392
rect 69480 3476 69532 3528
rect 70216 3476 70268 3528
rect 70676 3476 70728 3528
rect 71688 3476 71740 3528
rect 71872 3476 71924 3528
rect 72976 3476 73028 3528
rect 77484 3476 77536 3528
rect 554780 3476 554832 3528
rect 77576 3408 77628 3460
rect 569040 3408 569092 3460
rect 571432 3544 571484 3596
rect 572628 3544 572680 3596
rect 576216 3408 576268 3460
rect 68284 3340 68336 3392
rect 249156 3340 249208 3392
rect 249708 3340 249760 3392
rect 250352 3340 250404 3392
rect 251088 3340 251140 3392
rect 252652 3340 252704 3392
rect 253848 3340 253900 3392
rect 283656 3340 283708 3392
rect 284208 3340 284260 3392
rect 285956 3340 286008 3392
rect 286968 3340 287020 3392
rect 293132 3340 293184 3392
rect 293868 3340 293920 3392
rect 295524 3340 295576 3392
rect 296628 3340 296680 3392
rect 303804 3340 303856 3392
rect 304908 3340 304960 3392
rect 307760 3340 307812 3392
rect 321652 3340 321704 3392
rect 322756 3340 322808 3392
rect 324044 3340 324096 3392
rect 326436 3340 326488 3392
rect 326988 3340 327040 3392
rect 327632 3340 327684 3392
rect 328368 3340 328420 3392
rect 328828 3340 328880 3392
rect 329748 3340 329800 3392
rect 330024 3340 330076 3392
rect 331128 3340 331180 3392
rect 331220 3340 331272 3392
rect 332508 3340 332560 3392
rect 339500 3340 339552 3392
rect 340788 3340 340840 3392
rect 344284 3340 344336 3392
rect 388260 3340 388312 3392
rect 505100 3340 505152 3392
rect 54024 3272 54076 3324
rect 291292 3272 291344 3324
rect 307024 3272 307076 3324
rect 307392 3272 307444 3324
rect 493324 3272 493376 3324
rect 494152 3272 494204 3324
rect 9220 3204 9272 3256
rect 77392 3204 77444 3256
rect 65984 3136 66036 3188
rect 69664 3136 69716 3188
rect 78128 3136 78180 3188
rect 214656 3136 214708 3188
rect 265808 3204 265860 3256
rect 266268 3204 266320 3256
rect 74264 3068 74316 3120
rect 75184 3068 75236 3120
rect 85028 3068 85080 3120
rect 12440 3000 12492 3052
rect 13728 3000 13780 3052
rect 20720 3000 20772 3052
rect 22008 3000 22060 3052
rect 77208 3000 77260 3052
rect 129740 3068 129792 3120
rect 130200 3068 130252 3120
rect 136088 3068 136140 3120
rect 136548 3068 136600 3120
rect 122932 3000 122984 3052
rect 139676 3068 139728 3120
rect 140688 3068 140740 3120
rect 142160 3068 142212 3120
rect 143264 3068 143316 3120
rect 145656 3068 145708 3120
rect 146208 3068 146260 3120
rect 146392 3068 146444 3120
rect 146852 3068 146904 3120
rect 153200 3068 153252 3120
rect 153936 3068 153988 3120
rect 77760 2932 77812 2984
rect 99380 2932 99432 2984
rect 108948 2932 109000 2984
rect 118700 2932 118752 2984
rect 4068 2864 4120 2916
rect 8944 2864 8996 2916
rect 85120 2864 85172 2916
rect 157524 3000 157576 3052
rect 158628 3000 158680 3052
rect 164700 3000 164752 3052
rect 165528 3000 165580 3052
rect 167184 3000 167236 3052
rect 168196 3000 168248 3052
rect 172980 3000 173032 3052
rect 173808 3000 173860 3052
rect 176660 3000 176712 3052
rect 177764 3000 177816 3052
rect 165896 2932 165948 2984
rect 179420 3068 179472 3120
rect 180156 3068 180208 3120
rect 182548 3068 182600 3120
rect 183468 3068 183520 3120
rect 187700 3068 187752 3120
rect 188436 3068 188488 3120
rect 189632 3068 189684 3120
rect 190368 3068 190420 3120
rect 192024 3068 192076 3120
rect 193128 3068 193180 3120
rect 198004 3068 198056 3120
rect 198648 3068 198700 3120
rect 199200 3068 199252 3120
rect 199936 3068 199988 3120
rect 200396 3068 200448 3120
rect 201408 3068 201460 3120
rect 201500 3068 201552 3120
rect 202696 3068 202748 3120
rect 232504 3068 232556 3120
rect 233148 3068 233200 3120
rect 236000 3068 236052 3120
rect 237196 3068 237248 3120
rect 239588 3068 239640 3120
rect 240048 3068 240100 3120
rect 240784 3068 240836 3120
rect 241428 3068 241480 3120
rect 241980 3068 242032 3120
rect 242808 3068 242860 3120
rect 234804 3000 234856 3052
rect 255044 3136 255096 3188
rect 274088 3204 274140 3256
rect 274548 3204 274600 3256
rect 277676 3204 277728 3256
rect 278688 3204 278740 3256
rect 287152 3204 287204 3256
rect 479524 3204 479576 3256
rect 483480 3204 483532 3256
rect 484308 3204 484360 3256
rect 485780 3204 485832 3256
rect 487068 3204 487120 3256
rect 276480 3136 276532 3188
rect 305092 3136 305144 3188
rect 476764 3136 476816 3188
rect 477500 3136 477552 3188
rect 356152 3068 356204 3120
rect 387800 3068 387852 3120
rect 402244 3068 402296 3120
rect 411168 3068 411220 3120
rect 421564 3068 421616 3120
rect 422208 3068 422260 3120
rect 440608 3068 440660 3120
rect 447784 3068 447836 3120
rect 503076 3136 503128 3188
rect 510712 3204 510764 3256
rect 507952 3136 508004 3188
rect 508044 3068 508096 3120
rect 296720 3000 296772 3052
rect 297916 3000 297968 3052
rect 450176 3000 450228 3052
rect 509240 3000 509292 3052
rect 76932 2796 76984 2848
rect 133788 2796 133840 2848
rect 158720 2864 158772 2916
rect 451280 2932 451332 2984
rect 452476 2932 452528 2984
rect 456064 2932 456116 2984
rect 456708 2932 456760 2984
rect 466828 2932 466880 2984
rect 467748 2932 467800 2984
rect 471520 2932 471572 2984
rect 506388 2932 506440 2984
rect 471152 2864 471204 2916
rect 484584 2864 484636 2916
rect 489368 2864 489420 2916
rect 510620 2864 510672 2916
rect 571984 2864 572036 2916
rect 578608 2864 578660 2916
rect 142068 2796 142120 2848
rect 358820 2796 358872 2848
rect 384672 2796 384724 2848
rect 384948 2796 385000 2848
rect 481088 2796 481140 2848
rect 85580 2728 85632 2780
rect 95148 2728 95200 2780
rect 96896 2728 96948 2780
rect 161388 2728 161440 2780
rect 162308 2728 162360 2780
rect 359740 2728 359792 2780
rect 508228 2796 508280 2848
rect 563060 2728 563112 2780
rect 564348 2728 564400 2780
rect 305000 1232 305052 1284
rect 306196 1232 306248 1284
rect 80244 552 80296 604
rect 80336 552 80388 604
rect 92112 552 92164 604
rect 92388 552 92440 604
rect 100484 595 100536 604
rect 100484 561 100493 595
rect 100493 561 100527 595
rect 100527 561 100536 595
rect 100484 552 100536 561
rect 111156 595 111208 604
rect 111156 561 111165 595
rect 111165 561 111199 595
rect 111199 561 111208 595
rect 111156 552 111208 561
rect 134892 595 134944 604
rect 134892 561 134901 595
rect 134901 561 134935 595
rect 134935 561 134944 595
rect 134892 552 134944 561
rect 186044 595 186096 604
rect 186044 561 186053 595
rect 186053 561 186087 595
rect 186087 561 186096 595
rect 186044 552 186096 561
rect 190368 552 190420 604
rect 190828 552 190880 604
rect 205640 552 205692 604
rect 206284 552 206336 604
rect 212540 552 212592 604
rect 213460 552 213512 604
rect 247960 552 248012 604
rect 248328 552 248380 604
rect 258632 595 258684 604
rect 258632 561 258641 595
rect 258641 561 258675 595
rect 258675 561 258684 595
rect 258632 552 258684 561
rect 289544 552 289596 604
rect 289912 552 289964 604
rect 370412 595 370464 604
rect 370412 561 370421 595
rect 370421 561 370455 595
rect 370455 561 370464 595
rect 370412 552 370464 561
rect 371608 595 371660 604
rect 371608 561 371617 595
rect 371617 561 371651 595
rect 371651 561 371660 595
rect 371608 552 371660 561
rect 372804 595 372856 604
rect 372804 561 372813 595
rect 372813 561 372847 595
rect 372847 561 372856 595
rect 372804 552 372856 561
rect 377588 595 377640 604
rect 377588 561 377597 595
rect 377597 561 377631 595
rect 377631 561 377640 595
rect 377588 552 377640 561
rect 378784 595 378836 604
rect 378784 561 378793 595
rect 378793 561 378827 595
rect 378827 561 378836 595
rect 378784 552 378836 561
rect 396080 552 396132 604
rect 396632 552 396684 604
rect 412640 552 412692 604
rect 413284 552 413336 604
rect 428740 595 428792 604
rect 428740 561 428749 595
rect 428749 561 428783 595
rect 428783 561 428792 595
rect 428740 552 428792 561
rect 437020 595 437072 604
rect 437020 561 437029 595
rect 437029 561 437063 595
rect 437063 561 437072 595
rect 437020 552 437072 561
rect 437480 552 437532 604
rect 438216 552 438268 604
rect 444472 552 444524 604
rect 445392 552 445444 604
rect 445760 552 445812 604
rect 446588 552 446640 604
rect 448520 552 448572 604
rect 448980 552 449032 604
rect 453672 552 453724 604
rect 453948 552 454000 604
rect 454040 552 454092 604
rect 454868 552 454920 604
rect 473360 552 473412 604
rect 473912 552 473964 604
rect 492680 552 492732 604
rect 492956 552 493008 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 506664 552 506716 604
rect 507216 552 507268 604
rect 512092 552 512144 604
rect 513196 552 513248 604
rect 513380 552 513432 604
rect 514392 552 514444 604
rect 514760 552 514812 604
rect 515588 552 515640 604
rect 576860 552 576912 604
rect 577412 552 577464 604
rect 579620 552 579672 604
rect 579804 552 579856 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 19984 700324 20036 700330
rect 19984 700266 20036 700272
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 9312 681760 9364 681766
rect 9312 681702 9364 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 8852 610020 8904 610026
rect 8852 609962 8904 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 6184 582412 6236 582418
rect 6184 582354 6236 582360
rect 3424 581868 3476 581874
rect 3424 581810 3476 581816
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 2870 509960 2926 509969
rect 2870 509895 2926 509904
rect 2884 509318 2912 509895
rect 2872 509312 2924 509318
rect 2872 509254 2924 509260
rect 3332 481568 3384 481574
rect 3332 481510 3384 481516
rect 3344 481137 3372 481510
rect 3330 481128 3386 481137
rect 3330 481063 3386 481072
rect 2964 424244 3016 424250
rect 2964 424186 3016 424192
rect 2976 423745 3004 424186
rect 2962 423736 3018 423745
rect 2962 423671 3018 423680
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3344 394738 3372 394975
rect 3332 394732 3384 394738
rect 3332 394674 3384 394680
rect 3054 380624 3110 380633
rect 3054 380559 3110 380568
rect 3068 379574 3096 380559
rect 3056 379568 3108 379574
rect 3056 379510 3108 379516
rect 2962 337512 3018 337521
rect 2962 337447 3018 337456
rect 2976 336802 3004 337447
rect 2964 336796 3016 336802
rect 2964 336738 3016 336744
rect 3332 324284 3384 324290
rect 3332 324226 3384 324232
rect 3344 323105 3372 324226
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3240 294772 3292 294778
rect 3240 294714 3292 294720
rect 3252 294409 3280 294714
rect 3238 294400 3294 294409
rect 3238 294335 3294 294344
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 2792 200297 2820 280055
rect 2962 265704 3018 265713
rect 2962 265639 3018 265648
rect 2976 264994 3004 265639
rect 2964 264988 3016 264994
rect 2964 264930 3016 264936
rect 3330 251288 3386 251297
rect 3330 251223 3332 251232
rect 3384 251223 3386 251232
rect 3332 251194 3384 251200
rect 3240 237380 3292 237386
rect 3240 237322 3292 237328
rect 3252 237017 3280 237322
rect 3238 237008 3294 237017
rect 3238 236943 3294 236952
rect 3332 223576 3384 223582
rect 3332 223518 3384 223524
rect 3344 222601 3372 223518
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 3148 208344 3200 208350
rect 3148 208286 3200 208292
rect 3160 208185 3188 208286
rect 3146 208176 3202 208185
rect 3146 208111 3202 208120
rect 2778 200288 2834 200297
rect 2778 200223 2834 200232
rect 3436 193905 3464 581810
rect 4804 581596 4856 581602
rect 4804 581538 4856 581544
rect 3514 567352 3570 567361
rect 3514 567287 3570 567296
rect 3528 567254 3556 567287
rect 3516 567248 3568 567254
rect 3516 567190 3568 567196
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3528 538286 3556 538591
rect 3516 538280 3568 538286
rect 3516 538222 3568 538228
rect 3516 496800 3568 496806
rect 3516 496742 3568 496748
rect 3528 495553 3556 496742
rect 3514 495544 3570 495553
rect 3514 495479 3570 495488
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 3422 193896 3478 193905
rect 3422 193831 3478 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3424 165572 3476 165578
rect 3424 165514 3476 165520
rect 3436 165073 3464 165514
rect 3422 165064 3478 165073
rect 3422 164999 3478 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3422 136368 3478 136377
rect 3422 136303 3478 136312
rect 3436 120970 3464 136303
rect 3528 122210 3556 437951
rect 3606 366208 3662 366217
rect 3606 366143 3662 366152
rect 3620 365770 3648 366143
rect 3608 365764 3660 365770
rect 3608 365706 3660 365712
rect 3528 122182 3740 122210
rect 3514 122088 3570 122097
rect 3514 122023 3570 122032
rect 3528 121582 3556 122023
rect 3516 121576 3568 121582
rect 3516 121518 3568 121524
rect 3712 121174 3740 122182
rect 3700 121168 3752 121174
rect 3700 121110 3752 121116
rect 3424 120964 3476 120970
rect 3424 120906 3476 120912
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3422 80064 3478 80073
rect 3422 79999 3478 80008
rect 3436 78985 3464 79999
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 2780 64592 2832 64598
rect 2778 64560 2780 64569
rect 2832 64560 2834 64569
rect 2778 64495 2834 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3148 35896 3200 35902
rect 3146 35864 3148 35873
rect 3200 35864 3202 35873
rect 3146 35799 3202 35808
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 4816 3534 4844 581538
rect 4896 407176 4948 407182
rect 4896 407118 4948 407124
rect 4908 64598 4936 407118
rect 4896 64592 4948 64598
rect 4896 64534 4948 64540
rect 6196 35902 6224 582354
rect 8758 579728 8814 579737
rect 8758 579663 8814 579672
rect 8772 481574 8800 579663
rect 8760 481568 8812 481574
rect 8760 481510 8812 481516
rect 8864 478854 8892 609962
rect 8944 582752 8996 582758
rect 8944 582694 8996 582700
rect 8852 478848 8904 478854
rect 8852 478790 8904 478796
rect 8852 336796 8904 336802
rect 8852 336738 8904 336744
rect 6828 168428 6880 168434
rect 6828 168370 6880 168376
rect 6184 35896 6236 35902
rect 6184 35838 6236 35844
rect 5262 4856 5318 4865
rect 5262 4791 5318 4800
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 1676 3324 1728 3330
rect 1676 3266 1728 3272
rect 1688 480 1716 3266
rect 2884 480 2912 3470
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 480 4108 2858
rect 5276 480 5304 4791
rect 6840 626 6868 168370
rect 8864 121378 8892 336738
rect 8852 121372 8904 121378
rect 8852 121314 8904 121320
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 7656 3324 7708 3330
rect 7656 3266 7708 3272
rect 6472 598 6868 626
rect 6472 480 6500 598
rect 7668 480 7696 3266
rect 8864 480 8892 3402
rect 8956 2922 8984 582694
rect 9128 581664 9180 581670
rect 9128 581606 9180 581612
rect 9036 581256 9088 581262
rect 9036 581198 9088 581204
rect 9048 4146 9076 581198
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9140 3330 9168 581606
rect 9220 581392 9272 581398
rect 9220 581334 9272 581340
rect 9128 3324 9180 3330
rect 9128 3266 9180 3272
rect 9232 3262 9260 581334
rect 9324 121446 9352 681702
rect 15936 652792 15988 652798
rect 15936 652734 15988 652740
rect 14464 623824 14516 623830
rect 14464 623766 14516 623772
rect 10416 583228 10468 583234
rect 10416 583170 10468 583176
rect 9496 583160 9548 583166
rect 9496 583102 9548 583108
rect 9404 538280 9456 538286
rect 9404 538222 9456 538228
rect 9312 121440 9364 121446
rect 9312 121382 9364 121388
rect 9416 120902 9444 538222
rect 9508 294778 9536 583102
rect 9588 582480 9640 582486
rect 9588 582422 9640 582428
rect 9600 424250 9628 582422
rect 10324 581528 10376 581534
rect 10324 581470 10376 581476
rect 9588 424244 9640 424250
rect 9588 424186 9640 424192
rect 9588 394732 9640 394738
rect 9588 394674 9640 394680
rect 9496 294772 9548 294778
rect 9496 294714 9548 294720
rect 9600 121650 9628 394674
rect 10336 151774 10364 581470
rect 10428 165578 10456 583170
rect 10600 583092 10652 583098
rect 10600 583034 10652 583040
rect 10508 582276 10560 582282
rect 10508 582218 10560 582224
rect 10520 180810 10548 582218
rect 10612 208350 10640 583034
rect 10692 582684 10744 582690
rect 10692 582626 10744 582632
rect 10704 223582 10732 582626
rect 12348 436144 12400 436150
rect 12348 436086 12400 436092
rect 10968 372632 11020 372638
rect 10968 372574 11020 372580
rect 10692 223576 10744 223582
rect 10692 223518 10744 223524
rect 10600 208344 10652 208350
rect 10600 208286 10652 208292
rect 10508 180804 10560 180810
rect 10508 180746 10560 180752
rect 10416 165572 10468 165578
rect 10416 165514 10468 165520
rect 10324 151768 10376 151774
rect 10324 151710 10376 151716
rect 9588 121644 9640 121650
rect 9588 121586 9640 121592
rect 9404 120896 9456 120902
rect 9404 120838 9456 120844
rect 10980 3534 11008 372574
rect 12360 3534 12388 436086
rect 14476 278730 14504 623766
rect 15844 582820 15896 582826
rect 15844 582762 15896 582768
rect 14464 278724 14516 278730
rect 14464 278666 14516 278672
rect 14464 251252 14516 251258
rect 14464 251194 14516 251200
rect 14476 183530 14504 251194
rect 14464 183524 14516 183530
rect 14464 183466 14516 183472
rect 13728 164280 13780 164286
rect 13728 164222 13780 164228
rect 13634 101416 13690 101425
rect 13634 101351 13690 101360
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 9220 3256 9272 3262
rect 9220 3198 9272 3204
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 10060 480 10088 3470
rect 11256 480 11284 3470
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 480 12480 2994
rect 13648 480 13676 101351
rect 13740 3058 13768 164222
rect 15108 120080 15160 120086
rect 15108 120022 15160 120028
rect 15120 3346 15148 120022
rect 15856 51066 15884 582762
rect 15948 342242 15976 652734
rect 17224 509312 17276 509318
rect 17224 509254 17276 509260
rect 15936 342236 15988 342242
rect 15936 342178 15988 342184
rect 17236 333946 17264 509254
rect 17224 333940 17276 333946
rect 17224 333882 17276 333888
rect 17224 329860 17276 329866
rect 17224 329802 17276 329808
rect 17236 309126 17264 329802
rect 17224 309120 17276 309126
rect 17224 309062 17276 309068
rect 19996 176662 20024 700266
rect 24320 699718 24348 703520
rect 40512 700534 40540 703520
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 72988 700330 73016 703520
rect 78220 700732 78272 700738
rect 78220 700674 78272 700680
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 77944 700324 77996 700330
rect 77944 700266 77996 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 21364 379568 21416 379574
rect 21364 379510 21416 379516
rect 21376 362914 21404 379510
rect 21364 362908 21416 362914
rect 21364 362850 21416 362856
rect 19984 176656 20036 176662
rect 19984 176598 20036 176604
rect 24780 121242 24808 699654
rect 31116 594856 31168 594862
rect 31116 594798 31168 594804
rect 31024 584316 31076 584322
rect 31024 584258 31076 584264
rect 24768 121236 24820 121242
rect 24768 121178 24820 121184
rect 22008 119944 22060 119950
rect 22008 119886 22060 119892
rect 17224 119876 17276 119882
rect 17224 119818 17276 119824
rect 15844 51060 15896 51066
rect 15844 51002 15896 51008
rect 16026 4992 16082 5001
rect 16026 4927 16082 4936
rect 14844 3318 15148 3346
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14844 480 14872 3318
rect 16040 480 16068 4927
rect 17236 3534 17264 119818
rect 20628 119400 20680 119406
rect 20628 119342 20680 119348
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17328 1850 17356 3538
rect 17236 1822 17356 1850
rect 17236 480 17264 1822
rect 18340 480 18368 7822
rect 20640 3534 20668 119342
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 19536 480 19564 3470
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20732 480 20760 2994
rect 21928 480 21956 7686
rect 22020 3058 22048 119886
rect 28908 119536 28960 119542
rect 28908 119478 28960 119484
rect 26700 3868 26752 3874
rect 26700 3810 26752 3816
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 23124 480 23152 3470
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 24320 480 24348 3402
rect 25516 480 25544 3742
rect 26712 480 26740 3810
rect 28920 3398 28948 119478
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 480 27936 3334
rect 29104 480 29132 3606
rect 30300 480 30328 3878
rect 31036 3806 31064 584258
rect 31128 120358 31156 594798
rect 46204 585132 46256 585138
rect 46204 585074 46256 585080
rect 42064 583908 42116 583914
rect 42064 583850 42116 583856
rect 35808 583500 35860 583506
rect 35808 583442 35860 583448
rect 33784 567248 33836 567254
rect 33784 567190 33836 567196
rect 33796 121038 33824 567190
rect 33876 357468 33928 357474
rect 33876 357410 33928 357416
rect 33784 121032 33836 121038
rect 33784 120974 33836 120980
rect 31116 120352 31168 120358
rect 31116 120294 31168 120300
rect 33888 93838 33916 357410
rect 33876 93832 33928 93838
rect 33876 93774 33928 93780
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 31024 3800 31076 3806
rect 31024 3742 31076 3748
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31496 480 31524 3674
rect 32692 480 32720 4082
rect 33888 480 33916 7890
rect 35820 3398 35848 583442
rect 38568 427848 38620 427854
rect 38568 427790 38620 427796
rect 38476 119332 38528 119338
rect 38476 119274 38528 119280
rect 38488 3398 38516 119274
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 38476 3392 38528 3398
rect 38476 3334 38528 3340
rect 34992 480 35020 3334
rect 36176 3324 36228 3330
rect 36176 3266 36228 3272
rect 36188 480 36216 3266
rect 37384 480 37412 3334
rect 38580 480 38608 427790
rect 41328 248464 41380 248470
rect 41328 248406 41380 248412
rect 39764 3800 39816 3806
rect 39764 3742 39816 3748
rect 39776 480 39804 3742
rect 41340 3482 41368 248406
rect 42076 3670 42104 583850
rect 42156 552084 42208 552090
rect 42156 552026 42208 552032
rect 42168 120834 42196 552026
rect 42248 365764 42300 365770
rect 42248 365706 42300 365712
rect 42260 121310 42288 365706
rect 42248 121304 42300 121310
rect 42248 121246 42300 121252
rect 42156 120828 42208 120834
rect 42156 120770 42208 120776
rect 44548 7676 44600 7682
rect 44548 7618 44600 7624
rect 42156 4072 42208 4078
rect 42156 4014 42208 4020
rect 42064 3664 42116 3670
rect 42064 3606 42116 3612
rect 40972 3454 41368 3482
rect 40972 480 41000 3454
rect 42168 480 42196 4014
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 43364 480 43392 3946
rect 44560 480 44588 7618
rect 45744 3664 45796 3670
rect 45744 3606 45796 3612
rect 45756 480 45784 3606
rect 46216 3398 46244 585074
rect 71044 584996 71096 585002
rect 71044 584938 71096 584944
rect 57244 584928 57296 584934
rect 57244 584870 57296 584876
rect 50344 584452 50396 584458
rect 50344 584394 50396 584400
rect 48228 581936 48280 581942
rect 48228 581878 48280 581884
rect 46296 119468 46348 119474
rect 46296 119410 46348 119416
rect 46308 3602 46336 119410
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 46204 3392 46256 3398
rect 46204 3334 46256 3340
rect 46952 480 46980 3470
rect 48240 626 48268 581878
rect 48964 572756 49016 572762
rect 48964 572698 49016 572704
rect 48976 3534 49004 572698
rect 49608 379568 49660 379574
rect 49608 379510 49660 379516
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49620 626 49648 379510
rect 50356 3874 50384 584394
rect 53104 584384 53156 584390
rect 53104 584326 53156 584332
rect 51724 584180 51776 584186
rect 51724 584122 51776 584128
rect 50528 7608 50580 7614
rect 50528 7550 50580 7556
rect 50344 3868 50396 3874
rect 50344 3810 50396 3816
rect 48148 598 48268 626
rect 49344 598 49648 626
rect 48148 480 48176 598
rect 49344 480 49372 598
rect 50540 480 50568 7550
rect 51736 4146 51764 584122
rect 52368 581732 52420 581738
rect 52368 581674 52420 581680
rect 51816 119740 51868 119746
rect 51816 119682 51868 119688
rect 51724 4140 51776 4146
rect 51724 4082 51776 4088
rect 51828 3942 51856 119682
rect 51816 3936 51868 3942
rect 51816 3878 51868 3884
rect 52380 3534 52408 581674
rect 52828 3936 52880 3942
rect 52828 3878 52880 3884
rect 51632 3528 51684 3534
rect 51632 3470 51684 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 51644 480 51672 3470
rect 52840 480 52868 3878
rect 53116 3602 53144 584326
rect 56508 150476 56560 150482
rect 56508 150418 56560 150424
rect 56416 17264 56468 17270
rect 56416 17206 56468 17212
rect 56428 3602 56456 17206
rect 53104 3596 53156 3602
rect 53104 3538 53156 3544
rect 55220 3596 55272 3602
rect 55220 3538 55272 3544
rect 56416 3596 56468 3602
rect 56416 3538 56468 3544
rect 54024 3324 54076 3330
rect 54024 3266 54076 3272
rect 54036 480 54064 3266
rect 55232 480 55260 3538
rect 56520 3482 56548 150418
rect 57256 3942 57284 584870
rect 61384 584656 61436 584662
rect 61384 584598 61436 584604
rect 60004 584588 60056 584594
rect 60004 584530 60056 584536
rect 57888 280220 57940 280226
rect 57888 280162 57940 280168
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57900 3346 57928 280162
rect 59268 119672 59320 119678
rect 59268 119614 59320 119620
rect 59280 3534 59308 119614
rect 60016 3738 60044 584530
rect 60004 3732 60056 3738
rect 60004 3674 60056 3680
rect 60004 3596 60056 3602
rect 60004 3538 60056 3544
rect 58808 3528 58860 3534
rect 58808 3470 58860 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 57624 3318 57928 3346
rect 57624 480 57652 3318
rect 58820 480 58848 3470
rect 60016 480 60044 3538
rect 61396 3534 61424 584598
rect 64144 584520 64196 584526
rect 64144 584462 64196 584468
rect 63408 343664 63460 343670
rect 63408 343606 63460 343612
rect 63420 3534 63448 343606
rect 64156 4078 64184 584462
rect 64788 582548 64840 582554
rect 64788 582490 64840 582496
rect 64694 18592 64750 18601
rect 64694 18527 64750 18536
rect 64144 4072 64196 4078
rect 64144 4014 64196 4020
rect 64708 3534 64736 18527
rect 61384 3528 61436 3534
rect 61384 3470 61436 3476
rect 62396 3528 62448 3534
rect 62396 3470 62448 3476
rect 63408 3528 63460 3534
rect 63408 3470 63460 3476
rect 63592 3528 63644 3534
rect 63592 3470 63644 3476
rect 64696 3528 64748 3534
rect 64696 3470 64748 3476
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 61212 480 61240 3334
rect 62408 480 62436 3470
rect 63604 480 63632 3470
rect 64800 480 64828 582490
rect 67548 581460 67600 581466
rect 67548 581402 67600 581408
rect 65984 3188 66036 3194
rect 65984 3130 66036 3136
rect 65996 480 66024 3130
rect 67560 626 67588 581402
rect 70308 558952 70360 558958
rect 70308 558894 70360 558900
rect 69664 393372 69716 393378
rect 69664 393314 69716 393320
rect 69480 3528 69532 3534
rect 69480 3470 69532 3476
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3334
rect 69492 480 69520 3470
rect 69676 3194 69704 393314
rect 70216 309188 70268 309194
rect 70216 309130 70268 309136
rect 70228 3534 70256 309130
rect 70320 4049 70348 558894
rect 70306 4040 70362 4049
rect 70306 3975 70362 3984
rect 71056 3602 71084 584938
rect 77024 584724 77076 584730
rect 77024 584666 77076 584672
rect 76932 584248 76984 584254
rect 76932 584190 76984 584196
rect 75184 584112 75236 584118
rect 75184 584054 75236 584060
rect 73804 583976 73856 583982
rect 73804 583918 73856 583924
rect 73068 582140 73120 582146
rect 73068 582082 73120 582088
rect 71688 119808 71740 119814
rect 71688 119750 71740 119756
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 71700 3534 71728 119750
rect 72976 118924 73028 118930
rect 72976 118866 73028 118872
rect 72988 3534 73016 118866
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 70676 3528 70728 3534
rect 70676 3470 70728 3476
rect 71688 3528 71740 3534
rect 71688 3470 71740 3476
rect 71872 3528 71924 3534
rect 71872 3470 71924 3476
rect 72976 3528 73028 3534
rect 72976 3470 73028 3476
rect 69664 3188 69716 3194
rect 69664 3130 69716 3136
rect 70688 480 70716 3470
rect 71884 480 71912 3470
rect 73080 480 73108 582082
rect 73620 342236 73672 342242
rect 73620 342178 73672 342184
rect 73632 341057 73660 342178
rect 73618 341048 73674 341057
rect 73618 340983 73674 340992
rect 73816 3738 73844 583918
rect 74446 513768 74502 513777
rect 74446 513703 74502 513712
rect 74354 503160 74410 503169
rect 74354 503095 74410 503104
rect 74170 358728 74226 358737
rect 74170 358663 74226 358672
rect 74184 357474 74212 358663
rect 74172 357468 74224 357474
rect 74172 357410 74224 357416
rect 74368 6322 74396 503095
rect 74356 6316 74408 6322
rect 74356 6258 74408 6264
rect 74460 6186 74488 513703
rect 75090 436248 75146 436257
rect 75090 436183 75146 436192
rect 75104 436150 75132 436183
rect 75092 436144 75144 436150
rect 75092 436086 75144 436092
rect 74448 6180 74500 6186
rect 74448 6122 74500 6128
rect 73804 3732 73856 3738
rect 73804 3674 73856 3680
rect 75196 3126 75224 584054
rect 75828 583432 75880 583438
rect 75828 583374 75880 583380
rect 75276 583296 75328 583302
rect 75276 583238 75328 583244
rect 75288 324290 75316 583238
rect 75276 324284 75328 324290
rect 75276 324226 75328 324232
rect 75642 281208 75698 281217
rect 75642 281143 75698 281152
rect 75656 280226 75684 281143
rect 75644 280220 75696 280226
rect 75644 280162 75696 280168
rect 75460 278724 75512 278730
rect 75460 278666 75512 278672
rect 75472 277681 75500 278666
rect 75458 277672 75514 277681
rect 75458 277607 75514 277616
rect 75840 4842 75868 583374
rect 76838 450392 76894 450401
rect 76838 450327 76894 450336
rect 76746 418568 76802 418577
rect 76746 418503 76802 418512
rect 76470 333976 76526 333985
rect 76470 333911 76472 333920
rect 76524 333911 76526 333920
rect 76472 333882 76524 333888
rect 76654 288280 76710 288289
rect 76654 288215 76710 288224
rect 76010 249656 76066 249665
rect 76010 249591 76066 249600
rect 76024 248470 76052 249591
rect 76012 248464 76064 248470
rect 76012 248406 76064 248412
rect 76562 228440 76618 228449
rect 76562 228375 76618 228384
rect 76378 201920 76434 201929
rect 76378 201855 76434 201864
rect 76392 198121 76420 201855
rect 76472 200796 76524 200802
rect 76472 200738 76524 200744
rect 76378 198112 76434 198121
rect 76378 198047 76434 198056
rect 76484 191010 76512 200738
rect 76472 191004 76524 191010
rect 76472 190946 76524 190952
rect 76576 77246 76604 228375
rect 76564 77240 76616 77246
rect 76564 77182 76616 77188
rect 76564 11892 76616 11898
rect 76564 11834 76616 11840
rect 76576 6934 76604 11834
rect 76564 6928 76616 6934
rect 76564 6870 76616 6876
rect 76668 6882 76696 288215
rect 76760 11778 76788 418503
rect 76852 11898 76880 450327
rect 76944 200802 76972 584190
rect 76932 200796 76984 200802
rect 76932 200738 76984 200744
rect 76932 199572 76984 199578
rect 76932 199514 76984 199520
rect 76944 191146 76972 199514
rect 76932 191140 76984 191146
rect 76932 191082 76984 191088
rect 76932 191004 76984 191010
rect 76932 190946 76984 190952
rect 76944 122806 76972 190946
rect 76932 122800 76984 122806
rect 76932 122742 76984 122748
rect 76840 11892 76892 11898
rect 76840 11834 76892 11840
rect 76760 11750 76880 11778
rect 76668 6854 76788 6882
rect 75472 4814 75868 4842
rect 74264 3120 74316 3126
rect 74264 3062 74316 3068
rect 75184 3120 75236 3126
rect 75184 3062 75236 3068
rect 74276 480 74304 3062
rect 75472 480 75500 4814
rect 76656 4140 76708 4146
rect 76656 4082 76708 4088
rect 76668 480 76696 4082
rect 76760 4078 76788 6854
rect 76748 4072 76800 4078
rect 76748 4014 76800 4020
rect 76852 3942 76880 11750
rect 76932 6928 76984 6934
rect 76932 6870 76984 6876
rect 76840 3936 76892 3942
rect 76840 3878 76892 3884
rect 76944 2854 76972 6870
rect 77036 6662 77064 584666
rect 77208 584044 77260 584050
rect 77208 583986 77260 583992
rect 77116 583364 77168 583370
rect 77116 583306 77168 583312
rect 77128 199578 77156 583306
rect 77116 199572 77168 199578
rect 77116 199514 77168 199520
rect 77116 191140 77168 191146
rect 77116 191082 77168 191088
rect 77024 6656 77076 6662
rect 77024 6598 77076 6604
rect 77128 4146 77156 191082
rect 77116 4140 77168 4146
rect 77116 4082 77168 4088
rect 77220 3058 77248 583986
rect 77760 583024 77812 583030
rect 77760 582966 77812 582972
rect 77576 478848 77628 478854
rect 77576 478790 77628 478796
rect 77588 478417 77616 478790
rect 77574 478408 77630 478417
rect 77574 478343 77630 478352
rect 77574 429176 77630 429185
rect 77574 429111 77630 429120
rect 77588 427854 77616 429111
rect 77576 427848 77628 427854
rect 77576 427790 77628 427796
rect 77666 407960 77722 407969
rect 77666 407895 77722 407904
rect 77680 407182 77708 407895
rect 77668 407176 77720 407182
rect 77668 407118 77720 407124
rect 77574 379944 77630 379953
rect 77574 379879 77630 379888
rect 77588 379574 77616 379879
rect 77576 379568 77628 379574
rect 77576 379510 77628 379516
rect 77574 372872 77630 372881
rect 77574 372807 77630 372816
rect 77588 372638 77616 372807
rect 77576 372632 77628 372638
rect 77576 372574 77628 372580
rect 77576 362908 77628 362914
rect 77576 362850 77628 362856
rect 77588 362273 77616 362850
rect 77574 362264 77630 362273
rect 77574 362199 77630 362208
rect 77574 344584 77630 344593
rect 77574 344519 77630 344528
rect 77588 343670 77616 344519
rect 77576 343664 77628 343670
rect 77576 343606 77628 343612
rect 77574 330440 77630 330449
rect 77574 330375 77630 330384
rect 77588 329866 77616 330375
rect 77576 329860 77628 329866
rect 77576 329802 77628 329808
rect 77666 323640 77722 323649
rect 77666 323575 77722 323584
rect 77574 309496 77630 309505
rect 77574 309431 77630 309440
rect 77588 309194 77616 309431
rect 77576 309188 77628 309194
rect 77576 309130 77628 309136
rect 77574 295488 77630 295497
rect 77574 295423 77630 295432
rect 77588 284646 77616 295423
rect 77576 284640 77628 284646
rect 77576 284582 77628 284588
rect 77574 267064 77630 267073
rect 77574 266999 77630 267008
rect 77300 264988 77352 264994
rect 77300 264930 77352 264936
rect 77312 120766 77340 264930
rect 77482 256728 77538 256737
rect 77482 256663 77538 256672
rect 77390 247888 77446 247897
rect 77390 247823 77446 247832
rect 77404 237697 77432 247823
rect 77390 237688 77446 237697
rect 77390 237623 77446 237632
rect 77392 171148 77444 171154
rect 77392 171090 77444 171096
rect 77300 120760 77352 120766
rect 77300 120702 77352 120708
rect 77404 3262 77432 171090
rect 77496 3534 77524 256663
rect 77484 3528 77536 3534
rect 77484 3470 77536 3476
rect 77588 3466 77616 266999
rect 77680 3602 77708 323575
rect 77772 237386 77800 582966
rect 77852 400240 77904 400246
rect 77852 400182 77904 400188
rect 77760 237380 77812 237386
rect 77760 237322 77812 237328
rect 77760 216708 77812 216714
rect 77760 216650 77812 216656
rect 77772 6254 77800 216650
rect 77760 6248 77812 6254
rect 77760 6190 77812 6196
rect 77864 6066 77892 400182
rect 77956 129713 77984 700266
rect 78126 506696 78182 506705
rect 78126 506631 78182 506640
rect 78034 499624 78090 499633
rect 78034 499559 78090 499568
rect 77942 129704 77998 129713
rect 77942 129639 77998 129648
rect 77772 6038 77892 6066
rect 77668 3596 77720 3602
rect 77668 3538 77720 3544
rect 77576 3460 77628 3466
rect 77576 3402 77628 3408
rect 77392 3256 77444 3262
rect 77392 3198 77444 3204
rect 77208 3052 77260 3058
rect 77208 2994 77260 3000
rect 77772 2990 77800 6038
rect 78048 4842 78076 499559
rect 77864 4814 78076 4842
rect 77760 2984 77812 2990
rect 77760 2926 77812 2932
rect 76932 2848 76984 2854
rect 76932 2790 76984 2796
rect 77864 480 77892 4814
rect 78140 3194 78168 506631
rect 78232 121718 78260 700674
rect 81900 700596 81952 700602
rect 81900 700538 81952 700544
rect 81440 700460 81492 700466
rect 81440 700402 81492 700408
rect 79968 700392 80020 700398
rect 79968 700334 80020 700340
rect 78588 700324 78640 700330
rect 78588 700266 78640 700272
rect 78496 586560 78548 586566
rect 78496 586502 78548 586508
rect 78312 583840 78364 583846
rect 78312 583782 78364 583788
rect 78220 121712 78272 121718
rect 78220 121654 78272 121660
rect 78324 6594 78352 583782
rect 78404 583772 78456 583778
rect 78404 583714 78456 583720
rect 78312 6588 78364 6594
rect 78312 6530 78364 6536
rect 78416 6390 78444 583714
rect 78508 6526 78536 586502
rect 78600 119066 78628 700266
rect 78678 573608 78734 573617
rect 78678 573543 78734 573552
rect 78692 572762 78720 573543
rect 78680 572756 78732 572762
rect 78680 572698 78732 572704
rect 78678 559464 78734 559473
rect 78678 559399 78734 559408
rect 78692 558958 78720 559399
rect 78680 558952 78732 558958
rect 78680 558894 78732 558900
rect 79980 534721 80008 700334
rect 80704 582956 80756 582962
rect 80704 582898 80756 582904
rect 79966 534712 80022 534721
rect 79966 534647 80022 534656
rect 78678 520840 78734 520849
rect 78678 520775 78734 520784
rect 78692 172258 78720 520775
rect 80716 496806 80744 582898
rect 81346 563000 81402 563009
rect 81346 562935 81402 562944
rect 80704 496800 80756 496806
rect 80704 496742 80756 496748
rect 81162 489016 81218 489025
rect 81162 488951 81218 488960
rect 79874 481944 79930 481953
rect 79874 481879 79930 481888
rect 79690 446856 79746 446865
rect 79690 446791 79746 446800
rect 79414 411496 79470 411505
rect 79414 411431 79470 411440
rect 78770 400888 78826 400897
rect 78770 400823 78826 400832
rect 78784 400246 78812 400823
rect 78772 400240 78824 400246
rect 78772 400182 78824 400188
rect 78770 393816 78826 393825
rect 78770 393751 78826 393760
rect 78784 393378 78812 393751
rect 78772 393372 78824 393378
rect 78772 393314 78824 393320
rect 79138 348120 79194 348129
rect 79138 348055 79194 348064
rect 79046 253192 79102 253201
rect 79046 253127 79102 253136
rect 78954 231976 79010 231985
rect 78954 231911 79010 231920
rect 78862 196616 78918 196625
rect 78862 196551 78918 196560
rect 78772 188420 78824 188426
rect 78772 188362 78824 188368
rect 78784 184657 78812 188362
rect 78770 184648 78826 184657
rect 78770 184583 78826 184592
rect 78772 183524 78824 183530
rect 78772 183466 78824 183472
rect 78784 182753 78812 183466
rect 78770 182744 78826 182753
rect 78770 182679 78826 182688
rect 78692 172230 78812 172258
rect 78678 172136 78734 172145
rect 78678 172071 78734 172080
rect 78692 171154 78720 172071
rect 78680 171148 78732 171154
rect 78680 171090 78732 171096
rect 78678 168600 78734 168609
rect 78678 168535 78734 168544
rect 78692 168434 78720 168535
rect 78680 168428 78732 168434
rect 78680 168370 78732 168376
rect 78678 165064 78734 165073
rect 78678 164999 78734 165008
rect 78692 164286 78720 164999
rect 78680 164280 78732 164286
rect 78680 164222 78732 164228
rect 78784 162858 78812 172230
rect 78772 162852 78824 162858
rect 78772 162794 78824 162800
rect 78678 161528 78734 161537
rect 78678 161463 78734 161472
rect 78588 119060 78640 119066
rect 78588 119002 78640 119008
rect 78692 13394 78720 161463
rect 78772 157344 78824 157350
rect 78772 157286 78824 157292
rect 78784 151026 78812 157286
rect 78772 151020 78824 151026
rect 78772 150962 78824 150968
rect 78770 150920 78826 150929
rect 78770 150855 78826 150864
rect 78784 150482 78812 150855
rect 78772 150476 78824 150482
rect 78772 150418 78824 150424
rect 78772 150340 78824 150346
rect 78772 150282 78824 150288
rect 78784 147694 78812 150282
rect 78772 147688 78824 147694
rect 78772 147630 78824 147636
rect 78772 135720 78824 135726
rect 78772 135662 78824 135668
rect 78784 133346 78812 135662
rect 78772 133340 78824 133346
rect 78772 133282 78824 133288
rect 78770 133240 78826 133249
rect 78770 133175 78826 133184
rect 78784 122126 78812 133175
rect 78772 122120 78824 122126
rect 78772 122062 78824 122068
rect 78876 121786 78904 196551
rect 78864 121780 78916 121786
rect 78864 121722 78916 121728
rect 78968 118250 78996 231911
rect 79060 120698 79088 253127
rect 79152 203017 79180 348055
rect 79324 296132 79376 296138
rect 79324 296074 79376 296080
rect 79336 287366 79364 296074
rect 79324 287360 79376 287366
rect 79324 287302 79376 287308
rect 79322 274136 79378 274145
rect 79322 274071 79378 274080
rect 79230 259992 79286 260001
rect 79230 259927 79286 259936
rect 79138 203008 79194 203017
rect 79138 202943 79194 202952
rect 79140 202156 79192 202162
rect 79140 202098 79192 202104
rect 79048 120692 79100 120698
rect 79048 120634 79100 120640
rect 78956 118244 79008 118250
rect 78956 118186 79008 118192
rect 79152 116618 79180 202098
rect 79140 116612 79192 116618
rect 79140 116554 79192 116560
rect 79244 113830 79272 259927
rect 79232 113824 79284 113830
rect 79232 113766 79284 113772
rect 79336 111110 79364 274071
rect 79428 264654 79456 411431
rect 79600 328024 79652 328030
rect 79600 327966 79652 327972
rect 79612 319122 79640 327966
rect 79600 319116 79652 319122
rect 79600 319058 79652 319064
rect 79506 284744 79562 284753
rect 79506 284679 79562 284688
rect 79416 264648 79468 264654
rect 79416 264590 79468 264596
rect 79416 237516 79468 237522
rect 79416 237458 79468 237464
rect 79428 225690 79456 237458
rect 79416 225684 79468 225690
rect 79416 225626 79468 225632
rect 79414 210760 79470 210769
rect 79414 210695 79470 210704
rect 79324 111104 79376 111110
rect 79324 111046 79376 111052
rect 79324 91044 79376 91050
rect 79324 90986 79376 90992
rect 79336 81938 79364 90986
rect 79324 81932 79376 81938
rect 79324 81874 79376 81880
rect 79428 14482 79456 210695
rect 79416 14476 79468 14482
rect 79416 14418 79468 14424
rect 78680 13388 78732 13394
rect 78680 13330 78732 13336
rect 79520 10402 79548 284679
rect 79600 280832 79652 280838
rect 79600 280774 79652 280780
rect 79612 272202 79640 280774
rect 79600 272196 79652 272202
rect 79600 272138 79652 272144
rect 79600 260500 79652 260506
rect 79600 260442 79652 260448
rect 79612 252618 79640 260442
rect 79600 252612 79652 252618
rect 79600 252554 79652 252560
rect 79600 225684 79652 225690
rect 79600 225626 79652 225632
rect 79612 215286 79640 225626
rect 79600 215280 79652 215286
rect 79600 215222 79652 215228
rect 79600 205692 79652 205698
rect 79600 205634 79652 205640
rect 79612 196858 79640 205634
rect 79600 196852 79652 196858
rect 79600 196794 79652 196800
rect 79600 185700 79652 185706
rect 79600 185642 79652 185648
rect 79612 176594 79640 185642
rect 79600 176588 79652 176594
rect 79600 176530 79652 176536
rect 79600 167068 79652 167074
rect 79600 167010 79652 167016
rect 79612 157350 79640 167010
rect 79600 157344 79652 157350
rect 79600 157286 79652 157292
rect 79600 147688 79652 147694
rect 79600 147630 79652 147636
rect 79612 135726 79640 147630
rect 79600 135720 79652 135726
rect 79600 135662 79652 135668
rect 79598 130520 79654 130529
rect 79598 130455 79654 130464
rect 79612 123321 79640 130455
rect 79598 123312 79654 123321
rect 79598 123247 79654 123256
rect 79704 121854 79732 446791
rect 79782 351656 79838 351665
rect 79782 351591 79838 351600
rect 79796 287366 79824 351591
rect 79784 287360 79836 287366
rect 79784 287302 79836 287308
rect 79784 280832 79836 280838
rect 79784 280774 79836 280780
rect 79692 121848 79744 121854
rect 79692 121790 79744 121796
rect 79692 121508 79744 121514
rect 79692 121450 79744 121456
rect 79704 99346 79732 121450
rect 79692 99340 79744 99346
rect 79692 99282 79744 99288
rect 79692 69828 79744 69834
rect 79692 69770 79744 69776
rect 79704 56642 79732 69770
rect 79600 56636 79652 56642
rect 79600 56578 79652 56584
rect 79692 56636 79744 56642
rect 79692 56578 79744 56584
rect 79612 53446 79640 56578
rect 79600 53440 79652 53446
rect 79600 53382 79652 53388
rect 79796 10470 79824 280774
rect 79888 127906 79916 481879
rect 80978 471336 81034 471345
rect 80978 471271 81034 471280
rect 80886 460728 80942 460737
rect 80886 460663 80942 460672
rect 80794 443320 80850 443329
rect 80794 443255 80850 443264
rect 80702 439784 80758 439793
rect 80702 439719 80758 439728
rect 80610 404424 80666 404433
rect 80610 404359 80666 404368
rect 79966 337512 80022 337521
rect 79966 337447 80022 337456
rect 79980 328030 80008 337447
rect 79968 328024 80020 328030
rect 79968 327966 80020 327972
rect 80518 316568 80574 316577
rect 80518 316503 80574 316512
rect 79968 272196 80020 272202
rect 79968 272138 80020 272144
rect 79980 260506 80008 272138
rect 80060 264648 80112 264654
rect 80060 264590 80112 264596
rect 79968 260500 80020 260506
rect 79968 260442 80020 260448
rect 79968 252612 80020 252618
rect 79968 252554 80020 252560
rect 79980 237522 80008 252554
rect 79968 237516 80020 237522
rect 79968 237458 80020 237464
rect 79968 215280 80020 215286
rect 79968 215222 80020 215228
rect 79980 205698 80008 215222
rect 79968 205692 80020 205698
rect 79968 205634 80020 205640
rect 79968 196852 80020 196858
rect 79968 196794 80020 196800
rect 79980 185706 80008 196794
rect 79968 185700 80020 185706
rect 79968 185642 80020 185648
rect 79968 176656 80020 176662
rect 79968 176598 80020 176604
rect 79980 175681 80008 176598
rect 79966 175672 80022 175681
rect 79966 175607 80022 175616
rect 79968 175568 80020 175574
rect 79968 175510 80020 175516
rect 79980 167074 80008 175510
rect 79968 167068 80020 167074
rect 79968 167010 80020 167016
rect 79966 154456 80022 154465
rect 79966 154391 80022 154400
rect 79876 127900 79928 127906
rect 79876 127842 79928 127848
rect 79874 126168 79930 126177
rect 79874 126103 79930 126112
rect 79888 13190 79916 126103
rect 79980 123185 80008 154391
rect 79966 123176 80022 123185
rect 79966 123111 80022 123120
rect 80072 111790 80100 264590
rect 80426 241496 80482 241505
rect 80426 241431 80482 241440
rect 80440 239465 80468 241431
rect 80426 239456 80482 239465
rect 80426 239391 80482 239400
rect 80334 237008 80390 237017
rect 80334 236943 80390 236952
rect 80348 236201 80376 236943
rect 80334 236192 80390 236201
rect 80334 236127 80390 236136
rect 80334 217832 80390 217841
rect 80334 217767 80390 217776
rect 80348 216714 80376 217767
rect 80336 216708 80388 216714
rect 80336 216650 80388 216656
rect 80150 209128 80206 209137
rect 80150 209063 80206 209072
rect 80164 202745 80192 209063
rect 80242 207768 80298 207777
rect 80242 207703 80298 207712
rect 80150 202736 80206 202745
rect 80150 202671 80206 202680
rect 80150 202056 80206 202065
rect 80150 201991 80206 202000
rect 80164 199617 80192 201991
rect 80256 201657 80284 207703
rect 80334 203688 80390 203697
rect 80334 203623 80390 203632
rect 80348 202162 80376 203623
rect 80426 203008 80482 203017
rect 80426 202943 80482 202952
rect 80336 202156 80388 202162
rect 80336 202098 80388 202104
rect 80242 201648 80298 201657
rect 80242 201583 80298 201592
rect 80336 200252 80388 200258
rect 80336 200194 80388 200200
rect 80150 199608 80206 199617
rect 80150 199543 80206 199552
rect 80244 191140 80296 191146
rect 80244 191082 80296 191088
rect 80150 190360 80206 190369
rect 80150 190295 80206 190304
rect 80164 178401 80192 190295
rect 80256 180033 80284 191082
rect 80348 188465 80376 200194
rect 80334 188456 80390 188465
rect 80334 188391 80390 188400
rect 80334 186280 80390 186289
rect 80334 186215 80390 186224
rect 80242 180024 80298 180033
rect 80242 179959 80298 179968
rect 80242 179888 80298 179897
rect 80242 179823 80298 179832
rect 80150 178392 80206 178401
rect 80150 178327 80206 178336
rect 80150 171456 80206 171465
rect 80150 171391 80206 171400
rect 80164 165617 80192 171391
rect 80256 171193 80284 179823
rect 80242 171184 80298 171193
rect 80242 171119 80298 171128
rect 80150 165608 80206 165617
rect 80150 165543 80206 165552
rect 80150 149696 80206 149705
rect 80150 149631 80206 149640
rect 80164 143177 80192 149631
rect 80242 144120 80298 144129
rect 80242 144055 80244 144064
rect 80296 144055 80298 144064
rect 80244 144026 80296 144032
rect 80242 143848 80298 143857
rect 80242 143783 80298 143792
rect 80150 143168 80206 143177
rect 80150 143103 80206 143112
rect 80150 141944 80206 141953
rect 80150 141879 80206 141888
rect 80164 140418 80192 141879
rect 80152 140412 80204 140418
rect 80152 140354 80204 140360
rect 80150 140312 80206 140321
rect 80150 140247 80206 140256
rect 80164 123457 80192 140247
rect 80150 123448 80206 123457
rect 80150 123383 80206 123392
rect 80060 111784 80112 111790
rect 80060 111726 80112 111732
rect 80060 102196 80112 102202
rect 80060 102138 80112 102144
rect 79968 99340 80020 99346
rect 79968 99282 80020 99288
rect 79980 91050 80008 99282
rect 79968 91044 80020 91050
rect 79968 90986 80020 90992
rect 80072 82822 80100 102138
rect 80256 83502 80284 143783
rect 80348 115258 80376 186215
rect 80440 137329 80468 202943
rect 80426 137320 80482 137329
rect 80426 137255 80482 137264
rect 80428 137216 80480 137222
rect 80426 137184 80428 137193
rect 80480 137184 80482 137193
rect 80426 137119 80482 137128
rect 80428 137080 80480 137086
rect 80428 137022 80480 137028
rect 80440 136921 80468 137022
rect 80426 136912 80482 136921
rect 80426 136847 80482 136856
rect 80426 136776 80482 136785
rect 80426 136711 80482 136720
rect 80440 135969 80468 136711
rect 80426 135960 80482 135969
rect 80426 135895 80482 135904
rect 80428 127900 80480 127906
rect 80428 127842 80480 127848
rect 80336 115252 80388 115258
rect 80336 115194 80388 115200
rect 80244 83496 80296 83502
rect 80244 83438 80296 83444
rect 80060 82816 80112 82822
rect 80060 82758 80112 82764
rect 79968 81932 80020 81938
rect 79968 81874 80020 81880
rect 79980 69834 80008 81874
rect 80152 73228 80204 73234
rect 80152 73170 80204 73176
rect 79968 69828 80020 69834
rect 79968 69770 80020 69776
rect 80164 66298 80192 73170
rect 80060 66292 80112 66298
rect 80060 66234 80112 66240
rect 80152 66292 80204 66298
rect 80152 66234 80204 66240
rect 79968 53440 80020 53446
rect 79968 53382 80020 53388
rect 79980 44878 80008 53382
rect 79968 44872 80020 44878
rect 79968 44814 80020 44820
rect 79876 13184 79928 13190
rect 79876 13126 79928 13132
rect 79784 10464 79836 10470
rect 79784 10406 79836 10412
rect 79508 10396 79560 10402
rect 79508 10338 79560 10344
rect 80072 6905 80100 66234
rect 80058 6896 80114 6905
rect 80058 6831 80114 6840
rect 80334 6896 80390 6905
rect 80334 6831 80390 6840
rect 78496 6520 78548 6526
rect 78496 6462 78548 6468
rect 78404 6384 78456 6390
rect 78404 6326 78456 6332
rect 79046 3768 79102 3777
rect 79046 3703 79102 3712
rect 78128 3188 78180 3194
rect 78128 3130 78180 3136
rect 79060 480 79088 3703
rect 80348 610 80376 6831
rect 80440 3874 80468 127842
rect 80532 118318 80560 316503
rect 80624 119610 80652 404359
rect 80716 122262 80744 439719
rect 80808 122330 80836 443255
rect 80796 122324 80848 122330
rect 80796 122266 80848 122272
rect 80704 122256 80756 122262
rect 80704 122198 80756 122204
rect 80900 122058 80928 460663
rect 80992 136882 81020 471271
rect 81070 464264 81126 464273
rect 81070 464199 81126 464208
rect 80980 136876 81032 136882
rect 80980 136818 81032 136824
rect 80978 136776 81034 136785
rect 80978 136711 81034 136720
rect 80992 136678 81020 136711
rect 80980 136672 81032 136678
rect 80980 136614 81032 136620
rect 80980 136536 81032 136542
rect 80980 136478 81032 136484
rect 80888 122052 80940 122058
rect 80888 121994 80940 122000
rect 80992 120562 81020 136478
rect 80980 120556 81032 120562
rect 80980 120498 81032 120504
rect 80612 119604 80664 119610
rect 80612 119546 80664 119552
rect 80520 118312 80572 118318
rect 80520 118254 80572 118260
rect 81084 111178 81112 464199
rect 81176 122670 81204 488951
rect 81254 425640 81310 425649
rect 81254 425575 81310 425584
rect 81164 122664 81216 122670
rect 81164 122606 81216 122612
rect 81072 111172 81124 111178
rect 81072 111114 81124 111120
rect 81268 14550 81296 425575
rect 81360 122602 81388 562935
rect 81452 239057 81480 700402
rect 81532 673532 81584 673538
rect 81532 673474 81584 673480
rect 81438 239048 81494 239057
rect 81438 238983 81494 238992
rect 81438 233744 81494 233753
rect 81438 233679 81440 233688
rect 81492 233679 81494 233688
rect 81440 233650 81492 233656
rect 81440 230648 81492 230654
rect 81440 230590 81492 230596
rect 81452 229537 81480 230590
rect 81438 229528 81494 229537
rect 81438 229463 81494 229472
rect 81440 229288 81492 229294
rect 81438 229256 81440 229265
rect 81492 229256 81494 229265
rect 81438 229191 81494 229200
rect 81440 227928 81492 227934
rect 81438 227896 81440 227905
rect 81492 227896 81494 227905
rect 81438 227831 81494 227840
rect 81438 223408 81494 223417
rect 81438 223343 81494 223352
rect 81452 208049 81480 223343
rect 81544 221377 81572 673474
rect 81622 566536 81678 566545
rect 81622 566471 81678 566480
rect 81530 221368 81586 221377
rect 81530 221303 81586 221312
rect 81530 214296 81586 214305
rect 81530 214231 81586 214240
rect 81544 213450 81572 214231
rect 81532 213444 81584 213450
rect 81532 213386 81584 213392
rect 81530 210488 81586 210497
rect 81530 210423 81586 210432
rect 81438 208040 81494 208049
rect 81438 207975 81494 207984
rect 81544 207754 81572 210423
rect 81452 207726 81572 207754
rect 81452 200258 81480 207726
rect 81530 207224 81586 207233
rect 81530 207159 81586 207168
rect 81544 202502 81572 207159
rect 81532 202496 81584 202502
rect 81532 202438 81584 202444
rect 81530 201920 81586 201929
rect 81530 201855 81586 201864
rect 81544 201822 81572 201855
rect 81532 201816 81584 201822
rect 81532 201758 81584 201764
rect 81532 201272 81584 201278
rect 81530 201240 81532 201249
rect 81584 201240 81586 201249
rect 81530 201175 81586 201184
rect 81530 201104 81586 201113
rect 81530 201039 81586 201048
rect 81544 200326 81572 201039
rect 81532 200320 81584 200326
rect 81532 200262 81584 200268
rect 81440 200252 81492 200258
rect 81440 200194 81492 200200
rect 81532 200184 81584 200190
rect 81438 200152 81494 200161
rect 81532 200126 81584 200132
rect 81438 200087 81494 200096
rect 81348 122596 81400 122602
rect 81348 122538 81400 122544
rect 81256 14544 81308 14550
rect 81256 14486 81308 14492
rect 81452 9178 81480 200087
rect 81544 192438 81572 200126
rect 81532 192432 81584 192438
rect 81532 192374 81584 192380
rect 81530 192264 81586 192273
rect 81530 192199 81532 192208
rect 81584 192199 81586 192208
rect 81532 192170 81584 192176
rect 81530 191856 81586 191865
rect 81530 191791 81532 191800
rect 81584 191791 81586 191800
rect 81532 191762 81584 191768
rect 81532 190732 81584 190738
rect 81532 190674 81584 190680
rect 81544 170785 81572 190674
rect 81530 170776 81586 170785
rect 81530 170711 81586 170720
rect 81530 162208 81586 162217
rect 81530 162143 81532 162152
rect 81584 162143 81586 162152
rect 81532 162114 81584 162120
rect 81530 160848 81586 160857
rect 81530 160783 81586 160792
rect 81544 157486 81572 160783
rect 81532 157480 81584 157486
rect 81532 157422 81584 157428
rect 81532 157344 81584 157350
rect 81530 157312 81532 157321
rect 81584 157312 81586 157321
rect 81530 157247 81586 157256
rect 81532 157208 81584 157214
rect 81532 157150 81584 157156
rect 81544 144129 81572 157150
rect 81530 144120 81586 144129
rect 81530 144055 81586 144064
rect 81530 143984 81586 143993
rect 81530 143919 81586 143928
rect 81440 9172 81492 9178
rect 81440 9114 81492 9120
rect 81544 7546 81572 143919
rect 81636 118590 81664 566471
rect 81806 517304 81862 517313
rect 81806 517239 81862 517248
rect 81714 415032 81770 415041
rect 81714 414967 81770 414976
rect 81624 118584 81676 118590
rect 81624 118526 81676 118532
rect 81728 9382 81756 414967
rect 81820 118454 81848 517239
rect 81912 327457 81940 700538
rect 89180 699825 89208 703520
rect 105464 700330 105492 703520
rect 137848 700670 137876 703520
rect 154132 700777 154160 703520
rect 154118 700768 154174 700777
rect 154118 700703 154174 700712
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 170324 700602 170352 703520
rect 202800 700602 202828 703520
rect 218992 700641 219020 703520
rect 235184 700738 235212 703520
rect 235172 700732 235224 700738
rect 235172 700674 235224 700680
rect 218978 700632 219034 700641
rect 170312 700596 170364 700602
rect 170312 700538 170364 700544
rect 202788 700596 202840 700602
rect 218978 700567 219034 700576
rect 202788 700538 202840 700544
rect 267660 700505 267688 703520
rect 283852 700806 283880 703520
rect 283840 700800 283892 700806
rect 283840 700742 283892 700748
rect 300136 700738 300164 703520
rect 332520 700738 332548 703520
rect 335268 700868 335320 700874
rect 335268 700810 335320 700816
rect 269028 700732 269080 700738
rect 269028 700674 269080 700680
rect 300124 700732 300176 700738
rect 300124 700674 300176 700680
rect 332508 700732 332560 700738
rect 332508 700674 332560 700680
rect 267646 700496 267702 700505
rect 267646 700431 267702 700440
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 142068 700324 142120 700330
rect 142068 700266 142120 700272
rect 89166 699816 89222 699825
rect 89166 699751 89222 699760
rect 89534 695464 89590 695473
rect 89534 695399 89590 695408
rect 89548 689353 89576 695399
rect 89534 689344 89590 689353
rect 89534 689279 89590 689288
rect 89534 674792 89590 674801
rect 89534 674727 89590 674736
rect 89548 665281 89576 674727
rect 89534 665272 89590 665281
rect 89534 665207 89590 665216
rect 89534 655480 89590 655489
rect 89534 655415 89590 655424
rect 89548 645969 89576 655415
rect 89534 645960 89590 645969
rect 89534 645895 89590 645904
rect 89534 636168 89590 636177
rect 89534 636103 89590 636112
rect 89548 626657 89576 636103
rect 89534 626648 89590 626657
rect 82084 626612 82136 626618
rect 89534 626583 89590 626592
rect 82084 626554 82136 626560
rect 81990 467256 82046 467265
rect 81990 467191 82046 467200
rect 81898 327448 81954 327457
rect 81898 327383 81954 327392
rect 81898 291272 81954 291281
rect 81898 291207 81954 291216
rect 81808 118448 81860 118454
rect 81808 118390 81860 118396
rect 81716 9376 81768 9382
rect 81716 9318 81768 9324
rect 81532 7540 81584 7546
rect 81532 7482 81584 7488
rect 81912 4826 81940 291207
rect 82004 123554 82032 467191
rect 82096 391105 82124 626554
rect 83556 603152 83608 603158
rect 83556 603094 83608 603100
rect 83568 597553 83596 603094
rect 83554 597544 83610 597553
rect 83554 597479 83610 597488
rect 83738 597544 83794 597553
rect 83738 597479 83794 597488
rect 83752 590782 83780 597479
rect 89442 596184 89498 596193
rect 89442 596119 89498 596128
rect 89456 593366 89484 596119
rect 89352 593360 89404 593366
rect 89352 593302 89404 593308
rect 89444 593360 89496 593366
rect 89444 593302 89496 593308
rect 83556 590776 83608 590782
rect 83556 590718 83608 590724
rect 83740 590776 83792 590782
rect 83740 590718 83792 590724
rect 83568 586498 83596 590718
rect 83556 586492 83608 586498
rect 83556 586434 83608 586440
rect 83648 586424 83700 586430
rect 83648 586366 83700 586372
rect 82636 581324 82688 581330
rect 82636 581266 82688 581272
rect 82648 577697 82676 581266
rect 82634 577688 82690 577697
rect 82634 577623 82690 577632
rect 83660 574818 83688 586366
rect 89364 582865 89392 593302
rect 90916 585064 90968 585070
rect 90916 585006 90968 585012
rect 89350 582856 89406 582865
rect 89350 582791 89406 582800
rect 86316 582616 86368 582622
rect 86316 582558 86368 582564
rect 85212 582004 85264 582010
rect 85212 581946 85264 581952
rect 85224 581505 85252 581946
rect 85488 581800 85540 581806
rect 86328 581777 86356 582558
rect 90456 582344 90508 582350
rect 89074 582312 89130 582321
rect 90456 582286 90508 582292
rect 89074 582247 89130 582256
rect 85488 581742 85540 581748
rect 86314 581768 86370 581777
rect 85500 581505 85528 581742
rect 86314 581703 86370 581712
rect 89088 581641 89116 582247
rect 89720 582072 89772 582078
rect 89718 582040 89720 582049
rect 89772 582040 89774 582049
rect 89718 581975 89774 581984
rect 89810 581904 89866 581913
rect 89810 581839 89866 581848
rect 89824 581641 89852 581839
rect 89074 581632 89130 581641
rect 89074 581567 89130 581576
rect 89810 581632 89866 581641
rect 89810 581567 89866 581576
rect 85210 581496 85266 581505
rect 85210 581431 85266 581440
rect 85486 581496 85542 581505
rect 85486 581431 85542 581440
rect 90468 581369 90496 582286
rect 90928 581369 90956 585006
rect 92112 584860 92164 584866
rect 92112 584802 92164 584808
rect 92124 583817 92152 584802
rect 105360 584792 105412 584798
rect 105360 584734 105412 584740
rect 103520 584724 103572 584730
rect 103520 584666 103572 584672
rect 96344 584044 96396 584050
rect 96344 583986 96396 583992
rect 92110 583808 92166 583817
rect 92110 583743 92166 583752
rect 94226 582448 94282 582457
rect 93780 582406 94176 582434
rect 93674 582312 93730 582321
rect 93674 582247 93730 582256
rect 93216 582208 93268 582214
rect 93216 582150 93268 582156
rect 91928 582072 91980 582078
rect 91928 582014 91980 582020
rect 92664 582072 92716 582078
rect 92664 582014 92716 582020
rect 91940 581913 91968 582014
rect 91926 581904 91982 581913
rect 91926 581839 91982 581848
rect 92676 581369 92704 582014
rect 93228 581369 93256 582150
rect 93398 582040 93454 582049
rect 93688 582026 93716 582247
rect 93780 582185 93808 582406
rect 94148 582321 94176 582406
rect 94226 582383 94282 582392
rect 94134 582312 94190 582321
rect 93952 582276 94004 582282
rect 94134 582247 94190 582256
rect 93952 582218 94004 582224
rect 93766 582176 93822 582185
rect 93766 582111 93822 582120
rect 93688 581998 93808 582026
rect 93398 581975 93454 581984
rect 93412 581369 93440 581975
rect 93780 581505 93808 581998
rect 93964 581876 93992 582218
rect 94240 581777 94268 582383
rect 96356 581876 96384 583986
rect 96528 582616 96580 582622
rect 96528 582558 96580 582564
rect 96620 582616 96672 582622
rect 96620 582558 96672 582564
rect 101312 582616 101364 582622
rect 101312 582558 101364 582564
rect 96540 582026 96568 582558
rect 96632 582026 96660 582558
rect 101324 582457 101352 582558
rect 101310 582448 101366 582457
rect 101310 582383 101366 582392
rect 99840 582344 99892 582350
rect 99840 582286 99892 582292
rect 101586 582312 101642 582321
rect 96540 581998 96660 582026
rect 94226 581768 94282 581777
rect 94226 581703 94282 581712
rect 96894 581768 96950 581777
rect 96894 581703 96950 581712
rect 93766 581496 93822 581505
rect 93766 581431 93822 581440
rect 96908 581369 96936 581703
rect 99852 581505 99880 582286
rect 100024 582276 100076 582282
rect 101586 582247 101642 582256
rect 100024 582218 100076 582224
rect 99470 581496 99526 581505
rect 99470 581431 99526 581440
rect 99838 581496 99894 581505
rect 99838 581431 99894 581440
rect 99484 581398 99512 581431
rect 98460 581392 98512 581398
rect 84934 581360 84990 581369
rect 84594 581318 84934 581346
rect 84934 581295 84990 581304
rect 89258 581360 89314 581369
rect 90454 581360 90510 581369
rect 89314 581318 89378 581346
rect 89258 581295 89314 581304
rect 90454 581295 90510 581304
rect 90914 581360 90970 581369
rect 91742 581360 91798 581369
rect 91586 581318 91742 581346
rect 90914 581295 90970 581304
rect 91742 581295 91798 581304
rect 92662 581360 92718 581369
rect 92662 581295 92718 581304
rect 93214 581360 93270 581369
rect 93214 581295 93270 581304
rect 93398 581360 93454 581369
rect 93398 581295 93454 581304
rect 96894 581360 96950 581369
rect 99472 581392 99524 581398
rect 98512 581340 98762 581346
rect 98460 581334 98762 581340
rect 100036 581369 100064 582218
rect 101600 581890 101628 582247
rect 101154 581862 101628 581890
rect 103532 581876 103560 584666
rect 105372 582282 105400 584734
rect 117872 584724 117924 584730
rect 117872 584666 117924 584672
rect 105912 583840 105964 583846
rect 105912 583782 105964 583788
rect 107660 583840 107712 583846
rect 107660 583782 107712 583788
rect 105360 582276 105412 582282
rect 105360 582218 105412 582224
rect 105924 581876 105952 583782
rect 107672 582457 107700 583782
rect 113088 583772 113140 583778
rect 113088 583714 113140 583720
rect 110696 582820 110748 582826
rect 110696 582762 110748 582768
rect 107658 582448 107714 582457
rect 107658 582383 107714 582392
rect 110708 581876 110736 582762
rect 111064 582344 111116 582350
rect 111064 582286 111116 582292
rect 111076 581641 111104 582286
rect 113100 581876 113128 583714
rect 115848 582616 115900 582622
rect 115848 582558 115900 582564
rect 113270 582448 113326 582457
rect 113270 582383 113326 582392
rect 111062 581632 111118 581641
rect 111062 581567 111118 581576
rect 113284 581505 113312 582383
rect 113270 581496 113326 581505
rect 113270 581431 113326 581440
rect 103428 581392 103480 581398
rect 99472 581334 99524 581340
rect 100022 581360 100078 581369
rect 98472 581318 98762 581334
rect 96894 581295 96950 581304
rect 100022 581295 100078 581304
rect 103426 581360 103428 581369
rect 108672 581392 108724 581398
rect 103480 581360 103482 581369
rect 108330 581340 108672 581346
rect 115860 581369 115888 582558
rect 117884 581876 117912 584666
rect 131948 584112 132000 584118
rect 131948 584054 132000 584060
rect 127440 583976 127492 583982
rect 127440 583918 127492 583924
rect 125048 583840 125100 583846
rect 125048 583782 125100 583788
rect 123482 582312 123538 582321
rect 118700 582276 118752 582282
rect 123482 582247 123538 582256
rect 123758 582312 123814 582321
rect 123758 582247 123760 582256
rect 118700 582218 118752 582224
rect 118606 582040 118662 582049
rect 118528 581998 118606 582026
rect 118528 581641 118556 581998
rect 118606 581975 118662 581984
rect 118514 581632 118570 581641
rect 118514 581567 118570 581576
rect 118712 581369 118740 582218
rect 122656 582208 122708 582214
rect 122656 582150 122708 582156
rect 122668 581876 122696 582150
rect 120080 581664 120132 581670
rect 120132 581612 120290 581618
rect 120080 581606 120290 581612
rect 120092 581590 120290 581606
rect 123496 581505 123524 582247
rect 123812 582247 123814 582256
rect 123760 582218 123812 582224
rect 125060 581876 125088 583782
rect 127452 581876 127480 583918
rect 131960 583438 131988 584054
rect 142080 584050 142108 700266
rect 190368 650072 190420 650078
rect 190368 650014 190420 650020
rect 190380 585138 190408 650014
rect 236920 586560 236972 586566
rect 236920 586502 236972 586508
rect 163136 585132 163188 585138
rect 163136 585074 163188 585080
rect 189264 585132 189316 585138
rect 189264 585074 189316 585080
rect 190368 585132 190420 585138
rect 190368 585074 190420 585080
rect 197084 585132 197136 585138
rect 197084 585074 197136 585080
rect 148782 584896 148838 584905
rect 148782 584831 148838 584840
rect 157246 584896 157302 584905
rect 157430 584896 157486 584905
rect 157302 584854 157430 584882
rect 157246 584831 157302 584840
rect 157430 584831 157486 584840
rect 136824 584044 136876 584050
rect 136824 583986 136876 583992
rect 141608 584044 141660 584050
rect 141608 583986 141660 583992
rect 142068 584044 142120 584050
rect 142068 583986 142120 583992
rect 131948 583432 132000 583438
rect 131948 583374 132000 583380
rect 129832 582684 129884 582690
rect 129832 582626 129884 582632
rect 132224 582684 132276 582690
rect 132224 582626 132276 582632
rect 128360 582208 128412 582214
rect 128360 582150 128412 582156
rect 128372 582049 128400 582150
rect 128358 582040 128414 582049
rect 128358 581975 128414 581984
rect 129844 581876 129872 582626
rect 132236 581876 132264 582626
rect 132498 582448 132554 582457
rect 132498 582383 132554 582392
rect 123482 581496 123538 581505
rect 132512 581482 132540 582383
rect 132958 582312 133014 582321
rect 132958 582247 133014 582256
rect 132972 581505 133000 582247
rect 136836 581876 136864 583986
rect 139214 583808 139270 583817
rect 139214 583743 139270 583752
rect 137928 582208 137980 582214
rect 137928 582150 137980 582156
rect 137940 582049 137968 582150
rect 137926 582040 137982 582049
rect 137926 581975 137982 581984
rect 139228 581876 139256 583743
rect 141620 581876 141648 583986
rect 146392 582752 146444 582758
rect 146392 582694 146444 582700
rect 142802 582312 142858 582321
rect 142802 582247 142858 582256
rect 134340 581664 134392 581670
rect 134392 581612 134642 581618
rect 134340 581606 134642 581612
rect 134352 581590 134642 581606
rect 142816 581505 142844 582247
rect 146404 581876 146432 582694
rect 147678 582312 147734 582321
rect 147678 582247 147734 582256
rect 146944 582208 146996 582214
rect 146944 582150 146996 582156
rect 144368 581664 144420 581670
rect 144026 581612 144368 581618
rect 144026 581606 144420 581612
rect 144026 581590 144408 581606
rect 132590 581496 132646 581505
rect 132512 581454 132590 581482
rect 123482 581431 123538 581440
rect 132590 581431 132646 581440
rect 132958 581496 133014 581505
rect 132958 581431 133014 581440
rect 142802 581496 142858 581505
rect 142802 581431 142858 581440
rect 146956 581369 146984 582150
rect 147692 582049 147720 582247
rect 147678 582040 147734 582049
rect 147678 581975 147734 581984
rect 148796 581876 148824 584831
rect 158350 584760 158406 584769
rect 158350 584695 158406 584704
rect 156326 582448 156382 582457
rect 156326 582383 156382 582392
rect 150990 582312 151046 582321
rect 150990 582247 150992 582256
rect 151044 582247 151046 582256
rect 151174 582312 151230 582321
rect 151174 582247 151230 582256
rect 150992 582218 151044 582224
rect 151188 581876 151216 582247
rect 156340 582049 156368 582383
rect 156602 582312 156658 582321
rect 156602 582247 156658 582256
rect 157156 582276 157208 582282
rect 155866 582040 155922 582049
rect 155866 581975 155922 581984
rect 156326 582040 156382 582049
rect 156326 581975 156382 581984
rect 155880 581890 155908 581975
rect 155880 581862 155986 581890
rect 156616 581641 156644 582247
rect 157156 582218 157208 582224
rect 157248 582276 157300 582282
rect 157248 582218 157300 582224
rect 157168 582049 157196 582218
rect 157154 582040 157210 582049
rect 157154 581975 157210 581984
rect 157064 581664 157116 581670
rect 147862 581632 147918 581641
rect 153934 581632 153990 581641
rect 153594 581590 153934 581618
rect 147862 581567 147918 581576
rect 153934 581567 153990 581576
rect 156602 581632 156658 581641
rect 157064 581606 157116 581612
rect 156602 581567 156658 581576
rect 147876 581369 147904 581567
rect 157076 581505 157104 581606
rect 157062 581496 157118 581505
rect 157062 581431 157118 581440
rect 157260 581369 157288 582218
rect 158364 581876 158392 584695
rect 162490 582312 162546 582321
rect 162490 582247 162492 582256
rect 162544 582247 162546 582256
rect 162492 582218 162544 582224
rect 160468 582208 160520 582214
rect 160468 582150 160520 582156
rect 160480 581890 160508 582150
rect 160480 581862 160770 581890
rect 163148 581876 163176 585074
rect 167920 584860 167972 584866
rect 167920 584802 167972 584808
rect 182272 584860 182324 584866
rect 182272 584802 182324 584808
rect 166814 582312 166870 582321
rect 166998 582312 167054 582321
rect 166870 582270 166948 582298
rect 166814 582247 166870 582256
rect 157524 581664 157576 581670
rect 157524 581606 157576 581612
rect 157536 581505 157564 581606
rect 165252 581528 165304 581534
rect 157522 581496 157578 581505
rect 165304 581476 165554 581482
rect 165252 581470 165554 581476
rect 165264 581454 165554 581470
rect 157522 581431 157578 581440
rect 166920 581369 166948 582270
rect 166998 582247 167054 582256
rect 167012 581641 167040 582247
rect 167092 582208 167144 582214
rect 167092 582150 167144 582156
rect 167104 582049 167132 582150
rect 167090 582040 167146 582049
rect 167090 581975 167146 581984
rect 167932 581876 167960 584802
rect 182178 584760 182234 584769
rect 182178 584695 182234 584704
rect 182192 584610 182220 584695
rect 182284 584610 182312 584802
rect 182192 584582 182312 584610
rect 182270 584488 182326 584497
rect 182270 584423 182326 584432
rect 175094 584352 175150 584361
rect 175094 584287 175150 584296
rect 170312 584044 170364 584050
rect 170312 583986 170364 583992
rect 170324 581876 170352 583986
rect 171598 582312 171654 582321
rect 171598 582247 171654 582256
rect 171782 582312 171838 582321
rect 171782 582247 171838 582256
rect 166998 581632 167054 581641
rect 166998 581567 167054 581576
rect 108330 581334 108724 581340
rect 108946 581360 109002 581369
rect 108330 581318 108712 581334
rect 103426 581295 103482 581304
rect 109130 581360 109186 581369
rect 109002 581318 109130 581346
rect 108946 581295 109002 581304
rect 109130 581295 109186 581304
rect 115202 581360 115258 581369
rect 115846 581360 115902 581369
rect 115258 581318 115506 581346
rect 115202 581295 115258 581304
rect 115846 581295 115902 581304
rect 118698 581360 118754 581369
rect 118698 581295 118754 581304
rect 146942 581360 146998 581369
rect 146942 581295 146998 581304
rect 147862 581360 147918 581369
rect 147862 581295 147918 581304
rect 157246 581360 157302 581369
rect 157246 581295 157302 581304
rect 166906 581360 166962 581369
rect 171612 581346 171640 582247
rect 171796 581505 171824 582247
rect 175108 581876 175136 584287
rect 179878 583944 179934 583953
rect 179878 583879 179934 583888
rect 177488 582820 177540 582826
rect 177488 582762 177540 582768
rect 176568 582208 176620 582214
rect 176568 582150 176620 582156
rect 176580 582049 176608 582150
rect 176566 582040 176622 582049
rect 176566 581975 176622 581984
rect 177500 581876 177528 582762
rect 179892 581876 179920 583879
rect 181442 582312 181498 582321
rect 181442 582247 181498 582256
rect 172520 581800 172572 581806
rect 172572 581748 172730 581754
rect 172520 581742 172730 581748
rect 172532 581726 172730 581742
rect 176568 581528 176620 581534
rect 171782 581496 171838 581505
rect 171966 581496 172022 581505
rect 171782 581431 171838 581440
rect 171888 581454 171966 581482
rect 171888 581346 171916 581454
rect 176568 581470 176620 581476
rect 176752 581528 176804 581534
rect 181456 581505 181484 582247
rect 182284 581876 182312 584423
rect 186870 583944 186926 583953
rect 186870 583879 186926 583888
rect 184480 582888 184532 582894
rect 184480 582830 184532 582836
rect 184492 581876 184520 582830
rect 186318 582040 186374 582049
rect 186318 581975 186374 581984
rect 186332 581806 186360 581975
rect 186884 581876 186912 583879
rect 189276 581876 189304 585074
rect 191746 584896 191802 584905
rect 191746 584831 191748 584840
rect 191800 584831 191802 584840
rect 191748 584802 191800 584808
rect 197096 583370 197124 585074
rect 205638 585032 205694 585041
rect 205560 584990 205638 585018
rect 205560 584905 205588 584990
rect 205638 584967 205694 584976
rect 225142 585032 225198 585041
rect 225142 584967 225198 584976
rect 227732 584990 227852 585018
rect 205546 584896 205602 584905
rect 205546 584831 205602 584840
rect 218150 584896 218206 584905
rect 218150 584831 218206 584840
rect 215576 584792 215628 584798
rect 215576 584734 215628 584740
rect 218058 584760 218114 584769
rect 210792 584248 210844 584254
rect 210792 584190 210844 584196
rect 201222 584080 201278 584089
rect 201222 584015 201278 584024
rect 197084 583364 197136 583370
rect 197084 583306 197136 583312
rect 198832 582956 198884 582962
rect 198832 582898 198884 582904
rect 196438 582448 196494 582457
rect 196438 582383 196494 582392
rect 190826 582312 190882 582321
rect 190826 582247 190882 582256
rect 186320 581800 186372 581806
rect 186320 581742 186372 581748
rect 190840 581505 190868 582247
rect 191654 582176 191710 582185
rect 191654 582111 191710 582120
rect 192022 582176 192078 582185
rect 192022 582111 192078 582120
rect 191668 581876 191696 582111
rect 176752 581470 176804 581476
rect 181442 581496 181498 581505
rect 171966 581431 172022 581440
rect 176580 581369 176608 581470
rect 176764 581369 176792 581470
rect 181442 581431 181498 581440
rect 190826 581496 190882 581505
rect 190826 581431 190882 581440
rect 192036 581369 192064 582111
rect 195886 582040 195942 582049
rect 195886 581975 195942 581984
rect 192208 581800 192260 581806
rect 192208 581742 192260 581748
rect 192220 581369 192248 581742
rect 194416 581528 194468 581534
rect 194074 581476 194416 581482
rect 194074 581470 194468 581476
rect 194074 581454 194456 581470
rect 195900 581369 195928 581975
rect 196452 581876 196480 582383
rect 198844 581876 198872 582898
rect 200762 582312 200818 582321
rect 200762 582247 200818 582256
rect 200670 582176 200726 582185
rect 200670 582111 200726 582120
rect 198004 581664 198056 581670
rect 198002 581632 198004 581641
rect 198056 581632 198058 581641
rect 198002 581567 198058 581576
rect 200684 581369 200712 582111
rect 200776 581505 200804 582247
rect 200854 582176 200910 582185
rect 200854 582111 200910 582120
rect 200868 581670 200896 582111
rect 201236 581876 201264 584015
rect 206006 582584 206062 582593
rect 206006 582519 206062 582528
rect 203338 582040 203394 582049
rect 203338 581975 203394 581984
rect 203352 581890 203380 581975
rect 203352 581862 203642 581890
rect 206020 581876 206048 582519
rect 210330 582040 210386 582049
rect 210330 581975 210386 581984
rect 208306 581904 208362 581913
rect 208362 581862 208426 581890
rect 208306 581839 208362 581848
rect 200856 581664 200908 581670
rect 200856 581606 200908 581612
rect 200762 581496 200818 581505
rect 200762 581431 200818 581440
rect 210344 581369 210372 581975
rect 210422 581904 210478 581913
rect 210804 581876 210832 584190
rect 213182 582856 213238 582865
rect 213182 582791 213238 582800
rect 211158 582312 211214 582321
rect 211158 582247 211214 582256
rect 210422 581839 210478 581848
rect 210436 581505 210464 581839
rect 210422 581496 210478 581505
rect 210422 581431 210478 581440
rect 211172 581369 211200 582247
rect 213196 581876 213224 582791
rect 215588 581876 215616 584734
rect 218058 584695 218114 584704
rect 217968 584656 218020 584662
rect 218072 584644 218100 584695
rect 218164 584644 218192 584831
rect 218072 584616 218192 584644
rect 217968 584598 218020 584604
rect 217980 581876 218008 584598
rect 222750 584080 222806 584089
rect 222750 584015 222806 584024
rect 220360 582752 220412 582758
rect 220360 582694 220412 582700
rect 220082 581904 220138 581913
rect 220372 581876 220400 582694
rect 220910 582040 220966 582049
rect 220910 581975 220966 581984
rect 220726 581904 220782 581913
rect 220082 581839 220138 581848
rect 220726 581839 220782 581848
rect 220096 581505 220124 581839
rect 220082 581496 220138 581505
rect 220082 581431 220138 581440
rect 220740 581369 220768 581839
rect 220924 581369 220952 581975
rect 222764 581876 222792 584015
rect 225156 581876 225184 584967
rect 227732 584905 227760 584990
rect 227718 584896 227774 584905
rect 227718 584831 227774 584840
rect 226340 584792 226392 584798
rect 226340 584734 226392 584740
rect 226352 582146 226380 584734
rect 227824 584662 227852 584990
rect 234526 584760 234582 584769
rect 233240 584724 233292 584730
rect 234526 584695 234582 584704
rect 233240 584666 233292 584672
rect 227812 584656 227864 584662
rect 227812 584598 227864 584604
rect 233252 584497 233280 584666
rect 234540 584662 234568 584695
rect 234528 584656 234580 584662
rect 234528 584598 234580 584604
rect 233238 584488 233294 584497
rect 233238 584423 233294 584432
rect 234526 583808 234582 583817
rect 234526 583743 234582 583752
rect 229744 582956 229796 582962
rect 229744 582898 229796 582904
rect 229374 582176 229430 582185
rect 226340 582140 226392 582146
rect 229374 582111 229430 582120
rect 226340 582082 226392 582088
rect 227720 581664 227772 581670
rect 227562 581612 227720 581618
rect 227562 581606 227772 581612
rect 227562 581590 227760 581606
rect 229388 581369 229416 582111
rect 229466 582040 229522 582049
rect 229466 581975 229522 581984
rect 229480 581505 229508 581975
rect 229756 581876 229784 582898
rect 230110 581904 230166 581913
rect 234540 581876 234568 583743
rect 236458 582040 236514 582049
rect 236458 581975 236514 581984
rect 230110 581839 230166 581848
rect 229466 581496 229522 581505
rect 229466 581431 229522 581440
rect 230124 581369 230152 581839
rect 236472 581505 236500 581975
rect 236932 581876 236960 586502
rect 238758 584760 238814 584769
rect 238758 584695 238760 584704
rect 238812 584695 238814 584704
rect 244096 584724 244148 584730
rect 238760 584666 238812 584672
rect 244096 584666 244148 584672
rect 241702 584216 241758 584225
rect 241702 584151 241758 584160
rect 238758 582040 238814 582049
rect 238758 581975 238814 581984
rect 236458 581496 236514 581505
rect 236458 581431 236514 581440
rect 238772 581369 238800 581975
rect 239034 581904 239090 581913
rect 241716 581876 241744 584151
rect 244108 581876 244136 584666
rect 249708 584656 249760 584662
rect 249708 584598 249760 584604
rect 248880 584588 248932 584594
rect 248880 584530 248932 584536
rect 248892 581876 248920 584530
rect 249246 581904 249302 581913
rect 239034 581839 239090 581848
rect 249246 581839 249302 581848
rect 239048 581369 239076 581839
rect 246856 581800 246908 581806
rect 246514 581748 246856 581754
rect 246514 581742 246908 581748
rect 246514 581726 246896 581742
rect 249260 581369 249288 581839
rect 249720 581738 249748 584598
rect 258446 584216 258502 584225
rect 258446 584151 258502 584160
rect 256056 583228 256108 583234
rect 256056 583170 256108 583176
rect 256068 581876 256096 583170
rect 258354 582176 258410 582185
rect 258354 582111 258410 582120
rect 258170 582040 258226 582049
rect 258170 581975 258226 581984
rect 256238 581904 256294 581913
rect 256238 581839 256294 581848
rect 251298 581738 251680 581754
rect 249708 581732 249760 581738
rect 251298 581732 251692 581738
rect 251298 581726 251640 581732
rect 249708 581674 249760 581680
rect 251640 581674 251692 581680
rect 256252 581505 256280 581839
rect 256330 581632 256386 581641
rect 256330 581567 256386 581576
rect 253386 581496 253442 581505
rect 256238 581496 256294 581505
rect 253442 581454 253690 581482
rect 253386 581431 253442 581440
rect 256238 581431 256294 581440
rect 256344 581369 256372 581567
rect 258184 581369 258212 581975
rect 258368 581369 258396 582111
rect 258460 581876 258488 584151
rect 269040 583982 269068 700674
rect 294144 584792 294196 584798
rect 294144 584734 294196 584740
rect 291750 584624 291806 584633
rect 291750 584559 291806 584568
rect 270408 584520 270460 584526
rect 270408 584462 270460 584468
rect 275006 584488 275062 584497
rect 268016 583976 268068 583982
rect 268016 583918 268068 583924
rect 269028 583976 269080 583982
rect 269028 583918 269080 583924
rect 265624 583160 265676 583166
rect 265624 583102 265676 583108
rect 262968 581874 263258 581890
rect 265636 581876 265664 583102
rect 268028 581876 268056 583918
rect 270420 581876 270448 584462
rect 272800 584452 272852 584458
rect 275006 584423 275062 584432
rect 272800 584394 272852 584400
rect 272812 581876 272840 584394
rect 273166 582176 273222 582185
rect 273166 582111 273222 582120
rect 262956 581868 263258 581874
rect 263008 581862 263258 581868
rect 262956 581810 263008 581816
rect 273180 581641 273208 582111
rect 275020 581876 275048 584423
rect 277398 584352 277454 584361
rect 277398 584287 277454 584296
rect 277412 581876 277440 584287
rect 289360 583976 289412 583982
rect 289360 583918 289412 583924
rect 279792 583296 279844 583302
rect 279792 583238 279844 583244
rect 279804 581876 279832 583238
rect 284576 583092 284628 583098
rect 284576 583034 284628 583040
rect 282918 582312 282974 582321
rect 282918 582247 282974 582256
rect 282550 581904 282606 581913
rect 282210 581862 282550 581890
rect 282550 581839 282606 581848
rect 282932 581641 282960 582247
rect 284588 581876 284616 583034
rect 286692 582072 286744 582078
rect 286692 582014 286744 582020
rect 286704 581890 286732 582014
rect 286704 581862 286994 581890
rect 289372 581876 289400 583918
rect 291764 581876 291792 584559
rect 292486 582312 292542 582321
rect 292486 582247 292542 582256
rect 292500 581641 292528 582247
rect 294156 581876 294184 584734
rect 315670 584624 315726 584633
rect 315670 584559 315726 584568
rect 310888 584316 310940 584322
rect 310888 584258 310940 584264
rect 298926 583808 298982 583817
rect 298926 583743 298982 583752
rect 308496 583772 308548 583778
rect 296562 581874 296760 581890
rect 298940 581876 298968 583743
rect 308496 583714 308548 583720
rect 303710 582992 303766 583001
rect 303710 582927 303766 582936
rect 301318 582720 301374 582729
rect 301318 582655 301374 582664
rect 301332 581876 301360 582655
rect 302238 582312 302294 582321
rect 302238 582247 302294 582256
rect 296562 581868 296772 581874
rect 296562 581862 296720 581868
rect 296720 581810 296772 581816
rect 302252 581641 302280 582247
rect 303724 581876 303752 582927
rect 306286 582040 306342 582049
rect 306286 581975 306342 581984
rect 306300 581890 306328 581975
rect 306130 581862 306328 581890
rect 308508 581876 308536 583714
rect 310900 581876 310928 584258
rect 314660 583772 314712 583778
rect 314660 583714 314712 583720
rect 314672 583001 314700 583714
rect 314658 582992 314714 583001
rect 314658 582927 314714 582936
rect 311806 582312 311862 582321
rect 311806 582247 311862 582256
rect 311820 581641 311848 582247
rect 315684 581876 315712 584559
rect 322664 584384 322716 584390
rect 322664 584326 322716 584332
rect 318062 582856 318118 582865
rect 318062 582791 318118 582800
rect 318076 581876 318104 582791
rect 320180 582004 320232 582010
rect 320180 581946 320232 581952
rect 321560 582004 321612 582010
rect 321560 581946 321612 581952
rect 320192 581890 320220 581946
rect 320192 581862 320298 581890
rect 321572 581641 321600 581946
rect 322676 581876 322704 584326
rect 327448 583092 327500 583098
rect 327448 583034 327500 583040
rect 326434 582176 326490 582185
rect 326434 582111 326490 582120
rect 326448 582010 326476 582111
rect 326436 582004 326488 582010
rect 326436 581946 326488 581952
rect 327460 581876 327488 583034
rect 329838 582176 329894 582185
rect 329838 582111 329894 582120
rect 329852 581876 329880 582111
rect 331954 581768 332010 581777
rect 335280 581754 335308 700810
rect 343640 700800 343692 700806
rect 343640 700742 343692 700748
rect 341800 584316 341852 584322
rect 341800 584258 341852 584264
rect 339408 584248 339460 584254
rect 339408 584190 339460 584196
rect 337016 583160 337068 583166
rect 337016 583102 337068 583108
rect 337028 581876 337056 583102
rect 339420 581876 339448 584190
rect 341812 581876 341840 584258
rect 332010 581726 332258 581754
rect 334650 581726 335308 581754
rect 343652 581754 343680 700742
rect 348804 700369 348832 703520
rect 364996 700806 365024 703520
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 397472 700670 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 386420 700664 386472 700670
rect 386420 700606 386472 700612
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 348790 700360 348846 700369
rect 348790 700295 348846 700304
rect 372618 584760 372674 584769
rect 372618 584695 372674 584704
rect 348976 584588 349028 584594
rect 348976 584530 349028 584536
rect 348988 581876 349016 584530
rect 367928 584384 367980 584390
rect 367928 584326 367980 584332
rect 356152 584180 356204 584186
rect 356152 584122 356204 584128
rect 353760 583024 353812 583030
rect 353760 582966 353812 582972
rect 353772 581876 353800 582966
rect 356164 581876 356192 584122
rect 360936 583024 360988 583030
rect 360936 582966 360988 582972
rect 360948 581876 360976 582966
rect 363696 582004 363748 582010
rect 363696 581946 363748 581952
rect 363708 581890 363736 581946
rect 363354 581862 363736 581890
rect 367940 581876 367968 584326
rect 370320 584180 370372 584186
rect 370320 584122 370372 584128
rect 370332 581876 370360 584122
rect 372632 581942 372660 584695
rect 372712 584656 372764 584662
rect 372712 584598 372764 584604
rect 377496 584656 377548 584662
rect 377496 584598 377548 584604
rect 372620 581936 372672 581942
rect 372620 581878 372672 581884
rect 372724 581876 372752 584598
rect 377508 581876 377536 584598
rect 382280 584520 382332 584526
rect 382280 584462 382332 584468
rect 379888 583228 379940 583234
rect 379888 583170 379940 583176
rect 379900 581876 379928 583170
rect 382292 581876 382320 584462
rect 386432 581754 386460 700606
rect 402980 700528 403032 700534
rect 402980 700470 403032 700476
rect 401416 582208 401468 582214
rect 401416 582150 401468 582156
rect 394608 582072 394660 582078
rect 394608 582014 394660 582020
rect 394620 581890 394648 582014
rect 399392 581936 399444 581942
rect 394266 581862 394648 581890
rect 399050 581884 399392 581890
rect 399050 581878 399444 581884
rect 399050 581862 399432 581878
rect 401428 581876 401456 582150
rect 402992 581754 403020 700470
rect 413756 698290 413784 703446
rect 429856 700874 429884 703520
rect 429844 700868 429896 700874
rect 429844 700810 429896 700816
rect 462332 700466 462360 703520
rect 462320 700460 462372 700466
rect 462320 700402 462372 700408
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 508136 700800 508188 700806
rect 508136 700742 508188 700748
rect 501604 700732 501656 700738
rect 501604 700674 501656 700680
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 413112 659682 413140 666538
rect 412928 659654 413140 659682
rect 412928 647290 412956 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 412836 640422 412864 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 412928 630698 412956 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 412744 630578 412772 630634
rect 412744 630550 412864 630578
rect 412836 621058 412864 630550
rect 412836 621030 412956 621058
rect 412928 611386 412956 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 412744 611266 412772 611322
rect 412744 611238 412864 611266
rect 412836 608598 412864 611238
rect 412824 608592 412876 608598
rect 412824 608534 412876 608540
rect 413008 601724 413060 601730
rect 413008 601666 413060 601672
rect 413020 598942 413048 601666
rect 413008 598936 413060 598942
rect 413008 598878 413060 598884
rect 412916 589348 412968 589354
rect 412916 589290 412968 589296
rect 412928 585721 412956 589290
rect 412914 585712 412970 585721
rect 412914 585647 412970 585656
rect 477592 585132 477644 585138
rect 477592 585074 477644 585080
rect 487160 585132 487212 585138
rect 487160 585074 487212 585080
rect 432328 585064 432380 585070
rect 432328 585006 432380 585012
rect 439504 585064 439556 585070
rect 439504 585006 439556 585012
rect 427542 584896 427598 584905
rect 427542 584831 427598 584840
rect 413192 583908 413244 583914
rect 413192 583850 413244 583856
rect 422760 583908 422812 583914
rect 422760 583850 422812 583856
rect 408592 583772 408644 583778
rect 408592 583714 408644 583720
rect 406200 582140 406252 582146
rect 406200 582082 406252 582088
rect 406212 581876 406240 582082
rect 408604 581876 408632 583714
rect 410800 583296 410852 583302
rect 410800 583238 410852 583244
rect 410812 581876 410840 583238
rect 413204 581876 413232 583850
rect 415584 583840 415636 583846
rect 415584 583782 415636 583788
rect 415596 581876 415624 583782
rect 422772 581876 422800 583850
rect 424968 583772 425020 583778
rect 424968 583714 425020 583720
rect 424980 582185 425008 583714
rect 425152 582616 425204 582622
rect 425152 582558 425204 582564
rect 424966 582176 425022 582185
rect 424966 582111 425022 582120
rect 425164 581876 425192 582558
rect 427556 581876 427584 584831
rect 429936 583772 429988 583778
rect 429936 583714 429988 583720
rect 429948 581876 429976 583714
rect 432340 581876 432368 585006
rect 437112 584792 437164 584798
rect 437112 584734 437164 584740
rect 437124 581876 437152 584734
rect 439516 581876 439544 585006
rect 468024 584996 468076 585002
rect 468024 584938 468076 584944
rect 475200 584996 475252 585002
rect 475200 584938 475252 584944
rect 446680 584860 446732 584866
rect 446680 584802 446732 584808
rect 444288 584452 444340 584458
rect 444288 584394 444340 584400
rect 441896 583500 441948 583506
rect 441896 583442 441948 583448
rect 441908 581876 441936 583442
rect 444300 581876 444328 584394
rect 446692 581876 446720 584802
rect 465630 584760 465686 584769
rect 456064 584724 456116 584730
rect 465630 584695 465686 584704
rect 456064 584666 456116 584672
rect 449072 584112 449124 584118
rect 449072 584054 449124 584060
rect 453856 584112 453908 584118
rect 453856 584054 453908 584060
rect 449084 581876 449112 584054
rect 451462 583808 451518 583817
rect 451462 583743 451518 583752
rect 451476 581876 451504 583743
rect 453868 581876 453896 584054
rect 455328 583976 455380 583982
rect 455328 583918 455380 583924
rect 455340 583370 455368 583918
rect 455328 583364 455380 583370
rect 455328 583306 455380 583312
rect 456076 581876 456104 584666
rect 456800 584248 456852 584254
rect 456800 584190 456852 584196
rect 458456 584248 458508 584254
rect 458456 584190 458508 584196
rect 456812 583438 456840 584190
rect 456800 583432 456852 583438
rect 456800 583374 456852 583380
rect 458468 581876 458496 584190
rect 463240 582480 463292 582486
rect 463240 582422 463292 582428
rect 460848 582344 460900 582350
rect 460848 582286 460900 582292
rect 460860 581876 460888 582286
rect 463252 581876 463280 582422
rect 465644 581876 465672 584695
rect 468036 581876 468064 584938
rect 470416 584928 470468 584934
rect 470416 584870 470468 584876
rect 470428 581876 470456 584870
rect 472806 584760 472862 584769
rect 472806 584695 472862 584704
rect 472820 581876 472848 584695
rect 475212 581876 475240 584938
rect 477604 581876 477632 585074
rect 479984 584928 480036 584934
rect 479984 584870 480036 584876
rect 479996 581876 480024 584870
rect 485780 584588 485832 584594
rect 485780 584530 485832 584536
rect 484768 583976 484820 583982
rect 484768 583918 484820 583924
rect 482376 582480 482428 582486
rect 482376 582422 482428 582428
rect 482388 581876 482416 582422
rect 484780 581876 484808 583918
rect 485792 583506 485820 584530
rect 485780 583500 485832 583506
rect 485780 583442 485832 583448
rect 487172 581876 487200 585074
rect 494704 584656 494756 584662
rect 494704 584598 494756 584604
rect 491944 584588 491996 584594
rect 491944 584530 491996 584536
rect 490380 584044 490432 584050
rect 490380 583986 490432 583992
rect 489552 582412 489604 582418
rect 489552 582354 489604 582360
rect 490196 582412 490248 582418
rect 490196 582354 490248 582360
rect 489564 581876 489592 582354
rect 490208 582321 490236 582354
rect 490392 582321 490420 583986
rect 490194 582312 490250 582321
rect 490194 582247 490250 582256
rect 490378 582312 490434 582321
rect 490378 582247 490434 582256
rect 491850 582176 491906 582185
rect 491850 582111 491906 582120
rect 418158 581768 418214 581777
rect 343652 581726 344218 581754
rect 386432 581726 387090 581754
rect 402992 581726 403834 581754
rect 418002 581726 418158 581754
rect 331954 581703 332010 581712
rect 418158 581703 418214 581712
rect 273166 581632 273222 581641
rect 273166 581567 273222 581576
rect 282918 581632 282974 581641
rect 282918 581567 282974 581576
rect 292486 581632 292542 581641
rect 292486 581567 292542 581576
rect 302238 581632 302294 581641
rect 302238 581567 302294 581576
rect 311806 581632 311862 581641
rect 321558 581632 321614 581641
rect 313200 581602 313306 581618
rect 311806 581567 311862 581576
rect 313188 581596 313306 581602
rect 313240 581590 313306 581596
rect 321558 581567 321614 581576
rect 324778 581632 324834 581641
rect 346858 581632 346914 581641
rect 324834 581590 325082 581618
rect 346610 581590 346858 581618
rect 324778 581567 324834 581576
rect 351642 581632 351698 581641
rect 351394 581590 351642 581618
rect 346858 581567 346914 581576
rect 351642 581567 351698 581576
rect 365258 581632 365314 581641
rect 384854 581632 384910 581641
rect 365314 581590 365562 581618
rect 375130 581602 375328 581618
rect 375130 581596 375340 581602
rect 375130 581590 375288 581596
rect 365258 581567 365314 581576
rect 313188 581538 313240 581544
rect 384698 581590 384854 581618
rect 389730 581632 389786 581641
rect 389482 581590 389730 581618
rect 384854 581567 384910 581576
rect 389730 581567 389786 581576
rect 391754 581632 391810 581641
rect 396998 581632 397054 581641
rect 391810 581590 391874 581618
rect 396658 581590 396998 581618
rect 391754 581567 391810 581576
rect 396998 581567 397054 581576
rect 375288 581538 375340 581544
rect 263506 581496 263562 581505
rect 263690 581496 263746 581505
rect 263562 581454 263690 581482
rect 263506 581431 263562 581440
rect 420104 581466 420394 581482
rect 263690 581431 263746 581440
rect 420092 581460 420394 581466
rect 420144 581454 420394 581460
rect 434746 581466 435128 581482
rect 434746 581460 435140 581466
rect 434746 581454 435088 581460
rect 420092 581402 420144 581408
rect 435088 581402 435140 581408
rect 491864 581398 491892 582111
rect 491956 581876 491984 584530
rect 494336 584044 494388 584050
rect 494336 583986 494388 583992
rect 494348 581876 494376 583986
rect 494610 583944 494666 583953
rect 494610 583879 494666 583888
rect 494624 581398 494652 583879
rect 494716 582282 494744 584598
rect 501512 584316 501564 584322
rect 501512 584258 501564 584264
rect 496726 583944 496782 583953
rect 496726 583879 496782 583888
rect 494704 582276 494756 582282
rect 494704 582218 494756 582224
rect 496740 581876 496768 583879
rect 501328 583772 501380 583778
rect 501328 583714 501380 583720
rect 499120 582548 499172 582554
rect 499120 582490 499172 582496
rect 497556 582412 497608 582418
rect 497556 582354 497608 582360
rect 497568 582049 497596 582354
rect 497554 582040 497610 582049
rect 497554 581975 497610 581984
rect 499132 581876 499160 582490
rect 501340 581876 501368 583714
rect 491852 581392 491904 581398
rect 171612 581318 171916 581346
rect 176566 581360 176622 581369
rect 166906 581295 166962 581304
rect 176566 581295 176622 581304
rect 176750 581360 176806 581369
rect 176750 581295 176806 581304
rect 192022 581360 192078 581369
rect 192022 581295 192078 581304
rect 192206 581360 192262 581369
rect 192206 581295 192262 581304
rect 195886 581360 195942 581369
rect 195886 581295 195942 581304
rect 200670 581360 200726 581369
rect 200670 581295 200726 581304
rect 210330 581360 210386 581369
rect 210330 581295 210386 581304
rect 211158 581360 211214 581369
rect 211158 581295 211214 581304
rect 220726 581360 220782 581369
rect 220726 581295 220782 581304
rect 220910 581360 220966 581369
rect 220910 581295 220966 581304
rect 229374 581360 229430 581369
rect 229374 581295 229430 581304
rect 230110 581360 230166 581369
rect 230110 581295 230166 581304
rect 231950 581360 232006 581369
rect 238758 581360 238814 581369
rect 232006 581318 232162 581346
rect 231950 581295 232006 581304
rect 238758 581295 238814 581304
rect 239034 581360 239090 581369
rect 239678 581360 239734 581369
rect 239338 581318 239678 581346
rect 239034 581295 239090 581304
rect 239678 581295 239734 581304
rect 249246 581360 249302 581369
rect 249246 581295 249302 581304
rect 256330 581360 256386 581369
rect 256330 581295 256386 581304
rect 258170 581360 258226 581369
rect 258170 581295 258226 581304
rect 258354 581360 258410 581369
rect 258354 581295 258410 581304
rect 263506 581360 263562 581369
rect 263690 581360 263746 581369
rect 263562 581318 263690 581346
rect 263506 581295 263562 581304
rect 358726 581360 358782 581369
rect 358570 581318 358726 581346
rect 263690 581295 263746 581304
rect 491852 581334 491904 581340
rect 494612 581392 494664 581398
rect 494612 581334 494664 581340
rect 358726 581295 358782 581304
rect 83660 574790 83780 574818
rect 83752 547074 83780 574790
rect 83568 547046 83780 547074
rect 83568 545034 83596 547046
rect 83568 545006 83780 545034
rect 82634 541512 82690 541521
rect 82690 541470 82860 541498
rect 82634 541447 82690 541456
rect 82832 529922 82860 541470
rect 83752 530074 83780 545006
rect 83568 530046 83780 530074
rect 83568 529938 83596 530046
rect 82820 529916 82872 529922
rect 83568 529910 83688 529938
rect 82820 529858 82872 529864
rect 83660 528578 83688 529910
rect 83568 528550 83688 528578
rect 82912 520328 82964 520334
rect 82832 520276 82912 520282
rect 82832 520270 82964 520276
rect 82832 520254 82952 520270
rect 82358 518800 82414 518809
rect 82358 518735 82414 518744
rect 82372 509561 82400 518735
rect 82358 509552 82414 509561
rect 82358 509487 82414 509496
rect 82542 505744 82598 505753
rect 82542 505679 82598 505688
rect 82358 500848 82414 500857
rect 82358 500783 82414 500792
rect 82372 497185 82400 500783
rect 82556 498137 82584 505679
rect 82832 501090 82860 520254
rect 83568 518514 83596 528550
rect 83568 518486 83688 518514
rect 83660 518242 83688 518486
rect 83568 518214 83688 518242
rect 83568 516066 83596 518214
rect 83568 516038 83780 516066
rect 83752 504914 83780 516038
rect 83292 504886 83780 504914
rect 82820 501084 82872 501090
rect 82820 501026 82872 501032
rect 82912 501016 82964 501022
rect 82832 500964 82912 500970
rect 82832 500958 82964 500964
rect 82832 500954 82952 500958
rect 82820 500948 82952 500954
rect 82872 500942 82952 500948
rect 82820 500890 82872 500896
rect 82832 500859 82860 500890
rect 82542 498128 82598 498137
rect 82542 498063 82598 498072
rect 82358 497176 82414 497185
rect 82358 497111 82414 497120
rect 83292 493354 83320 504886
rect 83292 493326 83504 493354
rect 82820 491360 82872 491366
rect 82820 491302 82872 491308
rect 82542 486160 82598 486169
rect 82542 486095 82598 486104
rect 82358 481264 82414 481273
rect 82358 481199 82414 481208
rect 82372 473657 82400 481199
rect 82556 481137 82584 486095
rect 82542 481128 82598 481137
rect 82542 481063 82598 481072
rect 82542 475824 82598 475833
rect 82542 475759 82598 475768
rect 82450 474192 82506 474201
rect 82450 474127 82506 474136
rect 82358 473648 82414 473657
rect 82358 473583 82414 473592
rect 82464 466177 82492 474127
rect 82556 473521 82584 475759
rect 82634 474328 82690 474337
rect 82634 474263 82690 474272
rect 82648 474094 82676 474263
rect 82636 474088 82688 474094
rect 82636 474030 82688 474036
rect 82542 473512 82598 473521
rect 82542 473447 82598 473456
rect 82542 471064 82598 471073
rect 82542 470999 82598 471008
rect 82450 466168 82506 466177
rect 82450 466103 82506 466112
rect 82556 458017 82584 470999
rect 82542 458008 82598 458017
rect 82542 457943 82598 457952
rect 82634 453384 82690 453393
rect 82634 453319 82690 453328
rect 82648 450226 82676 453319
rect 82636 450220 82688 450226
rect 82636 450162 82688 450168
rect 82832 442950 82860 491302
rect 83476 483018 83504 493326
rect 83476 482990 83596 483018
rect 83568 478802 83596 482990
rect 83568 478774 83688 478802
rect 82912 474088 82964 474094
rect 82912 474030 82964 474036
rect 82924 473906 82952 474030
rect 82924 473878 83412 473906
rect 82912 450220 82964 450226
rect 82912 450162 82964 450168
rect 82820 442944 82872 442950
rect 82820 442886 82872 442892
rect 82820 442196 82872 442202
rect 82820 442138 82872 442144
rect 82832 439906 82860 442138
rect 82924 442082 82952 450162
rect 83384 447930 83412 473878
rect 83016 447902 83412 447930
rect 83016 447846 83044 447902
rect 83004 447840 83056 447846
rect 83004 447782 83056 447788
rect 83660 447658 83688 478774
rect 101586 456512 101642 456521
rect 101586 456447 101642 456456
rect 101600 452418 101628 456447
rect 101508 452390 101628 452418
rect 101508 451897 101536 452390
rect 101494 451888 101550 451897
rect 101494 451823 101550 451832
rect 83016 447630 83688 447658
rect 83016 442202 83044 447630
rect 83004 442196 83056 442202
rect 83004 442138 83056 442144
rect 83108 442190 83688 442218
rect 83108 442082 83136 442190
rect 82924 442054 83136 442082
rect 82832 439878 83596 439906
rect 82912 439544 82964 439550
rect 82964 439492 83412 439498
rect 82912 439486 83412 439492
rect 82924 439470 83412 439486
rect 82542 438968 82598 438977
rect 82542 438903 82598 438912
rect 82556 435441 82584 438903
rect 82820 438184 82872 438190
rect 82820 438126 82872 438132
rect 82542 435432 82598 435441
rect 82542 435367 82598 435376
rect 82542 431216 82598 431225
rect 82542 431151 82598 431160
rect 82556 406473 82584 431151
rect 82832 423638 82860 438126
rect 83384 425082 83412 439470
rect 83568 433378 83596 439878
rect 83476 433350 83596 433378
rect 83660 433378 83688 442190
rect 83660 433350 83780 433378
rect 83476 425218 83504 433350
rect 83752 433242 83780 433350
rect 83660 433214 83780 433242
rect 83476 425190 83596 425218
rect 83384 425054 83504 425082
rect 82820 423632 82872 423638
rect 82820 423574 82872 423580
rect 82912 423020 82964 423026
rect 83476 423008 83504 425054
rect 82964 422980 83504 423008
rect 82912 422962 82964 422968
rect 83568 422906 83596 425190
rect 83384 422878 83596 422906
rect 82912 419008 82964 419014
rect 82964 418956 83136 418962
rect 82912 418950 83136 418956
rect 82924 418934 83136 418950
rect 82820 414044 82872 414050
rect 82820 413986 82872 413992
rect 82542 406464 82598 406473
rect 82542 406399 82598 406408
rect 82542 401568 82598 401577
rect 82542 401503 82598 401512
rect 82358 400208 82414 400217
rect 82358 400143 82414 400152
rect 82266 391232 82322 391241
rect 82266 391167 82322 391176
rect 82082 391096 82138 391105
rect 82082 391031 82138 391040
rect 82280 388006 82308 391167
rect 82084 388000 82136 388006
rect 82084 387942 82136 387948
rect 82268 388000 82320 388006
rect 82268 387942 82320 387948
rect 82096 385665 82124 387942
rect 82372 385665 82400 400143
rect 82450 396808 82506 396817
rect 82450 396743 82506 396752
rect 82464 396137 82492 396743
rect 82450 396128 82506 396137
rect 82450 396063 82506 396072
rect 82556 385801 82584 401503
rect 82634 393136 82690 393145
rect 82634 393071 82690 393080
rect 82542 385792 82598 385801
rect 82542 385727 82598 385736
rect 82082 385656 82138 385665
rect 82082 385591 82138 385600
rect 82358 385656 82414 385665
rect 82358 385591 82414 385600
rect 82268 375352 82320 375358
rect 82268 375294 82320 375300
rect 82280 370870 82308 375294
rect 82450 371920 82506 371929
rect 82450 371855 82506 371864
rect 82268 370864 82320 370870
rect 82268 370806 82320 370812
rect 82358 369064 82414 369073
rect 82358 368999 82414 369008
rect 82372 364721 82400 368999
rect 82464 368121 82492 371855
rect 82542 369064 82598 369073
rect 82542 368999 82598 369008
rect 82450 368112 82506 368121
rect 82450 368047 82506 368056
rect 82556 366858 82584 368999
rect 82648 368937 82676 393071
rect 82832 385014 82860 413986
rect 83108 406314 83136 418934
rect 83384 415426 83412 422878
rect 83384 415398 83504 415426
rect 83476 414066 83504 415398
rect 82924 406298 83136 406314
rect 82912 406292 83136 406298
rect 82964 406286 83136 406292
rect 83384 414038 83504 414066
rect 82912 406234 82964 406240
rect 83384 404410 83412 414038
rect 83292 404382 83412 404410
rect 83292 400738 83320 404382
rect 83016 400722 83320 400738
rect 83004 400716 83320 400722
rect 83056 400710 83320 400716
rect 83004 400658 83056 400664
rect 83660 400602 83688 433214
rect 83016 400574 83688 400602
rect 83016 400382 83044 400574
rect 83004 400376 83056 400382
rect 83004 400318 83056 400324
rect 83004 400240 83056 400246
rect 83056 400200 83412 400228
rect 83004 400182 83056 400188
rect 83004 399560 83056 399566
rect 83004 399502 83056 399508
rect 83016 394754 83044 399502
rect 83384 398834 83412 400200
rect 83384 398806 83504 398834
rect 83016 394726 83136 394754
rect 83108 389994 83136 394726
rect 83108 389966 83228 389994
rect 83200 389586 83228 389966
rect 83476 389858 83504 398806
rect 83476 389830 83596 389858
rect 83200 389558 83504 389586
rect 83004 387932 83056 387938
rect 83004 387874 83056 387880
rect 82820 385008 82872 385014
rect 82820 384950 82872 384956
rect 83016 382922 83044 387874
rect 83476 383738 83504 389558
rect 83568 387818 83596 389830
rect 83568 387790 83688 387818
rect 83384 383710 83504 383738
rect 83016 382894 83320 382922
rect 82820 375488 82872 375494
rect 82820 375430 82872 375436
rect 82832 375358 82860 375430
rect 82820 375352 82872 375358
rect 82820 375294 82872 375300
rect 83292 373130 83320 382894
rect 82924 373102 83320 373130
rect 82924 369050 82952 373102
rect 83384 372858 83412 383710
rect 83016 372830 83412 372858
rect 83016 372774 83044 372830
rect 83004 372768 83056 372774
rect 83004 372710 83056 372716
rect 83004 372632 83056 372638
rect 83056 372592 83136 372620
rect 83004 372574 83056 372580
rect 83004 372496 83056 372502
rect 83004 372438 83056 372444
rect 83108 372450 83136 372592
rect 83660 372450 83688 387790
rect 83016 369866 83044 372438
rect 83108 372422 83688 372450
rect 83016 369838 83780 369866
rect 83004 369368 83056 369374
rect 83056 369316 83596 369322
rect 83004 369310 83596 369316
rect 83016 369294 83596 369310
rect 83200 369158 83412 369186
rect 83200 369050 83228 369158
rect 82924 369022 83228 369050
rect 82634 368928 82690 368937
rect 82634 368863 82690 368872
rect 82634 368792 82690 368801
rect 82634 368727 82690 368736
rect 82544 366852 82596 366858
rect 82544 366794 82596 366800
rect 82544 365288 82596 365294
rect 82544 365230 82596 365236
rect 82450 364848 82506 364857
rect 82450 364783 82506 364792
rect 82358 364712 82414 364721
rect 82358 364647 82414 364656
rect 82358 362944 82414 362953
rect 82358 362879 82414 362888
rect 82372 360233 82400 362879
rect 82358 360224 82414 360233
rect 82358 360159 82414 360168
rect 82464 359417 82492 364783
rect 82556 360210 82584 365230
rect 82648 362817 82676 368727
rect 82912 366852 82964 366858
rect 82912 366794 82964 366800
rect 82924 364698 82952 366794
rect 82924 364670 83228 364698
rect 82634 362808 82690 362817
rect 82634 362743 82690 362752
rect 82556 360182 82952 360210
rect 82634 360088 82690 360097
rect 82634 360023 82690 360032
rect 82450 359408 82506 359417
rect 82450 359343 82506 359352
rect 82648 358057 82676 360023
rect 82634 358048 82690 358057
rect 82634 357983 82690 357992
rect 82924 354770 82952 360182
rect 82832 354742 82952 354770
rect 82082 354648 82138 354657
rect 82082 354583 82138 354592
rect 82096 123690 82124 354583
rect 82542 347032 82598 347041
rect 82542 346967 82598 346976
rect 82174 339688 82230 339697
rect 82174 339623 82230 339632
rect 82188 338065 82216 339623
rect 82358 339008 82414 339017
rect 82358 338943 82414 338952
rect 82174 338056 82230 338065
rect 82174 337991 82230 338000
rect 82174 332208 82230 332217
rect 82174 332143 82230 332152
rect 82188 328137 82216 332143
rect 82372 331265 82400 338943
rect 82556 336977 82584 346967
rect 82832 345030 82860 354742
rect 83200 349874 83228 364670
rect 83108 349846 83228 349874
rect 83108 347154 83136 349846
rect 83016 347126 83136 347154
rect 83016 345114 83044 347126
rect 83016 345086 83320 345114
rect 82820 345024 82872 345030
rect 82820 344966 82872 344972
rect 82912 345024 82964 345030
rect 82912 344966 82964 344972
rect 82634 341728 82690 341737
rect 82634 341663 82690 341672
rect 82542 336968 82598 336977
rect 82542 336903 82598 336912
rect 82542 335064 82598 335073
rect 82542 334999 82598 335008
rect 82358 331256 82414 331265
rect 82358 331191 82414 331200
rect 82556 331129 82584 334999
rect 82648 331265 82676 341663
rect 82634 331256 82690 331265
rect 82634 331191 82690 331200
rect 82542 331120 82598 331129
rect 82542 331055 82598 331064
rect 82924 328574 82952 344966
rect 83292 342802 83320 345086
rect 83016 342774 83320 342802
rect 82912 328568 82964 328574
rect 82912 328510 82964 328516
rect 82820 328500 82872 328506
rect 82820 328442 82872 328448
rect 82174 328128 82230 328137
rect 82174 328063 82230 328072
rect 82634 319560 82690 319569
rect 82634 319495 82690 319504
rect 82450 317384 82506 317393
rect 82450 317319 82506 317328
rect 82464 316305 82492 317319
rect 82450 316296 82506 316305
rect 82450 316231 82506 316240
rect 82648 315994 82676 319495
rect 82728 316124 82780 316130
rect 82728 316066 82780 316072
rect 82636 315988 82688 315994
rect 82636 315930 82688 315936
rect 82634 312488 82690 312497
rect 82634 312423 82690 312432
rect 82450 312352 82506 312361
rect 82450 312287 82506 312296
rect 82464 307465 82492 312287
rect 82648 310758 82676 312423
rect 82636 310752 82688 310758
rect 82636 310694 82688 310700
rect 82740 310298 82768 316066
rect 82832 313342 82860 328442
rect 83016 328386 83044 342774
rect 83384 332602 83412 369158
rect 83384 332574 83504 332602
rect 83016 328358 83136 328386
rect 83108 328250 83136 328358
rect 83108 328222 83228 328250
rect 83200 327026 83228 328222
rect 83016 327010 83228 327026
rect 83004 327004 83228 327010
rect 83056 326998 83228 327004
rect 83004 326946 83056 326952
rect 83016 317490 83320 317506
rect 83004 317484 83320 317490
rect 83056 317478 83320 317484
rect 83004 317426 83056 317432
rect 83292 317370 83320 317478
rect 82924 317342 83320 317370
rect 82924 316130 82952 317342
rect 82912 316124 82964 316130
rect 82912 316066 82964 316072
rect 82912 315988 82964 315994
rect 82964 315948 83044 315976
rect 82912 315930 82964 315936
rect 82820 313336 82872 313342
rect 82820 313278 82872 313284
rect 83016 311386 83044 315948
rect 83476 312474 83504 332574
rect 82924 311370 83044 311386
rect 82912 311364 83044 311370
rect 82964 311358 83044 311364
rect 83384 312446 83504 312474
rect 82912 311306 82964 311312
rect 83384 311114 83412 312446
rect 82924 311086 83412 311114
rect 82924 310434 82952 311086
rect 83568 310978 83596 369294
rect 83016 310950 83596 310978
rect 83016 310894 83044 310950
rect 83004 310888 83056 310894
rect 83004 310830 83056 310836
rect 83004 310752 83056 310758
rect 83056 310712 83320 310740
rect 83004 310694 83056 310700
rect 83004 310616 83056 310622
rect 83056 310564 83228 310570
rect 83004 310558 83228 310564
rect 83016 310542 83228 310558
rect 82924 310406 83044 310434
rect 82740 310270 82952 310298
rect 82820 309120 82872 309126
rect 82820 309062 82872 309068
rect 82450 307456 82506 307465
rect 82450 307391 82506 307400
rect 82634 305416 82690 305425
rect 82634 305351 82690 305360
rect 82174 301880 82230 301889
rect 82174 301815 82230 301824
rect 82084 123684 82136 123690
rect 82084 123626 82136 123632
rect 82082 123584 82138 123593
rect 81992 123548 82044 123554
rect 82082 123519 82138 123528
rect 81992 123490 82044 123496
rect 82096 123486 82124 123519
rect 82084 123480 82136 123486
rect 82084 123422 82136 123428
rect 81992 123412 82044 123418
rect 81992 123354 82044 123360
rect 82004 118046 82032 123354
rect 82188 123298 82216 301815
rect 82648 300558 82676 305351
rect 82832 303346 82860 309062
rect 82924 303346 82952 310270
rect 82820 303340 82872 303346
rect 82820 303282 82872 303288
rect 82912 303340 82964 303346
rect 82912 303282 82964 303288
rect 83016 303090 83044 310406
rect 82924 303074 83044 303090
rect 82912 303068 83044 303074
rect 82964 303062 83044 303068
rect 82912 303010 82964 303016
rect 82820 302932 82872 302938
rect 82820 302874 82872 302880
rect 82912 302932 82964 302938
rect 82912 302874 82964 302880
rect 82636 300552 82688 300558
rect 82636 300494 82688 300500
rect 82728 298308 82780 298314
rect 82728 298250 82780 298256
rect 82542 297800 82598 297809
rect 82542 297735 82598 297744
rect 82358 296848 82414 296857
rect 82358 296783 82414 296792
rect 82266 294808 82322 294817
rect 82266 294743 82322 294752
rect 82280 123418 82308 294743
rect 82372 291281 82400 296783
rect 82358 291272 82414 291281
rect 82358 291207 82414 291216
rect 82556 289105 82584 297735
rect 82634 297528 82690 297537
rect 82634 297463 82690 297472
rect 82648 292097 82676 297463
rect 82634 292088 82690 292097
rect 82634 292023 82690 292032
rect 82542 289096 82598 289105
rect 82542 289031 82598 289040
rect 82740 286278 82768 298250
rect 82832 298110 82860 302874
rect 82924 300642 82952 302874
rect 83200 302274 83228 310542
rect 83292 303770 83320 310712
rect 83752 308122 83780 369838
rect 83660 308094 83780 308122
rect 83660 307986 83688 308094
rect 83568 307958 83688 307986
rect 83568 303906 83596 307958
rect 83568 303878 83780 303906
rect 83292 303742 83596 303770
rect 83200 302246 83320 302274
rect 82924 300614 83044 300642
rect 82912 300552 82964 300558
rect 82912 300494 82964 300500
rect 82820 298104 82872 298110
rect 82820 298046 82872 298052
rect 82924 293418 82952 300494
rect 82912 293412 82964 293418
rect 82912 293354 82964 293360
rect 83016 291938 83044 300614
rect 82820 291916 82872 291922
rect 82820 291858 82872 291864
rect 82924 291910 83044 291938
rect 82832 288946 82860 291858
rect 82924 291786 82952 291910
rect 82912 291780 82964 291786
rect 82912 291722 82964 291728
rect 83292 289082 83320 302246
rect 83568 293954 83596 303742
rect 83752 298738 83780 303878
rect 83660 298710 83780 298738
rect 83660 293954 83688 298710
rect 83568 293926 83780 293954
rect 83292 289054 83596 289082
rect 82832 288918 83504 288946
rect 82912 288856 82964 288862
rect 82964 288804 83412 288810
rect 82912 288798 83412 288804
rect 82924 288782 83412 288798
rect 82912 287768 82964 287774
rect 82964 287716 83320 287722
rect 82912 287710 83320 287716
rect 82924 287694 83320 287710
rect 82820 286408 82872 286414
rect 82820 286350 82872 286356
rect 82728 286272 82780 286278
rect 82728 286214 82780 286220
rect 82636 284640 82688 284646
rect 82636 284582 82688 284588
rect 82648 269657 82676 284582
rect 82634 269648 82690 269657
rect 82634 269583 82690 269592
rect 82450 266248 82506 266257
rect 82450 266183 82506 266192
rect 82464 260273 82492 266183
rect 82636 265940 82688 265946
rect 82636 265882 82688 265888
rect 82648 264081 82676 265882
rect 82634 264072 82690 264081
rect 82634 264007 82690 264016
rect 82450 260264 82506 260273
rect 82450 260199 82506 260208
rect 82542 254824 82598 254833
rect 82542 254759 82598 254768
rect 82556 252793 82584 254759
rect 82542 252784 82598 252793
rect 82542 252719 82598 252728
rect 82832 246226 82860 286350
rect 82912 286272 82964 286278
rect 82912 286214 82964 286220
rect 82924 282266 82952 286214
rect 82912 282260 82964 282266
rect 82912 282202 82964 282208
rect 82924 277438 82952 277469
rect 82912 277432 82964 277438
rect 82964 277380 83044 277386
rect 82912 277374 83044 277380
rect 82924 277358 83044 277374
rect 83016 273986 83044 277358
rect 82924 273958 83044 273986
rect 82924 273834 82952 273958
rect 82912 273828 82964 273834
rect 82912 273770 82964 273776
rect 83292 273714 83320 287694
rect 83016 273686 83320 273714
rect 83016 269906 83044 273686
rect 82924 269878 83044 269906
rect 82924 269822 82952 269878
rect 82912 269816 82964 269822
rect 83384 269804 83412 288782
rect 82912 269758 82964 269764
rect 83016 269776 83412 269804
rect 82912 269612 82964 269618
rect 83016 269600 83044 269776
rect 83476 269600 83504 288918
rect 82964 269572 83044 269600
rect 83384 269572 83504 269600
rect 82912 269554 82964 269560
rect 82912 269476 82964 269482
rect 83384 269464 83412 269572
rect 82964 269436 83412 269464
rect 82912 269418 82964 269424
rect 83568 269090 83596 289054
rect 83016 269062 83596 269090
rect 83016 265946 83044 269062
rect 83004 265940 83056 265946
rect 83004 265882 83056 265888
rect 82912 265872 82964 265878
rect 82964 265820 83504 265826
rect 82912 265814 83504 265820
rect 82924 265798 83504 265814
rect 83016 265526 83228 265554
rect 82912 265464 82964 265470
rect 83016 265418 83044 265526
rect 82964 265412 83044 265418
rect 82912 265406 83044 265412
rect 82924 265390 83044 265406
rect 83200 265418 83228 265526
rect 83200 265390 83412 265418
rect 82912 263560 82964 263566
rect 82964 263508 83320 263514
rect 82912 263502 83320 263508
rect 82924 263486 83320 263502
rect 82912 263152 82964 263158
rect 82964 263112 83044 263140
rect 82912 263094 82964 263100
rect 83016 260794 83044 263112
rect 83016 260766 83136 260794
rect 83108 251138 83136 260766
rect 83016 251110 83136 251138
rect 82912 248464 82964 248470
rect 83016 248452 83044 251110
rect 82964 248424 83044 248452
rect 82912 248406 82964 248412
rect 83292 246514 83320 263486
rect 82924 246486 83320 246514
rect 82924 246362 82952 246486
rect 82912 246356 82964 246362
rect 82912 246298 82964 246304
rect 82820 246220 82872 246226
rect 83384 246208 83412 265390
rect 82820 246162 82872 246168
rect 82924 246180 83412 246208
rect 82924 245954 82952 246180
rect 82912 245948 82964 245954
rect 82912 245890 82964 245896
rect 83476 245868 83504 265798
rect 83108 245840 83504 245868
rect 82358 245576 82414 245585
rect 82358 245511 82414 245520
rect 82372 125594 82400 245511
rect 83108 245154 83136 245840
rect 83660 245562 83688 293926
rect 83384 245534 83688 245562
rect 83384 245290 83412 245534
rect 83752 245426 83780 293926
rect 88706 248024 88762 248033
rect 88444 247982 88706 248010
rect 88444 247761 88472 247982
rect 88706 247959 88762 247968
rect 88430 247752 88486 247761
rect 88430 247687 88486 247696
rect 83660 245398 83780 245426
rect 83384 245262 83596 245290
rect 82740 245126 83136 245154
rect 82740 243846 82768 245126
rect 82912 245064 82964 245070
rect 83568 245018 83596 245262
rect 82912 245006 82964 245012
rect 82820 244996 82872 245002
rect 82820 244938 82872 244944
rect 82728 243840 82780 243846
rect 82728 243782 82780 243788
rect 82542 239456 82598 239465
rect 82542 239391 82598 239400
rect 82450 238368 82506 238377
rect 82450 238303 82506 238312
rect 82464 238134 82492 238303
rect 82452 238128 82504 238134
rect 82452 238070 82504 238076
rect 82450 235104 82506 235113
rect 82450 235039 82452 235048
rect 82504 235039 82506 235048
rect 82452 235010 82504 235016
rect 82450 234968 82506 234977
rect 82450 234903 82506 234912
rect 82360 125588 82412 125594
rect 82360 125530 82412 125536
rect 82464 125474 82492 234903
rect 82556 232506 82584 239391
rect 82832 238814 82860 244938
rect 82924 243930 82952 245006
rect 83384 244990 83596 245018
rect 83384 244066 83412 244990
rect 83660 244882 83688 245398
rect 83660 244854 83780 244882
rect 83384 244038 83688 244066
rect 82924 243902 83596 243930
rect 82912 243840 82964 243846
rect 82964 243788 83504 243794
rect 82912 243782 83504 243788
rect 82924 243766 83504 243782
rect 82912 243704 82964 243710
rect 82964 243652 83412 243658
rect 82912 243646 83412 243652
rect 82924 243630 83412 243646
rect 82912 243568 82964 243574
rect 82912 243510 82964 243516
rect 82820 238808 82872 238814
rect 82820 238750 82872 238756
rect 82924 238746 82952 243510
rect 83384 238762 83412 243630
rect 82912 238740 82964 238746
rect 82912 238682 82964 238688
rect 83016 238734 83412 238762
rect 82820 238672 82872 238678
rect 82820 238614 82872 238620
rect 82634 237008 82690 237017
rect 82634 236943 82690 236952
rect 82648 234841 82676 236943
rect 82728 235068 82780 235074
rect 82728 235010 82780 235016
rect 82634 234832 82690 234841
rect 82634 234767 82690 234776
rect 82634 233472 82690 233481
rect 82740 233458 82768 235010
rect 82690 233430 82768 233458
rect 82634 233407 82690 233416
rect 82728 232892 82780 232898
rect 82728 232834 82780 232840
rect 82634 232656 82690 232665
rect 82634 232591 82636 232600
rect 82688 232591 82690 232600
rect 82636 232562 82688 232568
rect 82556 232478 82676 232506
rect 82542 232384 82598 232393
rect 82542 232319 82598 232328
rect 82556 190874 82584 232319
rect 82648 225729 82676 232478
rect 82740 229022 82768 232834
rect 82728 229016 82780 229022
rect 82728 228958 82780 228964
rect 82634 225720 82690 225729
rect 82634 225655 82690 225664
rect 82634 224360 82690 224369
rect 82634 224295 82690 224304
rect 82648 209506 82676 224295
rect 82728 213444 82780 213450
rect 82728 213386 82780 213392
rect 82636 209500 82688 209506
rect 82636 209442 82688 209448
rect 82634 209400 82690 209409
rect 82634 209335 82690 209344
rect 82648 195265 82676 209335
rect 82740 195294 82768 213386
rect 82728 195288 82780 195294
rect 82634 195256 82690 195265
rect 82728 195230 82780 195236
rect 82634 195191 82690 195200
rect 82728 195152 82780 195158
rect 82634 195120 82690 195129
rect 82728 195094 82780 195100
rect 82634 195055 82636 195064
rect 82688 195055 82690 195064
rect 82636 195026 82688 195032
rect 82634 194984 82690 194993
rect 82634 194919 82636 194928
rect 82688 194919 82690 194928
rect 82636 194890 82688 194896
rect 82634 194848 82690 194857
rect 82634 194783 82636 194792
rect 82688 194783 82690 194792
rect 82636 194754 82688 194760
rect 82634 194712 82690 194721
rect 82634 194647 82690 194656
rect 82648 191282 82676 194647
rect 82636 191276 82688 191282
rect 82636 191218 82688 191224
rect 82634 191176 82690 191185
rect 82634 191111 82636 191120
rect 82688 191111 82690 191120
rect 82636 191082 82688 191088
rect 82636 191004 82688 191010
rect 82636 190946 82688 190952
rect 82648 190913 82676 190946
rect 82634 190904 82690 190913
rect 82544 190868 82596 190874
rect 82634 190839 82690 190848
rect 82544 190810 82596 190816
rect 82636 190800 82688 190806
rect 82542 190768 82598 190777
rect 82636 190742 82688 190748
rect 82542 190703 82544 190712
rect 82596 190703 82598 190712
rect 82544 190674 82596 190680
rect 82544 190528 82596 190534
rect 82542 190496 82544 190505
rect 82596 190496 82598 190505
rect 82542 190431 82598 190440
rect 82542 189272 82598 189281
rect 82542 189207 82598 189216
rect 82372 125446 82492 125474
rect 82268 123412 82320 123418
rect 82268 123354 82320 123360
rect 82096 123270 82216 123298
rect 81992 118040 82044 118046
rect 81992 117982 82044 117988
rect 82096 117978 82124 123270
rect 82176 123140 82228 123146
rect 82176 123082 82228 123088
rect 82188 118114 82216 123082
rect 82372 122534 82400 125446
rect 82452 125384 82504 125390
rect 82452 125326 82504 125332
rect 82464 123622 82492 125326
rect 82452 123616 82504 123622
rect 82452 123558 82504 123564
rect 82452 123208 82504 123214
rect 82452 123150 82504 123156
rect 82360 122528 82412 122534
rect 82360 122470 82412 122476
rect 82176 118108 82228 118114
rect 82176 118050 82228 118056
rect 82084 117972 82136 117978
rect 82084 117914 82136 117920
rect 82464 116822 82492 123150
rect 82556 123146 82584 189207
rect 82648 188737 82676 190742
rect 82634 188728 82690 188737
rect 82634 188663 82690 188672
rect 82636 188624 82688 188630
rect 82636 188566 82688 188572
rect 82648 187377 82676 188566
rect 82634 187368 82690 187377
rect 82634 187303 82690 187312
rect 82636 187264 82688 187270
rect 82636 187206 82688 187212
rect 82648 187105 82676 187206
rect 82634 187096 82690 187105
rect 82634 187031 82690 187040
rect 82636 186992 82688 186998
rect 82634 186960 82636 186969
rect 82688 186960 82690 186969
rect 82634 186895 82690 186904
rect 82740 186726 82768 195094
rect 82728 186720 82780 186726
rect 82728 186662 82780 186668
rect 82728 185700 82780 185706
rect 82728 185642 82780 185648
rect 82636 182436 82688 182442
rect 82636 182378 82688 182384
rect 82648 178770 82676 182378
rect 82636 178764 82688 178770
rect 82636 178706 82688 178712
rect 82636 178628 82688 178634
rect 82636 178570 82688 178576
rect 82648 170406 82676 178570
rect 82636 170400 82688 170406
rect 82636 170342 82688 170348
rect 82636 170264 82688 170270
rect 82634 170232 82636 170241
rect 82688 170232 82690 170241
rect 82634 170167 82690 170176
rect 82636 170128 82688 170134
rect 82634 170096 82636 170105
rect 82688 170096 82690 170105
rect 82634 170031 82690 170040
rect 82634 157448 82690 157457
rect 82634 157383 82690 157392
rect 82648 156398 82676 157383
rect 82636 156392 82688 156398
rect 82636 156334 82688 156340
rect 82636 156256 82688 156262
rect 82636 156198 82688 156204
rect 82648 129130 82676 156198
rect 82636 129124 82688 129130
rect 82636 129066 82688 129072
rect 82634 129024 82690 129033
rect 82740 129010 82768 185642
rect 82832 129146 82860 238614
rect 83016 238082 83044 238734
rect 82924 238054 83044 238082
rect 82924 233034 82952 238054
rect 83476 237946 83504 243766
rect 83108 237918 83504 237946
rect 82912 233028 82964 233034
rect 82912 232970 82964 232976
rect 83108 232914 83136 237918
rect 83568 237810 83596 243902
rect 83200 237782 83596 237810
rect 83200 233102 83228 237782
rect 83660 236994 83688 244038
rect 83476 236966 83688 236994
rect 83476 236178 83504 236966
rect 83752 236858 83780 244854
rect 83568 236830 83780 236858
rect 83568 236314 83596 236830
rect 83568 236286 83780 236314
rect 83476 236150 83688 236178
rect 83188 233096 83240 233102
rect 83188 233038 83240 233044
rect 82924 232898 83136 232914
rect 82912 232892 83136 232898
rect 82964 232886 83136 232892
rect 82912 232834 82964 232840
rect 82912 229016 82964 229022
rect 82964 228976 83504 229004
rect 82912 228958 82964 228964
rect 82912 228880 82964 228886
rect 82964 228828 83412 228834
rect 82912 228822 83412 228828
rect 82924 228806 83412 228822
rect 82912 226568 82964 226574
rect 82964 226516 83320 226522
rect 82912 226510 83320 226516
rect 82924 226494 83320 226510
rect 82912 225684 82964 225690
rect 82964 225644 83228 225672
rect 82912 225626 82964 225632
rect 82924 220918 83044 220946
rect 82924 220862 82952 220918
rect 82912 220856 82964 220862
rect 82912 220798 82964 220804
rect 83016 220810 83044 220918
rect 83200 220810 83228 225644
rect 83016 220782 83228 220810
rect 82912 219496 82964 219502
rect 82912 219438 82964 219444
rect 82924 211206 82952 219438
rect 82912 211200 82964 211206
rect 82912 211142 82964 211148
rect 83004 211200 83056 211206
rect 83004 211142 83056 211148
rect 83016 195378 83044 211142
rect 82924 195362 83044 195378
rect 82912 195356 83044 195362
rect 82964 195350 83044 195356
rect 82912 195298 82964 195304
rect 83292 195242 83320 226494
rect 82924 195226 83320 195242
rect 82912 195220 83320 195226
rect 82964 195214 83320 195220
rect 82912 195162 82964 195168
rect 83384 194970 83412 228806
rect 82924 194954 83412 194970
rect 82912 194948 83412 194954
rect 82964 194942 83412 194948
rect 82912 194890 82964 194896
rect 83476 194834 83504 228976
rect 82924 194818 83504 194834
rect 82912 194812 83504 194818
rect 82964 194806 83504 194812
rect 82912 194754 82964 194760
rect 82912 192228 82964 192234
rect 82912 192170 82964 192176
rect 82924 188306 82952 192170
rect 82924 188278 83596 188306
rect 82912 186992 82964 186998
rect 82964 186940 83044 186946
rect 82912 186934 83044 186940
rect 82924 186918 83044 186934
rect 82912 186720 82964 186726
rect 82912 186662 82964 186668
rect 82924 177274 82952 186662
rect 83016 184226 83044 186918
rect 83016 184198 83228 184226
rect 82912 177268 82964 177274
rect 82912 177210 82964 177216
rect 83200 177154 83228 184198
rect 82924 177138 83228 177154
rect 82912 177132 83228 177138
rect 82964 177126 83228 177132
rect 82912 177074 82964 177080
rect 82912 176996 82964 177002
rect 82964 176956 83504 176984
rect 82912 176938 82964 176944
rect 82912 176656 82964 176662
rect 82964 176616 83412 176644
rect 82912 176598 82964 176604
rect 82912 173188 82964 173194
rect 82912 173130 82964 173136
rect 82924 157622 82952 173130
rect 83004 168428 83056 168434
rect 83384 168416 83412 176616
rect 83056 168388 83412 168416
rect 83004 168370 83056 168376
rect 83476 167770 83504 176956
rect 83016 167742 83504 167770
rect 83016 167278 83044 167742
rect 83004 167272 83056 167278
rect 83004 167214 83056 167220
rect 83004 167136 83056 167142
rect 83004 167078 83056 167084
rect 83016 166954 83044 167078
rect 83016 166926 83320 166954
rect 83004 166728 83056 166734
rect 83056 166676 83228 166682
rect 83004 166670 83228 166676
rect 83016 166654 83228 166670
rect 83004 166048 83056 166054
rect 83004 165990 83056 165996
rect 82912 157616 82964 157622
rect 82912 157558 82964 157564
rect 83016 157554 83044 165990
rect 83200 157706 83228 166654
rect 83292 162874 83320 166926
rect 83292 162846 83412 162874
rect 83108 157678 83228 157706
rect 83004 157548 83056 157554
rect 83004 157490 83056 157496
rect 83108 157434 83136 157678
rect 83384 157570 83412 162846
rect 83384 157542 83504 157570
rect 83016 157406 83136 157434
rect 83016 157332 83044 157406
rect 82924 157304 83044 157332
rect 82924 157010 82952 157304
rect 83476 157162 83504 157542
rect 83292 157134 83504 157162
rect 83004 157072 83056 157078
rect 83292 157026 83320 157134
rect 83056 157020 83320 157026
rect 83004 157014 83320 157020
rect 82912 157004 82964 157010
rect 83016 156998 83320 157014
rect 82912 156946 82964 156952
rect 82912 156868 82964 156874
rect 82912 156810 82964 156816
rect 82924 156482 82952 156810
rect 83004 156800 83056 156806
rect 83004 156742 83056 156748
rect 83016 156618 83044 156742
rect 83016 156590 83504 156618
rect 82924 156454 83320 156482
rect 82912 156392 82964 156398
rect 82912 156334 82964 156340
rect 82924 152522 82952 156334
rect 82912 152516 82964 152522
rect 82912 152458 82964 152464
rect 82924 152386 83228 152402
rect 82912 152380 83228 152386
rect 82964 152374 83228 152380
rect 82912 152322 82964 152328
rect 82912 152176 82964 152182
rect 82964 152124 83044 152130
rect 82912 152118 83044 152124
rect 82924 152102 83044 152118
rect 83016 146010 83044 152102
rect 82924 145982 83044 146010
rect 82924 145926 82952 145982
rect 82912 145920 82964 145926
rect 82912 145862 82964 145868
rect 82912 145784 82964 145790
rect 82912 145726 82964 145732
rect 82924 145602 82952 145726
rect 82924 145574 83044 145602
rect 82912 145512 82964 145518
rect 82912 145454 82964 145460
rect 82924 138718 82952 145454
rect 82912 138712 82964 138718
rect 82912 138654 82964 138660
rect 83016 138530 83044 145574
rect 82924 138514 83044 138530
rect 82912 138508 83044 138514
rect 82964 138502 83044 138508
rect 82912 138450 82964 138456
rect 82912 137352 82964 137358
rect 83200 137340 83228 152374
rect 83292 151858 83320 156454
rect 83292 151830 83412 151858
rect 83384 147642 83412 151830
rect 82964 137312 83228 137340
rect 83292 147614 83412 147642
rect 82912 137294 82964 137300
rect 83292 137272 83320 147614
rect 83016 137244 83320 137272
rect 82912 137216 82964 137222
rect 83016 137204 83044 137244
rect 82964 137176 83044 137204
rect 82912 137158 82964 137164
rect 82912 137080 82964 137086
rect 82964 137040 83320 137068
rect 82912 137022 82964 137028
rect 82912 136944 82964 136950
rect 82964 136892 83228 136898
rect 82912 136886 83228 136892
rect 82924 136870 83228 136886
rect 82912 136672 82964 136678
rect 82912 136614 82964 136620
rect 82924 133906 82952 136614
rect 82924 133878 83044 133906
rect 83016 133210 83044 133878
rect 83004 133204 83056 133210
rect 83004 133146 83056 133152
rect 82924 133074 83136 133090
rect 82912 133068 83136 133074
rect 82964 133062 83136 133068
rect 82912 133010 82964 133016
rect 82912 132320 82964 132326
rect 82912 132262 82964 132268
rect 82924 129282 82952 132262
rect 82924 129254 83044 129282
rect 82832 129118 82952 129146
rect 82740 128982 82860 129010
rect 82634 128959 82690 128968
rect 82544 123140 82596 123146
rect 82544 123082 82596 123088
rect 82648 122913 82676 128959
rect 82728 128920 82780 128926
rect 82728 128862 82780 128868
rect 82634 122904 82690 122913
rect 82634 122839 82690 122848
rect 82556 118182 82584 122060
rect 82740 119474 82768 128862
rect 82832 122194 82860 128982
rect 82924 123690 82952 129118
rect 83016 123865 83044 129254
rect 83002 123856 83058 123865
rect 83002 123791 83058 123800
rect 83108 123729 83136 133062
rect 83094 123720 83150 123729
rect 82912 123684 82964 123690
rect 83094 123655 83150 123664
rect 82912 123626 82964 123632
rect 83200 123604 83228 136870
rect 83108 123576 83228 123604
rect 82820 122188 82872 122194
rect 82820 122130 82872 122136
rect 82728 119468 82780 119474
rect 82728 119410 82780 119416
rect 83108 118386 83136 123576
rect 83292 118522 83320 137040
rect 83370 123856 83426 123865
rect 83370 123791 83426 123800
rect 83280 118516 83332 118522
rect 83280 118458 83332 118464
rect 83096 118380 83148 118386
rect 83096 118322 83148 118328
rect 82544 118176 82596 118182
rect 82544 118118 82596 118124
rect 83186 118008 83242 118017
rect 83186 117943 83242 117952
rect 82452 116816 82504 116822
rect 82452 116758 82504 116764
rect 82728 113212 82780 113218
rect 82728 113154 82780 113160
rect 82740 111790 82768 113154
rect 82636 111784 82688 111790
rect 82636 111726 82688 111732
rect 82728 111784 82780 111790
rect 82728 111726 82780 111732
rect 82648 102218 82676 111726
rect 83200 106321 83228 117943
rect 83384 111790 83412 123791
rect 83476 122738 83504 156590
rect 83568 123865 83596 188278
rect 83554 123856 83610 123865
rect 83554 123791 83610 123800
rect 83660 123706 83688 236150
rect 83568 123678 83688 123706
rect 83464 122732 83516 122738
rect 83464 122674 83516 122680
rect 83568 122466 83596 123678
rect 83646 123312 83702 123321
rect 83646 123247 83702 123256
rect 83556 122460 83608 122466
rect 83556 122402 83608 122408
rect 83660 119270 83688 123247
rect 83648 119264 83700 119270
rect 83648 119206 83700 119212
rect 83752 111790 83780 236286
rect 88706 233064 88762 233073
rect 87892 233022 88706 233050
rect 87892 232801 87920 233022
rect 88706 232999 88762 233008
rect 87878 232792 87934 232801
rect 87878 232727 87934 232736
rect 84566 226808 84622 226817
rect 86130 226808 86186 226817
rect 84622 226766 86130 226794
rect 84566 226743 84622 226752
rect 86130 226743 86186 226752
rect 87326 179888 87382 179897
rect 88706 179888 88762 179897
rect 87382 179846 88706 179874
rect 87326 179823 87382 179832
rect 88706 179823 88762 179832
rect 87326 171592 87382 171601
rect 87602 171592 87658 171601
rect 87382 171550 87602 171578
rect 87326 171527 87382 171536
rect 87602 171527 87658 171536
rect 501524 151978 501552 584258
rect 501616 157622 501644 700674
rect 502524 700664 502576 700670
rect 502524 700606 502576 700612
rect 501788 700596 501840 700602
rect 501788 700538 501840 700544
rect 501696 581120 501748 581126
rect 501696 581062 501748 581068
rect 501708 159118 501736 581062
rect 501800 518129 501828 700538
rect 502340 583840 502392 583846
rect 502340 583782 502392 583788
rect 501972 582820 502024 582826
rect 501972 582762 502024 582768
rect 501880 582004 501932 582010
rect 501880 581946 501932 581952
rect 501892 581126 501920 581946
rect 501880 581120 501932 581126
rect 501880 581062 501932 581068
rect 501880 580984 501932 580990
rect 501880 580926 501932 580932
rect 501786 518120 501842 518129
rect 501786 518055 501842 518064
rect 501786 517304 501842 517313
rect 501786 517239 501842 517248
rect 501800 506977 501828 517239
rect 501786 506968 501842 506977
rect 501786 506903 501842 506912
rect 501786 474872 501842 474881
rect 501786 474807 501842 474816
rect 501800 464273 501828 474807
rect 501786 464264 501842 464273
rect 501786 464199 501842 464208
rect 501786 457192 501842 457201
rect 501786 457127 501842 457136
rect 501696 159112 501748 159118
rect 501696 159054 501748 159060
rect 501694 158944 501750 158953
rect 501694 158879 501750 158888
rect 501604 157616 501656 157622
rect 501604 157558 501656 157564
rect 501604 157480 501656 157486
rect 501602 157448 501604 157457
rect 501656 157448 501658 157457
rect 501602 157383 501658 157392
rect 501708 156641 501736 158879
rect 501694 156632 501750 156641
rect 501694 156567 501750 156576
rect 501604 154896 501656 154902
rect 501604 154838 501656 154844
rect 501512 151972 501564 151978
rect 501512 151914 501564 151920
rect 501510 151872 501566 151881
rect 501510 151807 501512 151816
rect 501564 151807 501566 151816
rect 501512 151778 501564 151784
rect 501512 151700 501564 151706
rect 501512 151642 501564 151648
rect 501524 124778 501552 151642
rect 501616 127362 501644 154838
rect 501696 154760 501748 154766
rect 501694 154728 501696 154737
rect 501748 154728 501750 154737
rect 501694 154663 501750 154672
rect 501696 154624 501748 154630
rect 501696 154566 501748 154572
rect 501708 136377 501736 154566
rect 501694 136368 501750 136377
rect 501694 136303 501750 136312
rect 501696 136196 501748 136202
rect 501696 136138 501748 136144
rect 501708 133346 501736 136138
rect 501696 133340 501748 133346
rect 501696 133282 501748 133288
rect 501696 133204 501748 133210
rect 501696 133146 501748 133152
rect 501604 127356 501656 127362
rect 501604 127298 501656 127304
rect 501602 126168 501658 126177
rect 501602 126103 501658 126112
rect 501512 124772 501564 124778
rect 501512 124714 501564 124720
rect 501512 124636 501564 124642
rect 501512 124578 501564 124584
rect 120540 122732 120592 122738
rect 120540 122674 120592 122680
rect 124312 122732 124364 122738
rect 124312 122674 124364 122680
rect 133788 122732 133840 122738
rect 133788 122674 133840 122680
rect 286968 122732 287020 122738
rect 286968 122674 287020 122680
rect 500144 122726 500540 122754
rect 87510 122632 87566 122641
rect 87170 122590 87510 122618
rect 87510 122567 87566 122576
rect 88982 122632 89038 122641
rect 88982 122567 89038 122576
rect 89258 122632 89314 122641
rect 89258 122567 89314 122576
rect 90638 122632 90694 122641
rect 90638 122567 90694 122576
rect 92294 122632 92350 122641
rect 92294 122567 92350 122576
rect 101034 122632 101090 122641
rect 101034 122567 101090 122576
rect 86866 122360 86922 122369
rect 86866 122295 86922 122304
rect 83830 122224 83886 122233
rect 83830 122159 83886 122168
rect 83844 116754 83872 122159
rect 84106 120728 84162 120737
rect 84106 120663 84162 120672
rect 84016 120624 84068 120630
rect 84016 120566 84068 120572
rect 83832 116748 83884 116754
rect 83832 116690 83884 116696
rect 83372 111784 83424 111790
rect 83372 111726 83424 111732
rect 83740 111784 83792 111790
rect 83740 111726 83792 111732
rect 83832 111784 83884 111790
rect 83832 111726 83884 111732
rect 83464 111716 83516 111722
rect 83464 111658 83516 111664
rect 83186 106312 83242 106321
rect 83186 106247 83242 106256
rect 83278 104816 83334 104825
rect 83278 104751 83334 104760
rect 82648 102190 82768 102218
rect 82740 53802 82768 102190
rect 83292 95305 83320 104751
rect 83278 95296 83334 95305
rect 83278 95231 83334 95240
rect 83278 86864 83334 86873
rect 83278 86799 83334 86808
rect 83292 77353 83320 86799
rect 83278 77344 83334 77353
rect 83278 77279 83334 77288
rect 83278 77072 83334 77081
rect 83278 77007 83334 77016
rect 83292 67697 83320 77007
rect 83278 67688 83334 67697
rect 83278 67623 83334 67632
rect 83278 57896 83334 57905
rect 83278 57831 83334 57840
rect 82648 53774 82768 53802
rect 82648 45626 82676 53774
rect 83292 48385 83320 57831
rect 83278 48376 83334 48385
rect 83278 48311 83334 48320
rect 82636 45620 82688 45626
rect 82636 45562 82688 45568
rect 83476 44198 83504 111658
rect 82636 44192 82688 44198
rect 82636 44134 82688 44140
rect 83372 44192 83424 44198
rect 83372 44134 83424 44140
rect 83464 44192 83516 44198
rect 83844 44180 83872 111726
rect 83464 44134 83516 44140
rect 83752 44152 83872 44180
rect 82648 29730 82676 44134
rect 83278 38584 83334 38593
rect 83278 38519 83334 38528
rect 82648 29702 82768 29730
rect 82740 13977 82768 29702
rect 83292 29209 83320 38519
rect 83384 35850 83412 44134
rect 83752 35902 83780 44152
rect 83740 35896 83792 35902
rect 83384 35822 83504 35850
rect 83740 35838 83792 35844
rect 83832 35896 83884 35902
rect 83832 35838 83884 35844
rect 83278 29200 83334 29209
rect 83278 29135 83334 29144
rect 83278 19136 83334 19145
rect 83278 19071 83334 19080
rect 83292 15881 83320 19071
rect 83278 15872 83334 15881
rect 83278 15807 83334 15816
rect 82726 13968 82782 13977
rect 82726 13903 82782 13912
rect 82634 13832 82690 13841
rect 82634 13767 82690 13776
rect 82648 6934 82676 13767
rect 83476 9246 83504 35822
rect 83844 9450 83872 35838
rect 83922 16008 83978 16017
rect 83922 15943 83978 15952
rect 83832 9444 83884 9450
rect 83832 9386 83884 9392
rect 83464 9240 83516 9246
rect 83464 9182 83516 9188
rect 83936 7562 83964 15943
rect 84028 11762 84056 120566
rect 84016 11756 84068 11762
rect 84016 11698 84068 11704
rect 84120 10606 84148 120663
rect 84764 120018 84792 122060
rect 86880 121990 86908 122295
rect 86868 121984 86920 121990
rect 86868 121926 86920 121932
rect 84936 121848 84988 121854
rect 88996 121825 89024 122567
rect 84936 121790 84988 121796
rect 88982 121816 89038 121825
rect 84752 120012 84804 120018
rect 84752 119954 84804 119960
rect 84844 118176 84896 118182
rect 84844 118118 84896 118124
rect 84290 106992 84346 107001
rect 84290 106927 84346 106936
rect 84304 98705 84332 106927
rect 84290 98696 84346 98705
rect 84290 98631 84346 98640
rect 84382 86320 84438 86329
rect 84382 86255 84438 86264
rect 84396 78033 84424 86255
rect 84382 78024 84438 78033
rect 84382 77959 84438 77968
rect 84382 23352 84438 23361
rect 84382 23287 84438 23296
rect 84396 13841 84424 23287
rect 84382 13832 84438 13841
rect 84382 13767 84438 13776
rect 84382 13696 84438 13705
rect 84382 13631 84438 13640
rect 84108 10600 84160 10606
rect 84108 10542 84160 10548
rect 83844 7534 83964 7562
rect 82636 6928 82688 6934
rect 82636 6870 82688 6876
rect 82544 6724 82596 6730
rect 82544 6666 82596 6672
rect 81900 4820 81952 4826
rect 81900 4762 81952 4768
rect 81438 3904 81494 3913
rect 80428 3868 80480 3874
rect 81438 3839 81494 3848
rect 80428 3810 80480 3816
rect 80244 604 80296 610
rect 80244 546 80296 552
rect 80336 604 80388 610
rect 80336 546 80388 552
rect 80256 480 80284 546
rect 81452 480 81480 3839
rect 82556 3505 82584 6666
rect 82634 5400 82690 5409
rect 82634 5335 82690 5344
rect 82542 3496 82598 3505
rect 82542 3431 82598 3440
rect 82648 480 82676 5335
rect 83844 480 83872 7534
rect 84396 4185 84424 13631
rect 84856 4962 84884 118118
rect 84948 7698 84976 121790
rect 88982 121751 89038 121760
rect 85028 121100 85080 121106
rect 85028 121042 85080 121048
rect 85040 7834 85068 121042
rect 88430 120728 88486 120737
rect 88430 120663 88486 120672
rect 87328 119264 87380 119270
rect 87328 119206 87380 119212
rect 86038 116920 86094 116929
rect 86038 116855 86094 116864
rect 85488 109744 85540 109750
rect 85488 109686 85540 109692
rect 85040 7806 85160 7834
rect 84948 7670 85068 7698
rect 84844 4956 84896 4962
rect 84844 4898 84896 4904
rect 84382 4176 84438 4185
rect 84382 4111 84438 4120
rect 84936 4140 84988 4146
rect 84936 4082 84988 4088
rect 84948 480 84976 4082
rect 85040 3126 85068 7670
rect 85028 3120 85080 3126
rect 85028 3062 85080 3068
rect 85132 2922 85160 7806
rect 85500 4146 85528 109686
rect 86052 106457 86080 116855
rect 87340 116793 87368 119206
rect 87142 116784 87198 116793
rect 87142 116719 87198 116728
rect 87326 116784 87382 116793
rect 87326 116719 87382 116728
rect 86590 111208 86646 111217
rect 86590 111143 86646 111152
rect 86604 107001 86632 111143
rect 86590 106992 86646 107001
rect 86590 106927 86646 106936
rect 86038 106448 86094 106457
rect 86038 106383 86094 106392
rect 87156 105913 87184 116719
rect 88444 106321 88472 120663
rect 89272 120057 89300 122567
rect 89258 120048 89314 120057
rect 89258 119983 89314 119992
rect 89548 113150 89576 122060
rect 90652 121854 90680 122567
rect 90640 121848 90692 121854
rect 90640 121790 90692 121796
rect 91940 119406 91968 122060
rect 92308 121786 92336 122567
rect 95330 122224 95386 122233
rect 95160 122182 95280 122210
rect 92296 121780 92348 121786
rect 92296 121722 92348 121728
rect 94332 119406 94360 122060
rect 95160 121990 95188 122182
rect 95148 121984 95200 121990
rect 95148 121926 95200 121932
rect 95252 121922 95280 122182
rect 95330 122159 95386 122168
rect 95344 121990 95372 122159
rect 95332 121984 95384 121990
rect 95332 121926 95384 121932
rect 95240 121916 95292 121922
rect 95240 121858 95292 121864
rect 91928 119400 91980 119406
rect 91928 119342 91980 119348
rect 94320 119400 94372 119406
rect 96724 119377 96752 122060
rect 99130 122046 99328 122074
rect 94320 119342 94372 119348
rect 96710 119368 96766 119377
rect 96710 119303 96766 119312
rect 92388 119196 92440 119202
rect 92388 119138 92440 119144
rect 91008 119128 91060 119134
rect 91008 119070 91060 119076
rect 89536 113144 89588 113150
rect 89536 113086 89588 113092
rect 89628 113076 89680 113082
rect 89628 113018 89680 113024
rect 88246 106312 88302 106321
rect 88246 106247 88302 106256
rect 88430 106312 88486 106321
rect 88430 106247 88486 106256
rect 87142 105904 87198 105913
rect 87142 105839 87198 105848
rect 88260 101561 88288 106247
rect 88246 101552 88302 101561
rect 88246 101487 88302 101496
rect 88154 96520 88210 96529
rect 88154 96455 88210 96464
rect 87970 96384 88026 96393
rect 87970 96319 88026 96328
rect 87984 92721 88012 96319
rect 88168 94625 88196 96455
rect 88154 94616 88210 94625
rect 88154 94551 88210 94560
rect 87970 92712 88026 92721
rect 87970 92647 88026 92656
rect 87142 86320 87198 86329
rect 87142 86255 87198 86264
rect 87156 78033 87184 86255
rect 87142 78024 87198 78033
rect 87142 77959 87198 77968
rect 87602 78024 87658 78033
rect 87602 77959 87658 77968
rect 88246 78024 88302 78033
rect 88246 77959 88302 77968
rect 87616 67697 87644 77959
rect 88260 69193 88288 77959
rect 88246 69184 88302 69193
rect 88246 69119 88302 69128
rect 87602 67688 87658 67697
rect 87602 67623 87658 67632
rect 85762 62792 85818 62801
rect 85762 62727 85818 62736
rect 85776 48521 85804 62727
rect 87510 57896 87566 57905
rect 87510 57831 87566 57840
rect 85762 48512 85818 48521
rect 85762 48447 85818 48456
rect 87524 48385 87552 57831
rect 87510 48376 87566 48385
rect 87510 48311 87566 48320
rect 89640 44282 89668 113018
rect 89640 44254 89760 44282
rect 89732 44180 89760 44254
rect 89640 44152 89760 44180
rect 85854 43480 85910 43489
rect 85854 43415 85910 43424
rect 85868 37505 85896 43415
rect 88248 37936 88300 37942
rect 88248 37878 88300 37884
rect 85854 37496 85910 37505
rect 85854 37431 85910 37440
rect 87510 35320 87566 35329
rect 87510 35255 87566 35264
rect 85854 27568 85910 27577
rect 85854 27503 85910 27512
rect 85868 18193 85896 27503
rect 87524 23497 87552 35255
rect 87510 23488 87566 23497
rect 87510 23423 87566 23432
rect 86406 22808 86462 22817
rect 86406 22743 86462 22752
rect 85946 19272 86002 19281
rect 85946 19207 86002 19216
rect 85854 18184 85910 18193
rect 85854 18119 85910 18128
rect 85960 9897 85988 19207
rect 85946 9888 86002 9897
rect 85946 9823 86002 9832
rect 86222 9480 86278 9489
rect 86222 9415 86278 9424
rect 86130 4720 86186 4729
rect 86130 4655 86186 4664
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 85578 3496 85634 3505
rect 85578 3431 85634 3440
rect 85120 2916 85172 2922
rect 85120 2858 85172 2864
rect 85592 2786 85620 3431
rect 85580 2780 85632 2786
rect 85580 2722 85632 2728
rect 86144 480 86172 4655
rect 86236 3233 86264 9415
rect 86420 4185 86448 22743
rect 87786 8120 87842 8129
rect 87786 8055 87842 8064
rect 87800 5817 87828 8055
rect 87786 5808 87842 5817
rect 87786 5743 87842 5752
rect 86406 4176 86462 4185
rect 88260 4146 88288 37878
rect 89640 22250 89668 44152
rect 89640 22222 89760 22250
rect 89732 13818 89760 22222
rect 89548 13790 89760 13818
rect 89548 9042 89576 13790
rect 89536 9036 89588 9042
rect 89536 8978 89588 8984
rect 86406 4111 86462 4120
rect 87328 4140 87380 4146
rect 87328 4082 87380 4088
rect 88248 4140 88300 4146
rect 88248 4082 88300 4088
rect 86222 3224 86278 3233
rect 86222 3159 86278 3168
rect 87340 480 87368 4082
rect 88522 3904 88578 3913
rect 88522 3839 88578 3848
rect 90730 3904 90786 3913
rect 90730 3839 90786 3848
rect 90914 3904 90970 3913
rect 90914 3839 90970 3848
rect 88536 480 88564 3839
rect 89720 3732 89772 3738
rect 89720 3674 89772 3680
rect 89732 480 89760 3674
rect 90744 3505 90772 3839
rect 90730 3496 90786 3505
rect 90730 3431 90786 3440
rect 90928 480 90956 3839
rect 91020 3738 91048 119070
rect 91008 3732 91060 3738
rect 91008 3674 91060 3680
rect 92400 610 92428 119138
rect 99196 17400 99248 17406
rect 99196 17342 99248 17348
rect 96528 17332 96580 17338
rect 96528 17274 96580 17280
rect 96540 4146 96568 17274
rect 99102 16144 99158 16153
rect 99102 16079 99158 16088
rect 99012 12436 99064 12442
rect 99012 12378 99064 12384
rect 95700 4140 95752 4146
rect 95700 4082 95752 4088
rect 96528 4140 96580 4146
rect 96528 4082 96580 4088
rect 98092 4140 98144 4146
rect 98092 4082 98144 4088
rect 93308 3732 93360 3738
rect 93308 3674 93360 3680
rect 92112 604 92164 610
rect 92112 546 92164 552
rect 92388 604 92440 610
rect 92388 546 92440 552
rect 92124 480 92152 546
rect 93320 480 93348 3674
rect 95146 3632 95202 3641
rect 95146 3567 95202 3576
rect 94502 2952 94558 2961
rect 94502 2887 94558 2896
rect 94516 480 94544 2887
rect 95160 2786 95188 3567
rect 95148 2780 95200 2786
rect 95148 2722 95200 2728
rect 95712 480 95740 4082
rect 96896 2780 96948 2786
rect 96896 2722 96948 2728
rect 96908 480 96936 2722
rect 98104 480 98132 4082
rect 99024 4026 99052 12378
rect 99116 4146 99144 16079
rect 99208 12442 99236 17342
rect 99196 12436 99248 12442
rect 99196 12378 99248 12384
rect 99300 6458 99328 122046
rect 99380 122052 99432 122058
rect 99380 121994 99432 122000
rect 99392 12424 99420 121994
rect 101048 121990 101076 122567
rect 101522 122046 101996 122074
rect 101036 121984 101088 121990
rect 101036 121926 101088 121932
rect 99392 12396 99512 12424
rect 99484 9654 99512 12396
rect 99472 9648 99524 9654
rect 99472 9590 99524 9596
rect 99288 6452 99340 6458
rect 99288 6394 99340 6400
rect 101968 4894 101996 122046
rect 103520 122052 103572 122058
rect 103520 121994 103572 122000
rect 102048 119264 102100 119270
rect 102048 119206 102100 119212
rect 101956 4888 102008 4894
rect 101956 4830 102008 4836
rect 99104 4140 99156 4146
rect 99104 4082 99156 4088
rect 99024 3998 99328 4026
rect 99300 480 99328 3998
rect 102060 3738 102088 119206
rect 102784 8016 102836 8022
rect 102784 7958 102836 7964
rect 101588 3732 101640 3738
rect 101588 3674 101640 3680
rect 102048 3732 102100 3738
rect 102048 3674 102100 3680
rect 99380 2984 99432 2990
rect 99380 2926 99432 2932
rect 99392 2825 99420 2926
rect 99378 2816 99434 2825
rect 99378 2751 99434 2760
rect 100484 604 100536 610
rect 100484 546 100536 552
rect 100496 480 100524 546
rect 101600 480 101628 3674
rect 102796 480 102824 7958
rect 103532 3738 103560 121994
rect 103900 119610 103928 122060
rect 105360 121916 105412 121922
rect 105360 121858 105412 121864
rect 105372 121145 105400 121858
rect 105358 121136 105414 121145
rect 105358 121071 105414 121080
rect 106292 119610 106320 122060
rect 108698 122046 108988 122074
rect 106464 120488 106516 120494
rect 106464 120430 106516 120436
rect 103888 119604 103940 119610
rect 103888 119546 103940 119552
rect 104808 119604 104860 119610
rect 104808 119546 104860 119552
rect 106280 119604 106332 119610
rect 106280 119546 106332 119552
rect 104820 11830 104848 119546
rect 106188 118992 106240 118998
rect 106188 118934 106240 118940
rect 104808 11824 104860 11830
rect 104808 11766 104860 11772
rect 106200 3738 106228 118934
rect 106476 12442 106504 120430
rect 107476 119604 107528 119610
rect 107476 119546 107528 119552
rect 106464 12436 106516 12442
rect 106464 12378 106516 12384
rect 107384 12436 107436 12442
rect 107384 12378 107436 12384
rect 103520 3732 103572 3738
rect 103520 3674 103572 3680
rect 103980 3732 104032 3738
rect 103980 3674 104032 3680
rect 105176 3732 105228 3738
rect 105176 3674 105228 3680
rect 106188 3732 106240 3738
rect 106188 3674 106240 3680
rect 106372 3732 106424 3738
rect 106372 3674 106424 3680
rect 103992 480 104020 3674
rect 105188 480 105216 3674
rect 106384 480 106412 3674
rect 107396 2938 107424 12378
rect 107488 5166 107516 119546
rect 107568 118788 107620 118794
rect 107568 118730 107620 118736
rect 107476 5160 107528 5166
rect 107476 5102 107528 5108
rect 107580 3738 107608 118730
rect 108960 8974 108988 122046
rect 111076 121718 111104 122060
rect 111064 121712 111116 121718
rect 111064 121654 111116 121660
rect 113468 119270 113496 122060
rect 113456 119264 113508 119270
rect 113456 119206 113508 119212
rect 114468 119264 114520 119270
rect 114468 119206 114520 119212
rect 113088 118856 113140 118862
rect 113088 118798 113140 118804
rect 110420 114572 110472 114578
rect 110420 114514 110472 114520
rect 110432 114442 110460 114514
rect 110420 114436 110472 114442
rect 110420 114378 110472 114384
rect 110328 112464 110380 112470
rect 110328 112406 110380 112412
rect 110340 13122 110368 112406
rect 110420 104916 110472 104922
rect 110420 104858 110472 104864
rect 110432 95418 110460 104858
rect 110432 95390 110552 95418
rect 110524 95282 110552 95390
rect 110432 95254 110552 95282
rect 110432 95198 110460 95254
rect 110420 95192 110472 95198
rect 110420 95134 110472 95140
rect 110420 85672 110472 85678
rect 110420 85614 110472 85620
rect 110432 85542 110460 85614
rect 110420 85536 110472 85542
rect 110420 85478 110472 85484
rect 110512 85536 110564 85542
rect 110512 85478 110564 85484
rect 110524 75970 110552 85478
rect 110432 75942 110552 75970
rect 110432 75886 110460 75942
rect 110420 75880 110472 75886
rect 110420 75822 110472 75828
rect 110420 66292 110472 66298
rect 110420 66234 110472 66240
rect 110432 56778 110460 66234
rect 110420 56772 110472 56778
rect 110420 56714 110472 56720
rect 110420 56636 110472 56642
rect 110420 56578 110472 56584
rect 110432 56506 110460 56578
rect 110420 56500 110472 56506
rect 110420 56442 110472 56448
rect 110420 46980 110472 46986
rect 110420 46922 110472 46928
rect 110432 37466 110460 46922
rect 110420 37460 110472 37466
rect 110420 37402 110472 37408
rect 110420 37324 110472 37330
rect 110420 37266 110472 37272
rect 110432 37194 110460 37266
rect 110420 37188 110472 37194
rect 110420 37130 110472 37136
rect 110420 27668 110472 27674
rect 110420 27610 110472 27616
rect 110432 18154 110460 27610
rect 110420 18148 110472 18154
rect 110420 18090 110472 18096
rect 110420 18012 110472 18018
rect 110420 17954 110472 17960
rect 110432 17898 110460 17954
rect 110432 17870 110552 17898
rect 109960 13116 110012 13122
rect 109960 13058 110012 13064
rect 110328 13116 110380 13122
rect 110328 13058 110380 13064
rect 108948 8968 109000 8974
rect 108948 8910 109000 8916
rect 107568 3732 107620 3738
rect 107568 3674 107620 3680
rect 107580 3182 108896 3210
rect 107580 3097 107608 3182
rect 107566 3088 107622 3097
rect 107566 3023 107622 3032
rect 108762 3088 108818 3097
rect 108868 3074 108896 3182
rect 108946 3088 109002 3097
rect 108868 3046 108946 3074
rect 108762 3023 108818 3032
rect 108946 3023 109002 3032
rect 107396 2910 107608 2938
rect 107580 480 107608 2910
rect 108776 480 108804 3023
rect 108948 2984 109000 2990
rect 108948 2926 109000 2932
rect 108960 2825 108988 2926
rect 108946 2816 109002 2825
rect 108946 2751 109002 2760
rect 109972 480 110000 13058
rect 110524 8378 110552 17870
rect 110432 8350 110552 8378
rect 110432 6866 110460 8350
rect 110420 6860 110472 6866
rect 110420 6802 110472 6808
rect 113100 3738 113128 118798
rect 113548 8152 113600 8158
rect 113548 8094 113600 8100
rect 112352 3732 112404 3738
rect 112352 3674 112404 3680
rect 113088 3732 113140 3738
rect 113088 3674 113140 3680
rect 111156 604 111208 610
rect 111156 546 111208 552
rect 111168 480 111196 546
rect 112364 480 112392 3674
rect 113560 480 113588 8094
rect 114480 5098 114508 119206
rect 115860 10538 115888 122060
rect 118266 122046 118648 122074
rect 117778 121544 117834 121553
rect 117778 121479 117834 121488
rect 117792 115818 117820 121479
rect 118424 120624 118476 120630
rect 118424 120566 118476 120572
rect 118436 115977 118464 120566
rect 118422 115968 118478 115977
rect 118422 115903 118478 115912
rect 117700 115790 117820 115818
rect 117700 110430 117728 115790
rect 117688 110424 117740 110430
rect 117688 110366 117740 110372
rect 117504 100836 117556 100842
rect 117504 100778 117556 100784
rect 117516 100706 117544 100778
rect 117504 100700 117556 100706
rect 117504 100642 117556 100648
rect 117780 100700 117832 100706
rect 117780 100642 117832 100648
rect 117792 99346 117820 100642
rect 117780 99340 117832 99346
rect 117780 99282 117832 99288
rect 117504 89752 117556 89758
rect 117504 89694 117556 89700
rect 117516 81462 117544 89694
rect 117504 81456 117556 81462
rect 117504 81398 117556 81404
rect 117596 81456 117648 81462
rect 117596 81398 117648 81404
rect 117608 80170 117636 81398
rect 117596 80164 117648 80170
rect 117596 80106 117648 80112
rect 117504 80028 117556 80034
rect 117504 79970 117556 79976
rect 117516 71777 117544 79970
rect 117318 71768 117374 71777
rect 117318 71703 117374 71712
rect 117502 71768 117558 71777
rect 117502 71703 117558 71712
rect 117332 62150 117360 71703
rect 117320 62144 117372 62150
rect 117320 62086 117372 62092
rect 117596 62144 117648 62150
rect 117596 62086 117648 62092
rect 117608 60858 117636 62086
rect 117596 60852 117648 60858
rect 117596 60794 117648 60800
rect 117504 60716 117556 60722
rect 117504 60658 117556 60664
rect 117516 52465 117544 60658
rect 117502 52456 117558 52465
rect 117502 52391 117558 52400
rect 117686 52456 117742 52465
rect 117686 52391 117742 52400
rect 117700 39370 117728 52391
rect 117688 39364 117740 39370
rect 117688 39306 117740 39312
rect 117596 27668 117648 27674
rect 117596 27610 117648 27616
rect 117608 24834 117636 27610
rect 117516 24806 117636 24834
rect 117516 22166 117544 24806
rect 117504 22160 117556 22166
rect 117504 22102 117556 22108
rect 117412 15224 117464 15230
rect 117412 15166 117464 15172
rect 115848 10532 115900 10538
rect 115848 10474 115900 10480
rect 117136 8220 117188 8226
rect 117136 8162 117188 8168
rect 114468 5092 114520 5098
rect 114468 5034 114520 5040
rect 115754 3768 115810 3777
rect 115754 3703 115756 3712
rect 115808 3703 115810 3712
rect 115938 3768 115994 3777
rect 115938 3703 115994 3712
rect 116858 3768 116914 3777
rect 116858 3703 116860 3712
rect 115756 3674 115808 3680
rect 114742 2952 114798 2961
rect 114742 2887 114798 2896
rect 114756 480 114784 2887
rect 115952 480 115980 3703
rect 116912 3703 116914 3712
rect 116860 3674 116912 3680
rect 117148 480 117176 8162
rect 117424 6866 117452 15166
rect 117412 6860 117464 6866
rect 117412 6802 117464 6808
rect 118240 6860 118292 6866
rect 118240 6802 118292 6808
rect 118252 480 118280 6802
rect 118620 5030 118648 122046
rect 120552 115818 120580 122674
rect 124218 122632 124274 122641
rect 124218 122567 124274 122576
rect 124232 122482 124260 122567
rect 124324 122482 124352 122674
rect 128360 122664 128412 122670
rect 133800 122641 133828 122674
rect 143632 122664 143684 122670
rect 128360 122606 128412 122612
rect 133786 122632 133842 122641
rect 124232 122454 124352 122482
rect 124232 122318 124352 122346
rect 124232 122233 124260 122318
rect 124218 122224 124274 122233
rect 124218 122159 124274 122168
rect 120644 118862 120672 122060
rect 123036 121786 123064 122060
rect 124324 122058 124352 122318
rect 124312 122052 124364 122058
rect 124312 121994 124364 122000
rect 123024 121780 123076 121786
rect 123024 121722 123076 121728
rect 125428 118930 125456 122060
rect 127820 121038 127848 122060
rect 127808 121032 127860 121038
rect 127808 120974 127860 120980
rect 125416 118924 125468 118930
rect 125416 118866 125468 118872
rect 120632 118856 120684 118862
rect 120632 118798 120684 118804
rect 120460 115790 120580 115818
rect 121366 115832 121422 115841
rect 120460 106298 120488 115790
rect 121366 115767 121422 115776
rect 121380 108934 121408 115767
rect 121368 108928 121420 108934
rect 121368 108870 121420 108876
rect 121552 108928 121604 108934
rect 121552 108870 121604 108876
rect 120368 106270 120488 106298
rect 121564 106298 121592 108870
rect 121564 106270 121684 106298
rect 120368 95334 120396 106270
rect 121472 99414 121500 99445
rect 121656 99414 121684 106270
rect 121460 99408 121512 99414
rect 121644 99408 121696 99414
rect 121512 99356 121644 99362
rect 121460 99350 121696 99356
rect 121472 99334 121684 99350
rect 120264 95328 120316 95334
rect 120264 95270 120316 95276
rect 120356 95328 120408 95334
rect 120356 95270 120408 95276
rect 120276 92478 120304 95270
rect 120264 92472 120316 92478
rect 120264 92414 120316 92420
rect 120356 92472 120408 92478
rect 120356 92414 120408 92420
rect 120368 82890 120396 92414
rect 121656 89758 121684 99334
rect 121460 89752 121512 89758
rect 121460 89694 121512 89700
rect 121644 89752 121696 89758
rect 121644 89694 121696 89700
rect 120356 82884 120408 82890
rect 120356 82826 120408 82832
rect 120356 81456 120408 81462
rect 120356 81398 120408 81404
rect 120368 80170 120396 81398
rect 120356 80164 120408 80170
rect 120356 80106 120408 80112
rect 121472 80050 121500 89694
rect 120264 80028 120316 80034
rect 121472 80022 121684 80050
rect 120264 79970 120316 79976
rect 120276 71777 120304 79970
rect 120078 71768 120134 71777
rect 120078 71703 120134 71712
rect 120262 71768 120318 71777
rect 120262 71703 120318 71712
rect 120092 62150 120120 71703
rect 120080 62144 120132 62150
rect 120080 62086 120132 62092
rect 120356 62144 120408 62150
rect 120356 62086 120408 62092
rect 120368 60858 120396 62086
rect 120356 60852 120408 60858
rect 120356 60794 120408 60800
rect 120264 60716 120316 60722
rect 120264 60658 120316 60664
rect 120276 52465 120304 60658
rect 120262 52456 120318 52465
rect 120262 52391 120318 52400
rect 120446 52456 120502 52465
rect 120446 52391 120502 52400
rect 120460 39370 120488 52391
rect 121656 45626 121684 80022
rect 121552 45620 121604 45626
rect 121552 45562 121604 45568
rect 121644 45620 121696 45626
rect 121644 45562 121696 45568
rect 121564 41426 121592 45562
rect 121564 41398 121684 41426
rect 120448 39364 120500 39370
rect 120448 39306 120500 39312
rect 121656 31634 121684 41398
rect 121564 31606 121684 31634
rect 120356 27668 120408 27674
rect 120356 27610 120408 27616
rect 120368 24857 120396 27610
rect 120078 24848 120134 24857
rect 120078 24783 120134 24792
rect 120354 24848 120410 24857
rect 120354 24783 120410 24792
rect 119528 17468 119580 17474
rect 119528 17410 119580 17416
rect 119540 12510 119568 17410
rect 120092 15230 120120 24783
rect 121564 22114 121592 31606
rect 121564 22086 121684 22114
rect 120080 15224 120132 15230
rect 120080 15166 120132 15172
rect 120172 15224 120224 15230
rect 120172 15166 120224 15172
rect 119528 12504 119580 12510
rect 119528 12446 119580 12452
rect 119436 12436 119488 12442
rect 119436 12378 119488 12384
rect 118608 5024 118660 5030
rect 118608 4966 118660 4972
rect 118700 2984 118752 2990
rect 118700 2926 118752 2932
rect 118712 2825 118740 2926
rect 118698 2816 118754 2825
rect 118698 2751 118754 2760
rect 119448 480 119476 12378
rect 120184 6934 120212 15166
rect 121656 12458 121684 22086
rect 121472 12430 121684 12458
rect 128372 12442 128400 122606
rect 133786 122567 133842 122576
rect 143538 122632 143594 122641
rect 153108 122664 153160 122670
rect 143632 122606 143684 122612
rect 149058 122632 149114 122641
rect 143538 122567 143594 122576
rect 143552 122482 143580 122567
rect 143644 122482 143672 122606
rect 149058 122567 149114 122576
rect 153106 122632 153108 122641
rect 249892 122664 249944 122670
rect 153160 122632 153162 122641
rect 153106 122567 153162 122576
rect 201314 122632 201370 122641
rect 201314 122567 201370 122576
rect 216586 122632 216642 122641
rect 249892 122606 249944 122612
rect 259368 122664 259420 122670
rect 259368 122606 259420 122612
rect 284208 122664 284260 122670
rect 284208 122606 284260 122612
rect 216586 122567 216642 122576
rect 143552 122454 143672 122482
rect 143552 122318 143672 122346
rect 143552 122233 143580 122318
rect 133786 122224 133842 122233
rect 133786 122159 133842 122168
rect 143538 122224 143594 122233
rect 143538 122159 143594 122168
rect 131210 122088 131266 122097
rect 129740 121848 129792 121854
rect 129740 121790 129792 121796
rect 128360 12436 128412 12442
rect 120276 6934 120304 6965
rect 120172 6928 120224 6934
rect 120172 6870 120224 6876
rect 120264 6928 120316 6934
rect 120316 6876 120396 6882
rect 120264 6870 120396 6876
rect 120276 6854 120396 6870
rect 120368 3346 120396 6854
rect 120368 3318 120672 3346
rect 120644 480 120672 3318
rect 121472 3074 121500 12430
rect 128360 12378 128412 12384
rect 129004 12436 129056 12442
rect 129004 12378 129056 12384
rect 126612 9308 126664 9314
rect 126612 9250 126664 9256
rect 124220 7812 124272 7818
rect 124220 7754 124272 7760
rect 122010 3496 122066 3505
rect 122010 3431 122066 3440
rect 123022 3496 123078 3505
rect 123022 3431 123078 3440
rect 121472 3046 121684 3074
rect 121656 2666 121684 3046
rect 122024 2961 122052 3431
rect 122932 3052 122984 3058
rect 122932 2994 122984 3000
rect 122010 2952 122066 2961
rect 122010 2887 122066 2896
rect 122944 2825 122972 2994
rect 122930 2816 122986 2825
rect 122930 2751 122986 2760
rect 121656 2638 121868 2666
rect 121840 480 121868 2638
rect 123036 480 123064 3431
rect 124232 480 124260 7754
rect 125414 2952 125470 2961
rect 125414 2887 125470 2896
rect 125428 480 125456 2887
rect 126624 480 126652 9250
rect 127808 5228 127860 5234
rect 127808 5170 127860 5176
rect 127820 480 127848 5170
rect 129016 480 129044 12378
rect 129752 3126 129780 121790
rect 130028 119649 130056 122060
rect 131210 122023 131266 122032
rect 130014 119640 130070 119649
rect 130014 119575 130070 119584
rect 131224 115938 131252 122023
rect 132420 118794 132448 122060
rect 133800 122058 133828 122159
rect 140686 122088 140742 122097
rect 133788 122052 133840 122058
rect 134826 122046 135208 122074
rect 133788 121994 133840 122000
rect 132408 118788 132460 118794
rect 132408 118730 132460 118736
rect 132592 118108 132644 118114
rect 132592 118050 132644 118056
rect 131212 115932 131264 115938
rect 131212 115874 131264 115880
rect 131212 106344 131264 106350
rect 131212 106286 131264 106292
rect 131224 96626 131252 106286
rect 131212 96620 131264 96626
rect 131212 96562 131264 96568
rect 131212 87032 131264 87038
rect 131212 86974 131264 86980
rect 131224 19310 131252 86974
rect 131212 19304 131264 19310
rect 131212 19246 131264 19252
rect 131212 9716 131264 9722
rect 131212 9658 131264 9664
rect 129740 3120 129792 3126
rect 129740 3062 129792 3068
rect 130200 3120 130252 3126
rect 130200 3062 130252 3068
rect 130212 480 130240 3062
rect 131224 2836 131252 9658
rect 131224 2808 131344 2836
rect 131316 2666 131344 2808
rect 131316 2638 131436 2666
rect 131408 480 131436 2638
rect 132604 480 132632 118050
rect 135076 86284 135128 86290
rect 135076 86226 135128 86232
rect 135088 12510 135116 86226
rect 135076 12504 135128 12510
rect 135076 12446 135128 12452
rect 134892 12436 134944 12442
rect 134892 12378 134944 12384
rect 134904 9654 134932 12378
rect 135180 10334 135208 122046
rect 137204 120086 137232 122060
rect 137192 120080 137244 120086
rect 137192 120022 137244 120028
rect 139596 119785 139624 122060
rect 140686 122023 140742 122032
rect 139582 119776 139638 119785
rect 139582 119711 139638 119720
rect 136548 116680 136600 116686
rect 136548 116622 136600 116628
rect 135168 10328 135220 10334
rect 135168 10270 135220 10276
rect 134892 9648 134944 9654
rect 134892 9590 134944 9596
rect 136560 3126 136588 116622
rect 138480 12096 138532 12102
rect 138480 12038 138532 12044
rect 137284 10532 137336 10538
rect 137284 10474 137336 10480
rect 136088 3120 136140 3126
rect 136088 3062 136140 3068
rect 136548 3120 136600 3126
rect 136548 3062 136600 3068
rect 133788 2848 133840 2854
rect 133788 2790 133840 2796
rect 133800 480 133828 2790
rect 134892 604 134944 610
rect 134892 546 134944 552
rect 134904 480 134932 546
rect 136100 480 136128 3062
rect 137296 480 137324 10474
rect 138492 480 138520 12038
rect 140700 3126 140728 122023
rect 141988 119513 142016 122060
rect 143644 122058 143672 122318
rect 143632 122052 143684 122058
rect 143632 121994 143684 122000
rect 142158 121680 142214 121689
rect 142158 121615 142214 121624
rect 141974 119504 142030 119513
rect 141974 119439 142030 119448
rect 140872 4956 140924 4962
rect 140872 4898 140924 4904
rect 139676 3120 139728 3126
rect 139676 3062 139728 3068
rect 140688 3120 140740 3126
rect 140688 3062 140740 3068
rect 139688 480 139716 3062
rect 140884 480 140912 4898
rect 142172 3126 142200 121615
rect 144380 121038 144408 122060
rect 146390 121816 146446 121825
rect 146390 121751 146446 121760
rect 144368 121032 144420 121038
rect 144368 120974 144420 120980
rect 146206 119640 146262 119649
rect 146206 119575 146262 119584
rect 144460 4956 144512 4962
rect 144460 4898 144512 4904
rect 143446 3632 143502 3641
rect 143446 3567 143502 3576
rect 142160 3120 142212 3126
rect 142160 3062 142212 3068
rect 143264 3120 143316 3126
rect 143264 3062 143316 3068
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 142080 480 142108 2790
rect 143276 480 143304 3062
rect 143460 2961 143488 3567
rect 143446 2952 143502 2961
rect 143446 2887 143502 2896
rect 144472 480 144500 4898
rect 146220 3126 146248 119575
rect 146404 3126 146432 121751
rect 146772 120970 146800 122060
rect 149072 121961 149100 122567
rect 179418 122496 179474 122505
rect 167000 122460 167052 122466
rect 167000 122402 167052 122408
rect 172612 122460 172664 122466
rect 201328 122482 201356 122567
rect 209686 122496 209742 122505
rect 179418 122431 179474 122440
rect 182088 122460 182140 122466
rect 172612 122402 172664 122408
rect 162872 122318 162992 122346
rect 162872 122233 162900 122318
rect 153106 122224 153162 122233
rect 153106 122159 153162 122168
rect 162858 122224 162914 122233
rect 162858 122159 162914 122168
rect 149058 121952 149114 121961
rect 149058 121887 149114 121896
rect 149058 121816 149114 121825
rect 149058 121751 149114 121760
rect 146760 120964 146812 120970
rect 146760 120906 146812 120912
rect 148046 3496 148102 3505
rect 148046 3431 148102 3440
rect 145656 3120 145708 3126
rect 145656 3062 145708 3068
rect 146208 3120 146260 3126
rect 146208 3062 146260 3068
rect 146392 3120 146444 3126
rect 146392 3062 146444 3068
rect 146852 3120 146904 3126
rect 146852 3062 146904 3068
rect 145668 480 145696 3062
rect 146864 480 146892 3062
rect 148060 480 148088 3431
rect 149072 1442 149100 121751
rect 149164 120086 149192 122060
rect 150624 120692 150676 120698
rect 150624 120634 150676 120640
rect 149152 120080 149204 120086
rect 149152 120022 149204 120028
rect 150348 120080 150400 120086
rect 150348 120022 150400 120028
rect 150360 9110 150388 120022
rect 150348 9104 150400 9110
rect 150348 9046 150400 9052
rect 150636 1442 150664 120634
rect 151556 119338 151584 122060
rect 153120 122058 153148 122159
rect 153108 122052 153160 122058
rect 153962 122046 154528 122074
rect 153108 121994 153160 122000
rect 153198 121952 153254 121961
rect 153198 121887 153254 121896
rect 153106 119776 153162 119785
rect 153106 119711 153162 119720
rect 151544 119332 151596 119338
rect 151544 119274 151596 119280
rect 153120 116006 153148 119711
rect 153016 116000 153068 116006
rect 153016 115942 153068 115948
rect 153108 116000 153160 116006
rect 153108 115942 153160 115948
rect 153028 115870 153056 115942
rect 153016 115864 153068 115870
rect 153016 115806 153068 115812
rect 153016 108928 153068 108934
rect 153016 108870 153068 108876
rect 153028 106298 153056 108870
rect 153028 106270 153148 106298
rect 153120 95266 153148 106270
rect 152924 95260 152976 95266
rect 152924 95202 152976 95208
rect 153108 95260 153160 95266
rect 153108 95202 153160 95208
rect 152936 70417 152964 95202
rect 152922 70408 152978 70417
rect 152922 70343 152978 70352
rect 152830 67688 152886 67697
rect 152830 67623 152886 67632
rect 152844 66230 152872 67623
rect 152832 66224 152884 66230
rect 152832 66166 152884 66172
rect 152924 66224 152976 66230
rect 152924 66166 152976 66172
rect 152936 61441 152964 66166
rect 152922 61432 152978 61441
rect 152922 61367 152978 61376
rect 153014 50960 153070 50969
rect 153014 50895 153070 50904
rect 153028 41426 153056 50895
rect 153028 41398 153148 41426
rect 153120 31822 153148 41398
rect 153108 31816 153160 31822
rect 153108 31758 153160 31764
rect 152924 29028 152976 29034
rect 152924 28970 152976 28976
rect 152936 27606 152964 28970
rect 152924 27600 152976 27606
rect 152924 27542 152976 27548
rect 153016 18012 153068 18018
rect 153016 17954 153068 17960
rect 153028 12510 153056 17954
rect 153016 12504 153068 12510
rect 153016 12446 153068 12452
rect 152740 12436 152792 12442
rect 152740 12378 152792 12384
rect 151726 10296 151782 10305
rect 151726 10231 151782 10240
rect 151740 1442 151768 10231
rect 149072 1414 149284 1442
rect 149256 480 149284 1414
rect 150452 1414 150664 1442
rect 151556 1414 151768 1442
rect 150452 480 150480 1414
rect 151556 480 151584 1414
rect 152752 480 152780 12378
rect 153106 3632 153162 3641
rect 153106 3567 153162 3576
rect 153120 2961 153148 3567
rect 153212 3126 153240 121887
rect 154500 12034 154528 122046
rect 156340 119950 156368 122060
rect 158732 121417 158760 122060
rect 158718 121408 158774 121417
rect 158718 121343 158774 121352
rect 156328 119944 156380 119950
rect 156328 119886 156380 119892
rect 161124 119066 161152 122060
rect 162964 122058 162992 122318
rect 162952 122052 163004 122058
rect 162952 121994 163004 122000
rect 163516 120834 163544 122060
rect 165908 120970 165936 122060
rect 165896 120964 165948 120970
rect 165896 120906 165948 120912
rect 163504 120828 163556 120834
rect 163504 120770 163556 120776
rect 161112 119060 161164 119066
rect 161112 119002 161164 119008
rect 156052 118652 156104 118658
rect 156052 118594 156104 118600
rect 156064 115954 156092 118594
rect 161480 116816 161532 116822
rect 161480 116758 161532 116764
rect 161296 116068 161348 116074
rect 161296 116010 161348 116016
rect 156064 115938 156184 115954
rect 161308 115938 161336 116010
rect 155868 115932 155920 115938
rect 156064 115932 156196 115938
rect 156064 115926 156144 115932
rect 155868 115874 155920 115880
rect 156144 115874 156196 115880
rect 161296 115932 161348 115938
rect 161296 115874 161348 115880
rect 155880 114510 155908 115874
rect 156156 115843 156184 115874
rect 155868 114504 155920 114510
rect 155868 114446 155920 114452
rect 161296 108928 161348 108934
rect 161296 108870 161348 108876
rect 161308 106298 161336 108870
rect 161308 106270 161428 106298
rect 156052 104916 156104 104922
rect 156052 104858 156104 104864
rect 156064 104802 156092 104858
rect 156064 104786 156184 104802
rect 156064 104780 156196 104786
rect 156064 104774 156144 104780
rect 156144 104722 156196 104728
rect 161400 99414 161428 106270
rect 161204 99408 161256 99414
rect 161204 99350 161256 99356
rect 161388 99408 161440 99414
rect 161388 99350 161440 99356
rect 161216 96626 161244 99350
rect 161204 96620 161256 96626
rect 161204 96562 161256 96568
rect 161296 96620 161348 96626
rect 161296 96562 161348 96568
rect 156236 95260 156288 95266
rect 156236 95202 156288 95208
rect 156248 89434 156276 95202
rect 156156 89406 156276 89434
rect 156156 76022 156184 89406
rect 161308 85610 161336 96562
rect 161020 85604 161072 85610
rect 161020 85546 161072 85552
rect 161296 85604 161348 85610
rect 161296 85546 161348 85552
rect 155960 76016 156012 76022
rect 155960 75958 156012 75964
rect 156144 76016 156196 76022
rect 156144 75958 156196 75964
rect 155972 70446 156000 75958
rect 161032 75954 161060 85546
rect 161020 75948 161072 75954
rect 161020 75890 161072 75896
rect 161204 75948 161256 75954
rect 161204 75890 161256 75896
rect 155960 70440 156012 70446
rect 155960 70382 156012 70388
rect 156144 70304 156196 70310
rect 156144 70246 156196 70252
rect 156156 66230 156184 70246
rect 161216 66314 161244 75890
rect 161032 66286 161244 66314
rect 156144 66224 156196 66230
rect 156144 66166 156196 66172
rect 161032 64870 161060 66286
rect 161020 64864 161072 64870
rect 161020 64806 161072 64812
rect 155960 56636 156012 56642
rect 155960 56578 156012 56584
rect 155972 50930 156000 56578
rect 161388 55276 161440 55282
rect 161388 55218 161440 55224
rect 155960 50924 156012 50930
rect 155960 50866 156012 50872
rect 156144 50924 156196 50930
rect 156144 50866 156196 50872
rect 156156 46918 156184 50866
rect 161400 48346 161428 55218
rect 161112 48340 161164 48346
rect 161112 48282 161164 48288
rect 161388 48340 161440 48346
rect 161388 48282 161440 48288
rect 161124 46918 161152 48282
rect 156144 46912 156196 46918
rect 156144 46854 156196 46860
rect 161112 46912 161164 46918
rect 161112 46854 161164 46860
rect 156052 41404 156104 41410
rect 156052 41346 156104 41352
rect 156064 31754 156092 41346
rect 161204 37324 161256 37330
rect 161204 37266 161256 37272
rect 161216 32502 161244 37266
rect 161204 32496 161256 32502
rect 161204 32438 161256 32444
rect 156052 31748 156104 31754
rect 156052 31690 156104 31696
rect 156236 31748 156288 31754
rect 156236 31690 156288 31696
rect 156248 28966 156276 31690
rect 161492 28966 161520 116758
rect 156236 28960 156288 28966
rect 156236 28902 156288 28908
rect 161480 28960 161532 28966
rect 161480 28902 161532 28908
rect 161204 27668 161256 27674
rect 161204 27610 161256 27616
rect 161216 27554 161244 27610
rect 161216 27526 161336 27554
rect 161308 20602 161336 27526
rect 161112 20596 161164 20602
rect 161112 20538 161164 20544
rect 161296 20596 161348 20602
rect 161296 20538 161348 20544
rect 156144 19372 156196 19378
rect 156144 19314 156196 19320
rect 156156 14618 156184 19314
rect 158628 15904 158680 15910
rect 158628 15846 158680 15852
rect 156144 14612 156196 14618
rect 156144 14554 156196 14560
rect 154488 12028 154540 12034
rect 154488 11970 154540 11976
rect 155132 11892 155184 11898
rect 155132 11834 155184 11840
rect 153200 3120 153252 3126
rect 153200 3062 153252 3068
rect 153936 3120 153988 3126
rect 153936 3062 153988 3068
rect 153106 2952 153162 2961
rect 153106 2887 153162 2896
rect 153948 480 153976 3062
rect 155144 480 155172 11834
rect 156236 9716 156288 9722
rect 156236 9658 156288 9664
rect 156248 2802 156276 9658
rect 158640 3058 158668 15846
rect 159916 6656 159968 6662
rect 159916 6598 159968 6604
rect 157524 3052 157576 3058
rect 157524 2994 157576 3000
rect 158628 3052 158680 3058
rect 158628 2994 158680 3000
rect 156156 2774 156276 2802
rect 156156 2666 156184 2774
rect 156156 2638 156368 2666
rect 156340 480 156368 2638
rect 157536 480 157564 2994
rect 158720 2916 158772 2922
rect 158720 2858 158772 2864
rect 158732 480 158760 2858
rect 159928 480 159956 6598
rect 161124 480 161152 20538
rect 161572 18012 161624 18018
rect 161572 17954 161624 17960
rect 161584 9722 161612 17954
rect 165526 17368 165582 17377
rect 165526 17303 165582 17312
rect 161480 9716 161532 9722
rect 161480 9658 161532 9664
rect 161572 9716 161624 9722
rect 161572 9658 161624 9664
rect 161492 2938 161520 9658
rect 162952 4208 163004 4214
rect 162952 4150 163004 4156
rect 164700 4208 164752 4214
rect 164700 4150 164752 4156
rect 162122 3768 162178 3777
rect 162122 3703 162178 3712
rect 162136 3505 162164 3703
rect 162766 3632 162822 3641
rect 162964 3618 162992 4150
rect 164712 3777 164740 4150
rect 163502 3768 163558 3777
rect 163502 3703 163558 3712
rect 164698 3768 164754 3777
rect 164698 3703 164754 3712
rect 162766 3567 162822 3576
rect 162872 3590 162992 3618
rect 162122 3496 162178 3505
rect 162122 3431 162178 3440
rect 162780 2961 162808 3567
rect 162872 3505 162900 3590
rect 162858 3496 162914 3505
rect 162858 3431 162914 3440
rect 162858 3360 162914 3369
rect 162858 3295 162914 3304
rect 163318 3360 163374 3369
rect 163318 3295 163374 3304
rect 162872 3210 162900 3295
rect 163332 3210 163360 3295
rect 162872 3182 163360 3210
rect 161400 2910 161520 2938
rect 162766 2952 162822 2961
rect 161400 2786 161428 2910
rect 162766 2887 162822 2896
rect 161388 2780 161440 2786
rect 161388 2722 161440 2728
rect 162308 2780 162360 2786
rect 162308 2722 162360 2728
rect 162320 480 162348 2722
rect 163516 480 163544 3703
rect 165540 3058 165568 17303
rect 167012 3482 167040 122402
rect 167090 122360 167146 122369
rect 167090 122295 167146 122304
rect 169666 122360 169722 122369
rect 169666 122295 169722 122304
rect 167104 3618 167132 122295
rect 168300 121553 168328 122060
rect 168286 121544 168342 121553
rect 168286 121479 168342 121488
rect 167104 3590 167224 3618
rect 167012 3454 167132 3482
rect 164700 3052 164752 3058
rect 164700 2994 164752 3000
rect 165528 3052 165580 3058
rect 165528 2994 165580 3000
rect 164712 480 164740 2994
rect 165896 2984 165948 2990
rect 165896 2926 165948 2932
rect 165908 480 165936 2926
rect 167104 480 167132 3454
rect 167196 3058 167224 3590
rect 169680 3482 169708 122295
rect 172624 122233 172652 122402
rect 172426 122224 172482 122233
rect 172426 122159 172482 122168
rect 172610 122224 172666 122233
rect 172610 122159 172666 122168
rect 170706 122046 171088 122074
rect 172440 122058 172468 122159
rect 172518 122088 172574 122097
rect 169760 118856 169812 118862
rect 169760 118798 169812 118804
rect 169772 3618 169800 118798
rect 171060 8090 171088 122046
rect 172428 122052 172480 122058
rect 172518 122023 172520 122032
rect 172428 121994 172480 122000
rect 172572 122023 172574 122032
rect 172794 122088 172850 122097
rect 172794 122023 172796 122032
rect 172520 121994 172572 122000
rect 172848 122023 172850 122032
rect 172796 121994 172848 122000
rect 173084 121174 173112 122060
rect 173898 121816 173954 121825
rect 173898 121751 173954 121760
rect 173072 121168 173124 121174
rect 173072 121110 173124 121116
rect 173808 10532 173860 10538
rect 173808 10474 173860 10480
rect 171784 9444 171836 9450
rect 171784 9386 171836 9392
rect 171048 8084 171100 8090
rect 171048 8026 171100 8032
rect 169772 3590 170628 3618
rect 169404 3454 169708 3482
rect 167184 3052 167236 3058
rect 167184 2994 167236 3000
rect 168196 3052 168248 3058
rect 168196 2994 168248 3000
rect 168208 480 168236 2994
rect 169404 480 169432 3454
rect 170600 480 170628 3590
rect 171796 480 171824 9386
rect 173820 3058 173848 10474
rect 173912 3482 173940 121751
rect 175292 121650 175320 122060
rect 175280 121644 175332 121650
rect 175280 121586 175332 121592
rect 179328 119944 179380 119950
rect 179328 119886 179380 119892
rect 176658 118824 176714 118833
rect 176658 118759 176714 118768
rect 176568 5296 176620 5302
rect 176568 5238 176620 5244
rect 175370 3496 175426 3505
rect 173912 3454 174216 3482
rect 172980 3052 173032 3058
rect 172980 2994 173032 3000
rect 173808 3052 173860 3058
rect 173808 2994 173860 3000
rect 172992 480 173020 2994
rect 174188 480 174216 3454
rect 175370 3431 175426 3440
rect 175384 480 175412 3431
rect 176580 480 176608 5238
rect 176672 3058 176700 118759
rect 179340 115938 179368 119886
rect 179328 115932 179380 115938
rect 179328 115874 179380 115880
rect 179328 106412 179380 106418
rect 179328 106354 179380 106360
rect 179340 104854 179368 106354
rect 179328 104848 179380 104854
rect 179328 104790 179380 104796
rect 179328 87100 179380 87106
rect 179328 87042 179380 87048
rect 179340 85542 179368 87042
rect 179328 85536 179380 85542
rect 179328 85478 179380 85484
rect 179328 75948 179380 75954
rect 179328 75890 179380 75896
rect 179340 67833 179368 75890
rect 179326 67824 179382 67833
rect 179326 67759 179382 67768
rect 179326 67688 179382 67697
rect 179326 67623 179382 67632
rect 179340 66230 179368 67623
rect 179328 66224 179380 66230
rect 179328 66166 179380 66172
rect 179328 56636 179380 56642
rect 179328 56578 179380 56584
rect 179340 48498 179368 56578
rect 179248 48470 179368 48498
rect 179248 48362 179276 48470
rect 179248 48334 179368 48362
rect 179340 46918 179368 48334
rect 179328 46912 179380 46918
rect 179328 46854 179380 46860
rect 179236 37324 179288 37330
rect 179236 37266 179288 37272
rect 179248 29050 179276 37266
rect 179248 29022 179368 29050
rect 179340 27606 179368 29022
rect 179328 27600 179380 27606
rect 179328 27542 179380 27548
rect 178960 9716 179012 9722
rect 178960 9658 179012 9664
rect 176660 3052 176712 3058
rect 176660 2994 176712 3000
rect 177764 3052 177816 3058
rect 177764 2994 177816 3000
rect 177776 480 177804 2994
rect 178972 480 179000 9658
rect 179432 3126 179460 122431
rect 201328 122454 201448 122482
rect 182088 122402 182140 122408
rect 182100 122233 182128 122402
rect 201420 122369 201448 122454
rect 209686 122431 209742 122440
rect 201406 122360 201462 122369
rect 201406 122295 201462 122304
rect 205640 122256 205692 122262
rect 182086 122224 182142 122233
rect 182086 122159 182142 122168
rect 182362 122224 182418 122233
rect 182362 122159 182418 122168
rect 191746 122224 191802 122233
rect 205640 122198 205692 122204
rect 191746 122159 191802 122168
rect 196072 122188 196124 122194
rect 180076 119066 180104 122060
rect 182376 122058 182404 122159
rect 182364 122052 182416 122058
rect 182364 121994 182416 122000
rect 182468 121281 182496 122060
rect 183572 122046 184874 122074
rect 182454 121272 182510 121281
rect 182454 121207 182510 121216
rect 180064 119060 180116 119066
rect 180064 119002 180116 119008
rect 183468 115320 183520 115326
rect 183468 115262 183520 115268
rect 181352 12164 181404 12170
rect 181352 12106 181404 12112
rect 179420 3120 179472 3126
rect 179420 3062 179472 3068
rect 180156 3120 180208 3126
rect 180156 3062 180208 3068
rect 180168 480 180196 3062
rect 181364 480 181392 12106
rect 182086 3632 182142 3641
rect 182086 3567 182142 3576
rect 182100 2961 182128 3567
rect 183480 3126 183508 115262
rect 183572 5302 183600 122046
rect 187252 121281 187280 122060
rect 187238 121272 187294 121281
rect 187238 121207 187294 121216
rect 189644 121174 189672 122060
rect 191760 122058 191788 122159
rect 196072 122130 196124 122136
rect 198648 122188 198700 122194
rect 198648 122130 198700 122136
rect 191748 122052 191800 122058
rect 191748 121994 191800 122000
rect 191852 122046 192050 122074
rect 189632 121168 189684 121174
rect 189632 121110 189684 121116
rect 190458 119232 190514 119241
rect 190458 119167 190514 119176
rect 187698 118960 187754 118969
rect 187698 118895 187754 118904
rect 186228 114572 186280 114578
rect 186228 114514 186280 114520
rect 186240 104854 186268 114514
rect 186228 104848 186280 104854
rect 186228 104790 186280 104796
rect 186228 95260 186280 95266
rect 186228 95202 186280 95208
rect 186240 85542 186268 95202
rect 186228 85536 186280 85542
rect 186228 85478 186280 85484
rect 186228 75948 186280 75954
rect 186228 75890 186280 75896
rect 186240 66230 186268 75890
rect 186228 66224 186280 66230
rect 186228 66166 186280 66172
rect 186228 56636 186280 56642
rect 186228 56578 186280 56584
rect 186240 46918 186268 56578
rect 186228 46912 186280 46918
rect 186228 46854 186280 46860
rect 186228 37324 186280 37330
rect 186228 37266 186280 37272
rect 186240 27606 186268 37266
rect 186228 27600 186280 27606
rect 186228 27542 186280 27548
rect 184848 13320 184900 13326
rect 184848 13262 184900 13268
rect 183744 7540 183796 7546
rect 183744 7482 183796 7488
rect 183560 5296 183612 5302
rect 183560 5238 183612 5244
rect 182548 3120 182600 3126
rect 182548 3062 182600 3068
rect 183468 3120 183520 3126
rect 183468 3062 183520 3068
rect 182086 2952 182142 2961
rect 182086 2887 182142 2896
rect 182560 480 182588 3062
rect 183756 480 183784 7482
rect 184860 480 184888 13262
rect 186044 9784 186096 9790
rect 186044 9726 186096 9732
rect 186056 9654 186084 9726
rect 186044 9648 186096 9654
rect 186044 9590 186096 9596
rect 187240 5092 187292 5098
rect 187240 5034 187292 5040
rect 186044 604 186096 610
rect 186044 546 186096 552
rect 186056 480 186084 546
rect 187252 480 187280 5034
rect 187712 3126 187740 118895
rect 190366 17504 190422 17513
rect 190366 17439 190422 17448
rect 190380 3126 190408 17439
rect 187700 3120 187752 3126
rect 187700 3062 187752 3068
rect 188436 3120 188488 3126
rect 188436 3062 188488 3068
rect 189632 3120 189684 3126
rect 189632 3062 189684 3068
rect 190368 3120 190420 3126
rect 190368 3062 190420 3068
rect 188448 480 188476 3062
rect 189644 480 189672 3062
rect 190472 2938 190500 119167
rect 191852 10538 191880 122046
rect 194428 119542 194456 122060
rect 194416 119536 194468 119542
rect 194416 119478 194468 119484
rect 193218 119096 193274 119105
rect 193218 119031 193274 119040
rect 193128 13524 193180 13530
rect 193128 13466 193180 13472
rect 191840 10532 191892 10538
rect 191840 10474 191892 10480
rect 193140 3126 193168 13466
rect 192024 3120 192076 3126
rect 192024 3062 192076 3068
rect 193128 3120 193180 3126
rect 193128 3062 193180 3068
rect 190380 2910 190500 2938
rect 190380 610 190408 2910
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 190828 604 190880 610
rect 190828 546 190880 552
rect 190840 480 190868 546
rect 192036 480 192064 3062
rect 193232 480 193260 119031
rect 195426 14648 195482 14657
rect 195426 14583 195482 14592
rect 194416 10532 194468 10538
rect 194416 10474 194468 10480
rect 194428 480 194456 10474
rect 195440 9761 195468 14583
rect 196084 12442 196112 122130
rect 196622 122088 196678 122097
rect 196622 122023 196678 122032
rect 196636 121825 196664 122023
rect 196622 121816 196678 121825
rect 196622 121751 196678 121760
rect 196820 119134 196848 122060
rect 196808 119128 196860 119134
rect 196808 119070 196860 119076
rect 196072 12436 196124 12442
rect 196072 12378 196124 12384
rect 196808 12436 196860 12442
rect 196808 12378 196860 12384
rect 195426 9752 195482 9761
rect 195426 9687 195482 9696
rect 195610 9752 195666 9761
rect 195610 9687 195666 9696
rect 195624 9654 195652 9687
rect 195612 9648 195664 9654
rect 195612 9590 195664 9596
rect 195612 9512 195664 9518
rect 195612 9454 195664 9460
rect 195624 480 195652 9454
rect 196820 480 196848 12378
rect 198660 3126 198688 122130
rect 199212 120086 199240 122060
rect 201604 120086 201632 122060
rect 199200 120080 199252 120086
rect 199200 120022 199252 120028
rect 200028 120080 200080 120086
rect 200028 120022 200080 120028
rect 201592 120080 201644 120086
rect 201592 120022 201644 120028
rect 199934 16280 199990 16289
rect 199934 16215 199990 16224
rect 199948 3126 199976 16215
rect 200040 14618 200068 120022
rect 201498 119912 201554 119921
rect 201498 119847 201554 119856
rect 201408 118788 201460 118794
rect 201408 118730 201460 118736
rect 200028 14612 200080 14618
rect 200028 14554 200080 14560
rect 201420 3126 201448 118730
rect 201512 3126 201540 119847
rect 203996 118998 204024 122060
rect 203984 118992 204036 118998
rect 203984 118934 204036 118940
rect 204166 16416 204222 16425
rect 204166 16351 204222 16360
rect 201592 5296 201644 5302
rect 201592 5238 201644 5244
rect 198004 3120 198056 3126
rect 198004 3062 198056 3068
rect 198648 3120 198700 3126
rect 198648 3062 198700 3068
rect 199200 3120 199252 3126
rect 199200 3062 199252 3068
rect 199936 3120 199988 3126
rect 199936 3062 199988 3068
rect 200396 3120 200448 3126
rect 200396 3062 200448 3068
rect 201408 3120 201460 3126
rect 201408 3062 201460 3068
rect 201500 3120 201552 3126
rect 201500 3062 201552 3068
rect 198016 480 198044 3062
rect 199212 480 199240 3062
rect 200408 480 200436 3062
rect 201604 2666 201632 5238
rect 202696 3120 202748 3126
rect 202696 3062 202748 3068
rect 201512 2638 201632 2666
rect 201512 480 201540 2638
rect 202708 480 202736 3062
rect 204180 626 204208 16351
rect 205088 5024 205140 5030
rect 205088 4966 205140 4972
rect 203904 598 204208 626
rect 203904 480 203932 598
rect 205100 480 205128 4966
rect 205652 610 205680 122198
rect 206388 119134 206416 122060
rect 208780 119202 208808 122060
rect 208768 119196 208820 119202
rect 208768 119138 208820 119144
rect 206376 119128 206428 119134
rect 206376 119070 206428 119076
rect 209700 3874 209728 122431
rect 212540 122392 212592 122398
rect 212262 122360 212318 122369
rect 212446 122360 212502 122369
rect 212318 122318 212446 122346
rect 212262 122295 212318 122304
rect 212540 122334 212592 122340
rect 212446 122295 212502 122304
rect 212448 122256 212500 122262
rect 212448 122198 212500 122204
rect 211172 119542 211200 122060
rect 211160 119536 211212 119542
rect 211160 119478 211212 119484
rect 212356 119536 212408 119542
rect 212356 119478 212408 119484
rect 211068 119196 211120 119202
rect 211068 119138 211120 119144
rect 210976 82136 211028 82142
rect 210976 82078 211028 82084
rect 210988 3874 211016 82078
rect 208676 3868 208728 3874
rect 208676 3810 208728 3816
rect 209688 3868 209740 3874
rect 209688 3810 209740 3816
rect 209872 3868 209924 3874
rect 209872 3810 209924 3816
rect 210976 3868 211028 3874
rect 210976 3810 211028 3816
rect 206926 3768 206982 3777
rect 206926 3703 206982 3712
rect 207478 3768 207534 3777
rect 207478 3703 207534 3712
rect 206940 3505 206968 3703
rect 206926 3496 206982 3505
rect 206926 3431 206982 3440
rect 205640 604 205692 610
rect 205640 546 205692 552
rect 206284 604 206336 610
rect 206284 546 206336 552
rect 206296 480 206324 546
rect 207492 480 207520 3703
rect 208688 480 208716 3810
rect 209884 480 209912 3810
rect 211080 480 211108 119138
rect 212368 5030 212396 119478
rect 212356 5024 212408 5030
rect 212356 4966 212408 4972
rect 212460 4842 212488 122198
rect 212276 4814 212488 4842
rect 212276 480 212304 4814
rect 212552 610 212580 122334
rect 213578 122046 213868 122074
rect 215970 122046 216536 122074
rect 213840 5438 213868 122046
rect 216508 11966 216536 122046
rect 216496 11960 216548 11966
rect 216496 11902 216548 11908
rect 213828 5432 213880 5438
rect 213828 5374 213880 5380
rect 216600 3874 216628 122567
rect 241428 122460 241480 122466
rect 241428 122402 241480 122408
rect 229008 122392 229060 122398
rect 229008 122334 229060 122340
rect 223580 122324 223632 122330
rect 223580 122266 223632 122272
rect 227628 122324 227680 122330
rect 227628 122266 227680 122272
rect 218348 119202 218376 122060
rect 218336 119196 218388 119202
rect 218336 119138 218388 119144
rect 219348 119196 219400 119202
rect 219348 119138 219400 119144
rect 217966 115288 218022 115297
rect 217966 115223 218022 115232
rect 217980 3874 218008 115223
rect 219360 13122 219388 119138
rect 220556 109154 220584 122060
rect 222948 119202 222976 122060
rect 222936 119196 222988 119202
rect 222936 119138 222988 119144
rect 222108 118856 222160 118862
rect 222108 118798 222160 118804
rect 220728 118108 220780 118114
rect 220728 118050 220780 118056
rect 220464 109126 220584 109154
rect 220464 109018 220492 109126
rect 220464 108990 220584 109018
rect 220556 99634 220584 108990
rect 220740 104854 220768 118050
rect 220728 104848 220780 104854
rect 220728 104790 220780 104796
rect 220464 99606 220584 99634
rect 220464 95282 220492 99606
rect 220464 95254 220584 95282
rect 220556 95198 220584 95254
rect 220728 95260 220780 95266
rect 220728 95202 220780 95208
rect 220544 95192 220596 95198
rect 220544 95134 220596 95140
rect 220544 85604 220596 85610
rect 220544 85546 220596 85552
rect 220556 80170 220584 85546
rect 220740 85542 220768 95202
rect 220728 85536 220780 85542
rect 220728 85478 220780 85484
rect 220544 80164 220596 80170
rect 220544 80106 220596 80112
rect 220544 80028 220596 80034
rect 220544 79970 220596 79976
rect 220556 70394 220584 79970
rect 220728 75948 220780 75954
rect 220728 75890 220780 75896
rect 220464 70366 220584 70394
rect 220464 70258 220492 70366
rect 220464 70230 220584 70258
rect 220556 51134 220584 70230
rect 220740 66230 220768 75890
rect 220728 66224 220780 66230
rect 220728 66166 220780 66172
rect 220728 56636 220780 56642
rect 220728 56578 220780 56584
rect 220544 51128 220596 51134
rect 220544 51070 220596 51076
rect 220360 51060 220412 51066
rect 220360 51002 220412 51008
rect 220372 42106 220400 51002
rect 220740 46918 220768 56578
rect 220728 46912 220780 46918
rect 220728 46854 220780 46860
rect 220280 42078 220400 42106
rect 220280 37369 220308 42078
rect 220266 37360 220322 37369
rect 220266 37295 220322 37304
rect 220450 37360 220506 37369
rect 220450 37295 220506 37304
rect 220728 37324 220780 37330
rect 220464 37262 220492 37295
rect 220728 37266 220780 37272
rect 220452 37256 220504 37262
rect 220452 37198 220504 37204
rect 220544 27668 220596 27674
rect 220544 27610 220596 27616
rect 220556 27554 220584 27610
rect 220740 27606 220768 37266
rect 220728 27600 220780 27606
rect 220556 27526 220676 27554
rect 220728 27542 220780 27548
rect 220648 22080 220676 27526
rect 220464 22052 220676 22080
rect 220464 13258 220492 22052
rect 220728 18012 220780 18018
rect 220728 17954 220780 17960
rect 220452 13252 220504 13258
rect 220452 13194 220504 13200
rect 219348 13116 219400 13122
rect 219348 13058 219400 13064
rect 220740 12578 220768 17954
rect 220728 12572 220780 12578
rect 220728 12514 220780 12520
rect 222120 12510 222148 118798
rect 223592 104854 223620 122266
rect 225052 120080 225104 120086
rect 225052 120022 225104 120028
rect 223580 104848 223632 104854
rect 223580 104790 223632 104796
rect 223580 95260 223632 95266
rect 223580 95202 223632 95208
rect 223592 85542 223620 95202
rect 223580 85536 223632 85542
rect 223580 85478 223632 85484
rect 223580 75948 223632 75954
rect 223580 75890 223632 75896
rect 223592 66230 223620 75890
rect 223580 66224 223632 66230
rect 223580 66166 223632 66172
rect 223580 56636 223632 56642
rect 223580 56578 223632 56584
rect 223592 46918 223620 56578
rect 223580 46912 223632 46918
rect 223580 46854 223632 46860
rect 223580 37324 223632 37330
rect 223580 37266 223632 37272
rect 223592 27606 223620 37266
rect 223580 27600 223632 27606
rect 223580 27542 223632 27548
rect 223580 18012 223632 18018
rect 223580 17954 223632 17960
rect 222108 12504 222160 12510
rect 222108 12446 222160 12452
rect 223592 9897 223620 17954
rect 223578 9888 223634 9897
rect 223578 9823 223634 9832
rect 220544 9716 220596 9722
rect 220544 9658 220596 9664
rect 221740 9716 221792 9722
rect 221740 9658 221792 9664
rect 223578 9718 223634 9727
rect 215852 3868 215904 3874
rect 215852 3810 215904 3816
rect 216588 3868 216640 3874
rect 216588 3810 216640 3816
rect 217048 3868 217100 3874
rect 217048 3810 217100 3816
rect 217968 3868 218020 3874
rect 217968 3810 218020 3816
rect 214656 3188 214708 3194
rect 214656 3130 214708 3136
rect 212540 604 212592 610
rect 212540 546 212592 552
rect 213460 604 213512 610
rect 213460 546 213512 552
rect 213472 480 213500 546
rect 214668 480 214696 3130
rect 215864 480 215892 3810
rect 217060 480 217088 3810
rect 219346 3768 219402 3777
rect 219346 3703 219402 3712
rect 220082 3768 220138 3777
rect 220082 3703 220138 3712
rect 218150 2952 218206 2961
rect 218150 2887 218206 2896
rect 218164 480 218192 2887
rect 219360 480 219388 3703
rect 220096 3505 220124 3703
rect 220082 3496 220138 3505
rect 220082 3431 220138 3440
rect 220266 3496 220322 3505
rect 220266 3431 220322 3440
rect 220280 2961 220308 3431
rect 220266 2952 220322 2961
rect 220266 2887 220322 2896
rect 220556 480 220584 9658
rect 221752 480 221780 9658
rect 223578 9653 223634 9662
rect 222936 9376 222988 9382
rect 222936 9318 222988 9324
rect 222948 480 222976 9318
rect 223592 8265 223620 9653
rect 223578 8256 223634 8265
rect 223578 8191 223634 8200
rect 224222 8120 224278 8129
rect 224222 8055 224278 8064
rect 224236 2666 224264 8055
rect 225064 3482 225092 120022
rect 225340 118726 225368 122060
rect 225328 118720 225380 118726
rect 225328 118662 225380 118668
rect 226248 118720 226300 118726
rect 226248 118662 226300 118668
rect 226260 14686 226288 118662
rect 226248 14680 226300 14686
rect 226248 14622 226300 14628
rect 227640 3874 227668 122266
rect 227732 119678 227760 122060
rect 227720 119672 227772 119678
rect 227720 119614 227772 119620
rect 226524 3868 226576 3874
rect 226524 3810 226576 3816
rect 227628 3868 227680 3874
rect 227628 3810 227680 3816
rect 227720 3868 227772 3874
rect 227720 3810 227772 3816
rect 225064 3454 225368 3482
rect 224144 2638 224264 2666
rect 224144 480 224172 2638
rect 225340 480 225368 3454
rect 226536 480 226564 3810
rect 227732 480 227760 3810
rect 229020 3482 229048 122334
rect 239876 122318 240088 122346
rect 230124 119678 230152 122060
rect 230112 119672 230164 119678
rect 230112 119614 230164 119620
rect 232516 119270 232544 122060
rect 234908 119814 234936 122060
rect 237102 121952 237158 121961
rect 237102 121887 237158 121896
rect 234896 119808 234948 119814
rect 234896 119750 234948 119756
rect 232504 119264 232556 119270
rect 232504 119206 232556 119212
rect 233148 118992 233200 118998
rect 233148 118934 233200 118940
rect 230480 12028 230532 12034
rect 230480 11970 230532 11976
rect 230110 5808 230166 5817
rect 230110 5743 230166 5752
rect 228928 3454 229048 3482
rect 228928 480 228956 3454
rect 230124 480 230152 5743
rect 230492 3482 230520 11970
rect 230492 3454 231348 3482
rect 231320 480 231348 3454
rect 233160 3126 233188 118934
rect 233700 5024 233752 5030
rect 233700 4966 233752 4972
rect 232504 3120 232556 3126
rect 232504 3062 232556 3068
rect 233148 3120 233200 3126
rect 233148 3062 233200 3068
rect 232516 480 232544 3062
rect 233712 480 233740 4966
rect 236000 3120 236052 3126
rect 236000 3062 236052 3068
rect 234804 3052 234856 3058
rect 234804 2994 234856 3000
rect 234816 480 234844 2994
rect 236012 480 236040 3062
rect 237116 2938 237144 121887
rect 239692 120834 239720 122060
rect 239876 121689 239904 122318
rect 240060 122233 240088 122318
rect 240046 122224 240102 122233
rect 240046 122159 240102 122168
rect 240322 122224 240378 122233
rect 240322 122159 240378 122168
rect 240336 122058 240364 122159
rect 240324 122052 240376 122058
rect 240324 121994 240376 122000
rect 239862 121680 239918 121689
rect 239862 121615 239918 121624
rect 239680 120828 239732 120834
rect 239680 120770 239732 120776
rect 240048 119264 240100 119270
rect 240048 119206 240100 119212
rect 237196 118856 237248 118862
rect 237196 118798 237248 118804
rect 237208 3126 237236 118798
rect 240060 3126 240088 119206
rect 241440 3126 241468 122402
rect 241518 122224 241574 122233
rect 241518 122159 241574 122168
rect 249798 122224 249854 122233
rect 249798 122159 249854 122168
rect 241532 122058 241560 122159
rect 249812 122074 249840 122159
rect 249904 122074 249932 122606
rect 253848 122596 253900 122602
rect 253848 122538 253900 122544
rect 241520 122052 241572 122058
rect 241520 121994 241572 122000
rect 242084 119814 242112 122060
rect 242806 120728 242862 120737
rect 242806 120663 242862 120672
rect 242072 119808 242124 119814
rect 242072 119750 242124 119756
rect 241518 3632 241574 3641
rect 241518 3567 241574 3576
rect 237196 3120 237248 3126
rect 239588 3120 239640 3126
rect 237196 3062 237248 3068
rect 238390 3088 238446 3097
rect 239588 3062 239640 3068
rect 240048 3120 240100 3126
rect 240048 3062 240100 3068
rect 240784 3120 240836 3126
rect 240784 3062 240836 3068
rect 241428 3120 241480 3126
rect 241428 3062 241480 3068
rect 238390 3023 238446 3032
rect 237116 2910 237236 2938
rect 237208 480 237236 2910
rect 238404 480 238432 3023
rect 239600 480 239628 3062
rect 240796 480 240824 3062
rect 241532 2825 241560 3567
rect 242820 3126 242848 120663
rect 244476 120086 244504 122060
rect 245672 122046 246882 122074
rect 249274 122046 249656 122074
rect 249812 122046 249932 122074
rect 251192 122046 251666 122074
rect 244464 120080 244516 120086
rect 244464 120022 244516 120028
rect 245568 120080 245620 120086
rect 245568 120022 245620 120028
rect 242900 120012 242952 120018
rect 242900 119954 242952 119960
rect 241980 3120 242032 3126
rect 241980 3062 242032 3068
rect 242808 3120 242860 3126
rect 242808 3062 242860 3068
rect 241518 2816 241574 2825
rect 241518 2751 241574 2760
rect 241992 480 242020 3062
rect 242912 626 242940 119954
rect 244372 118176 244424 118182
rect 244372 118118 244424 118124
rect 244384 115954 244412 118118
rect 244292 115938 244412 115954
rect 244280 115932 244412 115938
rect 244332 115926 244412 115932
rect 244280 115874 244332 115880
rect 244292 115843 244320 115874
rect 244280 106344 244332 106350
rect 244280 106286 244332 106292
rect 244292 96626 244320 106286
rect 244280 96620 244332 96626
rect 244280 96562 244332 96568
rect 244280 87032 244332 87038
rect 244280 86974 244332 86980
rect 244292 77178 244320 86974
rect 244280 77172 244332 77178
rect 244280 77114 244332 77120
rect 244280 67652 244332 67658
rect 244280 67594 244332 67600
rect 244292 57934 244320 67594
rect 244280 57928 244332 57934
rect 244280 57870 244332 57876
rect 244280 48340 244332 48346
rect 244280 48282 244332 48288
rect 244292 38622 244320 48282
rect 244280 38616 244332 38622
rect 244280 38558 244332 38564
rect 244280 29028 244332 29034
rect 244280 28970 244332 28976
rect 244292 19310 244320 28970
rect 244280 19304 244332 19310
rect 244280 19246 244332 19252
rect 245476 11552 245528 11558
rect 245476 11494 245528 11500
rect 244280 9716 244332 9722
rect 244280 9658 244332 9664
rect 244292 2938 244320 9658
rect 245488 9654 245516 11494
rect 245476 9648 245528 9654
rect 245476 9590 245528 9596
rect 245580 5370 245608 120022
rect 245672 12170 245700 122046
rect 248326 121952 248382 121961
rect 248326 121887 248382 121896
rect 246948 118924 247000 118930
rect 246948 118866 247000 118872
rect 245660 12164 245712 12170
rect 245660 12106 245712 12112
rect 245660 9648 245712 9654
rect 245660 9590 245712 9596
rect 245568 5364 245620 5370
rect 245568 5306 245620 5312
rect 245672 4842 245700 9590
rect 244200 2910 244320 2938
rect 245580 4814 245700 4842
rect 244200 2530 244228 2910
rect 244200 2502 244412 2530
rect 242912 598 243216 626
rect 243188 480 243216 598
rect 244384 480 244412 2502
rect 245580 480 245608 4814
rect 246960 626 246988 118866
rect 246776 598 246988 626
rect 248340 610 248368 121887
rect 249628 12034 249656 122046
rect 251088 120080 251140 120086
rect 251088 120022 251140 120028
rect 249708 118176 249760 118182
rect 249708 118118 249760 118124
rect 249616 12028 249668 12034
rect 249616 11970 249668 11976
rect 249720 3398 249748 118118
rect 251100 3398 251128 120022
rect 251192 12102 251220 122046
rect 251180 12096 251232 12102
rect 251180 12038 251232 12044
rect 251456 5024 251508 5030
rect 251456 4966 251508 4972
rect 249156 3392 249208 3398
rect 249156 3334 249208 3340
rect 249708 3392 249760 3398
rect 249708 3334 249760 3340
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 247960 604 248012 610
rect 246776 480 246804 598
rect 247960 546 248012 552
rect 248328 604 248380 610
rect 248328 546 248380 552
rect 247972 480 248000 546
rect 249168 480 249196 3334
rect 250364 480 250392 3334
rect 251468 480 251496 4966
rect 253860 3398 253888 122538
rect 259380 122233 259408 122606
rect 259366 122224 259422 122233
rect 259366 122159 259422 122168
rect 278686 122224 278742 122233
rect 278686 122159 278742 122168
rect 253952 122046 254058 122074
rect 256450 122046 256648 122074
rect 258842 122046 259408 122074
rect 253952 8226 253980 122046
rect 256620 14822 256648 122046
rect 258172 118584 258224 118590
rect 258172 118526 258224 118532
rect 258184 115954 258212 118526
rect 258092 115938 258212 115954
rect 258080 115932 258212 115938
rect 258132 115926 258212 115932
rect 258080 115874 258132 115880
rect 258092 115843 258120 115874
rect 258080 102944 258132 102950
rect 258080 102886 258132 102892
rect 258092 96626 258120 102886
rect 258080 96620 258132 96626
rect 258080 96562 258132 96568
rect 258080 87032 258132 87038
rect 258080 86974 258132 86980
rect 258092 77178 258120 86974
rect 258080 77172 258132 77178
rect 258080 77114 258132 77120
rect 258080 67652 258132 67658
rect 258080 67594 258132 67600
rect 258092 57934 258120 67594
rect 258080 57928 258132 57934
rect 258080 57870 258132 57876
rect 258080 48340 258132 48346
rect 258080 48282 258132 48288
rect 258092 38622 258120 48282
rect 258080 38616 258132 38622
rect 258080 38558 258132 38564
rect 258080 29028 258132 29034
rect 258080 28970 258132 28976
rect 258092 19310 258120 28970
rect 258080 19304 258132 19310
rect 258080 19246 258132 19252
rect 258264 19304 258316 19310
rect 258264 19246 258316 19252
rect 256608 14816 256660 14822
rect 256608 14758 256660 14764
rect 258276 9761 258304 19246
rect 259380 16046 259408 122046
rect 261220 120018 261248 122060
rect 261208 120012 261260 120018
rect 261208 119954 261260 119960
rect 262128 120012 262180 120018
rect 262128 119954 262180 119960
rect 259368 16040 259420 16046
rect 259368 15982 259420 15988
rect 258078 9752 258134 9761
rect 258078 9687 258134 9696
rect 258262 9752 258318 9761
rect 258262 9687 258318 9696
rect 258092 9654 258120 9687
rect 258080 9648 258132 9654
rect 258080 9590 258132 9596
rect 262140 8226 262168 119954
rect 263612 118726 263640 122060
rect 265820 120018 265848 122060
rect 265808 120012 265860 120018
rect 265808 119954 265860 119960
rect 268212 118794 268240 122060
rect 270604 119882 270632 122060
rect 270592 119876 270644 119882
rect 270592 119818 270644 119824
rect 272996 118810 273024 122060
rect 273166 120864 273222 120873
rect 273166 120799 273222 120808
rect 268200 118788 268252 118794
rect 272996 118782 273116 118810
rect 268200 118730 268252 118736
rect 263600 118720 263652 118726
rect 263600 118662 263652 118668
rect 267740 118516 267792 118522
rect 267740 118458 267792 118464
rect 266082 111208 266138 111217
rect 263600 111172 263652 111178
rect 266082 111143 266138 111152
rect 263600 111114 263652 111120
rect 253940 8220 253992 8226
rect 253940 8162 253992 8168
rect 262128 8220 262180 8226
rect 262128 8162 262180 8168
rect 261024 6588 261076 6594
rect 261024 6530 261076 6536
rect 256240 5500 256292 5506
rect 256240 5442 256292 5448
rect 252652 3392 252704 3398
rect 252652 3334 252704 3340
rect 253848 3392 253900 3398
rect 253848 3334 253900 3340
rect 252664 480 252692 3334
rect 255044 3188 255096 3194
rect 255044 3130 255096 3136
rect 253846 3088 253902 3097
rect 253846 3023 253902 3032
rect 253860 480 253888 3023
rect 255056 480 255084 3130
rect 256252 480 256280 5442
rect 257434 3768 257490 3777
rect 257434 3703 257490 3712
rect 259826 3768 259882 3777
rect 259826 3703 259882 3712
rect 257448 480 257476 3703
rect 259366 3632 259422 3641
rect 259366 3567 259422 3576
rect 259380 2825 259408 3567
rect 259366 2816 259422 2825
rect 259366 2751 259422 2760
rect 258632 604 258684 610
rect 258632 546 258684 552
rect 258644 480 258672 546
rect 259840 480 259868 3703
rect 261036 480 261064 6530
rect 262220 5092 262272 5098
rect 262220 5034 262272 5040
rect 262232 480 262260 5034
rect 263414 3904 263470 3913
rect 263414 3839 263470 3848
rect 263428 480 263456 3839
rect 263612 3346 263640 111114
rect 266096 102202 266124 111143
rect 266084 102196 266136 102202
rect 266084 102138 266136 102144
rect 266268 102196 266320 102202
rect 266268 102138 266320 102144
rect 263612 3318 264652 3346
rect 264624 480 264652 3318
rect 266280 3262 266308 102138
rect 267002 5264 267058 5273
rect 267002 5199 267058 5208
rect 265808 3256 265860 3262
rect 265808 3198 265860 3204
rect 266268 3256 266320 3262
rect 266268 3198 266320 3204
rect 265820 480 265848 3198
rect 267016 480 267044 5199
rect 267752 3482 267780 118458
rect 269120 118448 269172 118454
rect 269120 118390 269172 118396
rect 269132 3482 269160 118390
rect 273088 114578 273116 118782
rect 272984 114572 273036 114578
rect 272984 114514 273036 114520
rect 273076 114572 273128 114578
rect 273076 114514 273128 114520
rect 272996 109206 273024 114514
rect 272984 109200 273036 109206
rect 272984 109142 273036 109148
rect 272892 108928 272944 108934
rect 272892 108870 272944 108876
rect 272904 106185 272932 108870
rect 272614 106176 272670 106185
rect 272614 106111 272670 106120
rect 272890 106176 272946 106185
rect 272890 106111 272946 106120
rect 272628 99278 272656 106111
rect 272616 99272 272668 99278
rect 272616 99214 272668 99220
rect 272984 99272 273036 99278
rect 272984 99214 273036 99220
rect 272996 96626 273024 99214
rect 272984 96620 273036 96626
rect 272984 96562 273036 96568
rect 272984 87032 273036 87038
rect 272984 86974 273036 86980
rect 272996 80170 273024 86974
rect 272984 80164 273036 80170
rect 272984 80106 273036 80112
rect 272984 80028 273036 80034
rect 272984 79970 273036 79976
rect 272996 70394 273024 79970
rect 272904 70366 273024 70394
rect 272904 70258 272932 70366
rect 272904 70230 273024 70258
rect 272996 51082 273024 70230
rect 272904 51066 273024 51082
rect 272892 51060 273024 51066
rect 272944 51054 273024 51060
rect 273076 51060 273128 51066
rect 272892 51002 272944 51008
rect 273076 51002 273128 51008
rect 272904 50971 272932 51002
rect 273088 48278 273116 51002
rect 273076 48272 273128 48278
rect 273076 48214 273128 48220
rect 272984 38684 273036 38690
rect 272984 38626 273036 38632
rect 272996 31770 273024 38626
rect 272904 31742 273024 31770
rect 272904 26874 272932 31742
rect 272904 26846 273024 26874
rect 272996 22114 273024 26846
rect 272996 22098 273116 22114
rect 272892 22092 272944 22098
rect 272996 22092 273128 22098
rect 272996 22086 273076 22092
rect 272892 22034 272944 22040
rect 273076 22034 273128 22040
rect 272904 14754 272932 22034
rect 272892 14748 272944 14754
rect 272892 14690 272944 14696
rect 271510 4040 271566 4049
rect 271510 3975 271566 3984
rect 271694 4040 271750 4049
rect 271694 3975 271750 3984
rect 270498 3768 270554 3777
rect 270498 3703 270554 3712
rect 267752 3454 268148 3482
rect 269132 3454 269344 3482
rect 268120 480 268148 3454
rect 269316 480 269344 3454
rect 270512 480 270540 3703
rect 271524 3097 271552 3975
rect 271510 3088 271566 3097
rect 271510 3023 271566 3032
rect 271708 480 271736 3975
rect 273180 3482 273208 120799
rect 274548 120692 274600 120698
rect 274548 120634 274600 120640
rect 272904 3454 273208 3482
rect 272904 480 272932 3454
rect 274560 3262 274588 120634
rect 275388 119882 275416 122060
rect 277780 121582 277808 122060
rect 278700 121825 278728 122159
rect 278686 121816 278742 121825
rect 278686 121751 278742 121760
rect 277768 121576 277820 121582
rect 277768 121518 277820 121524
rect 275376 119876 275428 119882
rect 275376 119818 275428 119824
rect 280172 118794 280200 122060
rect 281552 122046 282578 122074
rect 280160 118788 280212 118794
rect 280160 118730 280212 118736
rect 278688 115456 278740 115462
rect 278688 115398 278740 115404
rect 276018 111208 276074 111217
rect 276018 111143 276020 111152
rect 276072 111143 276074 111152
rect 276020 111114 276072 111120
rect 275282 4040 275338 4049
rect 275282 3975 275338 3984
rect 274088 3256 274140 3262
rect 274088 3198 274140 3204
rect 274548 3256 274600 3262
rect 274548 3198 274600 3204
rect 274100 480 274128 3198
rect 275296 480 275324 3975
rect 278700 3262 278728 115398
rect 281264 6520 281316 6526
rect 281264 6462 281316 6468
rect 278870 4040 278926 4049
rect 278870 3975 278926 3984
rect 277676 3256 277728 3262
rect 277676 3198 277728 3204
rect 278688 3256 278740 3262
rect 278688 3198 278740 3204
rect 276480 3188 276532 3194
rect 276480 3130 276532 3136
rect 276492 480 276520 3130
rect 277688 480 277716 3198
rect 278884 480 278912 3975
rect 280066 3088 280122 3097
rect 280066 3023 280122 3032
rect 280080 480 280108 3023
rect 281276 480 281304 6462
rect 281552 5234 281580 122046
rect 281540 5228 281592 5234
rect 281540 5170 281592 5176
rect 282458 5128 282514 5137
rect 282458 5063 282514 5072
rect 282472 480 282500 5063
rect 284220 3398 284248 122606
rect 284956 120630 284984 122060
rect 284944 120624 284996 120630
rect 284944 120566 284996 120572
rect 285494 111208 285550 111217
rect 285494 111143 285496 111152
rect 285548 111143 285550 111152
rect 285496 111114 285548 111120
rect 284300 13252 284352 13258
rect 284300 13194 284352 13200
rect 283656 3392 283708 3398
rect 283656 3334 283708 3340
rect 284208 3392 284260 3398
rect 284208 3334 284260 3340
rect 283668 480 283696 3334
rect 284312 626 284340 13194
rect 286980 3398 287008 122674
rect 500144 122641 500172 122726
rect 500512 122641 500540 122726
rect 500130 122632 500186 122641
rect 500130 122567 500186 122576
rect 500314 122632 500370 122641
rect 500314 122567 500370 122576
rect 500498 122632 500554 122641
rect 500498 122567 500554 122576
rect 365628 122528 365680 122534
rect 365628 122470 365680 122476
rect 298006 122224 298062 122233
rect 298006 122159 298062 122168
rect 318614 122224 318670 122233
rect 318798 122224 318854 122233
rect 318670 122182 318798 122210
rect 318614 122159 318670 122168
rect 318798 122159 318854 122168
rect 336646 122224 336702 122233
rect 355966 122224 356022 122233
rect 351762 122182 351960 122210
rect 336646 122159 336702 122168
rect 287164 122046 287362 122074
rect 289648 122046 289754 122074
rect 291304 122046 292146 122074
rect 294538 122046 295288 122074
rect 287060 118380 287112 118386
rect 287060 118322 287112 118328
rect 287072 7546 287100 118322
rect 287164 9314 287192 122046
rect 289544 96620 289596 96626
rect 289544 96562 289596 96568
rect 289556 87009 289584 96562
rect 289542 87000 289598 87009
rect 289542 86935 289598 86944
rect 289544 57928 289596 57934
rect 289544 57870 289596 57876
rect 289556 53922 289584 57870
rect 289544 53916 289596 53922
rect 289544 53858 289596 53864
rect 289648 48482 289676 122046
rect 289726 119912 289782 119921
rect 289726 119847 289782 119856
rect 289740 97073 289768 119847
rect 289726 97064 289782 97073
rect 289726 96999 289782 97008
rect 289726 96656 289782 96665
rect 289726 96591 289728 96600
rect 289780 96591 289782 96600
rect 289728 96562 289780 96568
rect 289726 87000 289782 87009
rect 289726 86935 289782 86944
rect 289740 77586 289768 86935
rect 289728 77580 289780 77586
rect 289728 77522 289780 77528
rect 289728 77308 289780 77314
rect 289728 77250 289780 77256
rect 289740 57934 289768 77250
rect 289728 57928 289780 57934
rect 289728 57870 289780 57876
rect 289728 53916 289780 53922
rect 289728 53858 289780 53864
rect 289636 48476 289688 48482
rect 289636 48418 289688 48424
rect 289636 48272 289688 48278
rect 289636 48214 289688 48220
rect 289648 13258 289676 48214
rect 289740 46918 289768 53858
rect 289728 46912 289780 46918
rect 289728 46854 289780 46860
rect 289728 37324 289780 37330
rect 289728 37266 289780 37272
rect 289740 27606 289768 37266
rect 289728 27600 289780 27606
rect 289728 27542 289780 27548
rect 289636 13252 289688 13258
rect 289636 13194 289688 13200
rect 289728 12504 289780 12510
rect 289728 12446 289780 12452
rect 287152 9308 287204 9314
rect 287152 9250 287204 9256
rect 289740 8265 289768 12446
rect 290738 8936 290794 8945
rect 290738 8871 290794 8880
rect 289726 8256 289782 8265
rect 289726 8191 289782 8200
rect 289910 8256 289966 8265
rect 289910 8191 289966 8200
rect 287060 7540 287112 7546
rect 287060 7482 287112 7488
rect 288348 7540 288400 7546
rect 288348 7482 288400 7488
rect 285956 3392 286008 3398
rect 285956 3334 286008 3340
rect 286968 3392 287020 3398
rect 286968 3334 287020 3340
rect 284312 598 284800 626
rect 284772 480 284800 598
rect 285968 480 285996 3334
rect 287152 3256 287204 3262
rect 287152 3198 287204 3204
rect 287164 480 287192 3198
rect 288360 480 288388 7482
rect 289924 610 289952 8191
rect 289544 604 289596 610
rect 289544 546 289596 552
rect 289912 604 289964 610
rect 289912 546 289964 552
rect 289556 480 289584 546
rect 290752 480 290780 8871
rect 291304 3330 291332 122046
rect 293868 15972 293920 15978
rect 293868 15914 293920 15920
rect 291936 5228 291988 5234
rect 291936 5170 291988 5176
rect 291292 3324 291344 3330
rect 291292 3266 291344 3272
rect 291948 480 291976 5170
rect 293880 3398 293908 15914
rect 295260 14890 295288 122046
rect 296732 122046 296930 122074
rect 296626 119232 296682 119241
rect 296626 119167 296682 119176
rect 295340 111240 295392 111246
rect 295338 111208 295340 111217
rect 295392 111208 295394 111217
rect 295338 111143 295394 111152
rect 295248 14884 295300 14890
rect 295248 14826 295300 14832
rect 294328 5432 294380 5438
rect 294328 5374 294380 5380
rect 293132 3392 293184 3398
rect 293132 3334 293184 3340
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 293144 480 293172 3334
rect 294340 480 294368 5374
rect 296640 3398 296668 119167
rect 296732 5506 296760 122046
rect 298020 121689 298048 122159
rect 298006 121680 298062 121689
rect 298006 121615 298062 121624
rect 299308 99482 299336 122060
rect 301700 118998 301728 122060
rect 301688 118992 301740 118998
rect 301688 118934 301740 118940
rect 304092 118862 304120 122060
rect 304908 120556 304960 120562
rect 304908 120498 304960 120504
rect 304080 118856 304132 118862
rect 304080 118798 304132 118804
rect 304920 111314 304948 120498
rect 306484 119746 306512 122060
rect 307772 122046 308890 122074
rect 306472 119740 306524 119746
rect 306472 119682 306524 119688
rect 307024 118720 307076 118726
rect 307024 118662 307076 118668
rect 305000 118312 305052 118318
rect 305000 118254 305052 118260
rect 304908 111308 304960 111314
rect 304908 111250 304960 111256
rect 304816 111240 304868 111246
rect 304906 111208 304962 111217
rect 304868 111188 304906 111194
rect 304816 111182 304906 111188
rect 304828 111166 304906 111182
rect 304906 111143 304962 111152
rect 304908 105528 304960 105534
rect 304908 105470 304960 105476
rect 299296 99476 299348 99482
rect 299296 99418 299348 99424
rect 299296 99340 299348 99346
rect 299296 99282 299348 99288
rect 299308 96626 299336 99282
rect 299296 96620 299348 96626
rect 299296 96562 299348 96568
rect 299296 87032 299348 87038
rect 299296 86974 299348 86980
rect 299308 80170 299336 86974
rect 299296 80164 299348 80170
rect 299296 80106 299348 80112
rect 299296 80028 299348 80034
rect 299296 79970 299348 79976
rect 299308 70394 299336 79970
rect 299216 70366 299336 70394
rect 299216 70258 299244 70366
rect 299216 70230 299336 70258
rect 299308 51082 299336 70230
rect 299216 51066 299336 51082
rect 299204 51060 299336 51066
rect 299256 51054 299336 51060
rect 299388 51060 299440 51066
rect 299204 51002 299256 51008
rect 299388 51002 299440 51008
rect 299216 50971 299244 51002
rect 299400 48278 299428 51002
rect 299388 48272 299440 48278
rect 299388 48214 299440 48220
rect 299296 38684 299348 38690
rect 299296 38626 299348 38632
rect 299308 33810 299336 38626
rect 299032 33782 299336 33810
rect 299032 29050 299060 33782
rect 299032 29022 299152 29050
rect 299124 27606 299152 29022
rect 299112 27600 299164 27606
rect 299112 27542 299164 27548
rect 297914 19136 297970 19145
rect 297914 19071 297970 19080
rect 296720 5500 296772 5506
rect 296720 5442 296772 5448
rect 297824 5500 297876 5506
rect 297824 5442 297876 5448
rect 295524 3392 295576 3398
rect 295524 3334 295576 3340
rect 296628 3392 296680 3398
rect 296628 3334 296680 3340
rect 295536 480 295564 3334
rect 296720 3052 296772 3058
rect 296720 2994 296772 3000
rect 296732 480 296760 2994
rect 297836 2802 297864 5442
rect 297928 3058 297956 19071
rect 299204 18012 299256 18018
rect 299204 17954 299256 17960
rect 299216 6526 299244 17954
rect 302240 14884 302292 14890
rect 302240 14826 302292 14832
rect 299204 6520 299256 6526
rect 299204 6462 299256 6468
rect 300308 5432 300360 5438
rect 300308 5374 300360 5380
rect 298006 3632 298062 3641
rect 298006 3567 298062 3576
rect 298020 3097 298048 3567
rect 299110 3224 299166 3233
rect 299110 3159 299166 3168
rect 298006 3088 298062 3097
rect 297916 3052 297968 3058
rect 298006 3023 298062 3032
rect 297916 2994 297968 3000
rect 297836 2774 297956 2802
rect 297928 480 297956 2774
rect 299124 480 299152 3159
rect 300320 480 300348 5374
rect 301410 3224 301466 3233
rect 301410 3159 301466 3168
rect 301424 480 301452 3159
rect 302252 626 302280 14826
rect 304920 3398 304948 105470
rect 303804 3392 303856 3398
rect 303804 3334 303856 3340
rect 304908 3392 304960 3398
rect 304908 3334 304960 3340
rect 302252 598 302648 626
rect 302620 480 302648 598
rect 303816 480 303844 3334
rect 305012 1290 305040 118254
rect 307036 3330 307064 118662
rect 307772 3398 307800 122046
rect 311084 119746 311112 122060
rect 313476 120766 313504 122060
rect 313464 120760 313516 120766
rect 313464 120702 313516 120708
rect 311072 119740 311124 119746
rect 311072 119682 311124 119688
rect 313924 118992 313976 118998
rect 313924 118934 313976 118940
rect 310520 118788 310572 118794
rect 310520 118730 310572 118736
rect 309140 10600 309192 10606
rect 309140 10542 309192 10548
rect 308588 9240 308640 9246
rect 308588 9182 308640 9188
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307024 3324 307076 3330
rect 307024 3266 307076 3272
rect 307392 3324 307444 3330
rect 307392 3266 307444 3272
rect 305092 3188 305144 3194
rect 305092 3130 305144 3136
rect 305000 1284 305052 1290
rect 305000 1226 305052 1232
rect 305104 1170 305132 3130
rect 306196 1284 306248 1290
rect 306196 1226 306248 1232
rect 305012 1142 305132 1170
rect 305012 480 305040 1142
rect 306208 480 306236 1226
rect 307404 480 307432 3266
rect 308600 480 308628 9182
rect 309152 3346 309180 10542
rect 310532 3346 310560 118730
rect 313280 14816 313332 14822
rect 313280 14758 313332 14764
rect 312176 5160 312228 5166
rect 312176 5102 312228 5108
rect 309152 3318 309824 3346
rect 310532 3318 311020 3346
rect 309796 480 309824 3318
rect 310992 480 311020 3318
rect 312188 480 312216 5102
rect 313292 1578 313320 14758
rect 313936 3806 313964 118934
rect 315868 118726 315896 122060
rect 318260 120766 318288 122060
rect 318248 120760 318300 120766
rect 318248 120702 318300 120708
rect 320652 120057 320680 122060
rect 325450 122046 325648 122074
rect 322846 121816 322902 121825
rect 322846 121751 322902 121760
rect 320638 120048 320694 120057
rect 320638 119983 320694 119992
rect 317326 119096 317382 119105
rect 317326 119031 317382 119040
rect 315856 118720 315908 118726
rect 315856 118662 315908 118668
rect 314658 111208 314714 111217
rect 314658 111143 314660 111152
rect 314712 111143 314714 111152
rect 314660 111114 314712 111120
rect 315946 19136 316002 19145
rect 315946 19071 316002 19080
rect 314566 19000 314622 19009
rect 314566 18935 314622 18944
rect 313924 3800 313976 3806
rect 313924 3742 313976 3748
rect 313292 1550 313412 1578
rect 313384 480 313412 1550
rect 314580 480 314608 18935
rect 315960 18873 315988 19071
rect 315946 18864 316002 18873
rect 315946 18799 316002 18808
rect 315764 3800 315816 3806
rect 315764 3742 315816 3748
rect 315776 480 315804 3742
rect 317340 3482 317368 119031
rect 320180 118244 320232 118250
rect 320180 118186 320232 118192
rect 318062 5944 318118 5953
rect 318062 5879 318118 5888
rect 316972 3454 317368 3482
rect 316972 480 317000 3454
rect 318076 480 318104 5879
rect 318890 4176 318946 4185
rect 318812 4134 318890 4162
rect 318812 4049 318840 4134
rect 320192 4162 320220 118186
rect 322756 116816 322808 116822
rect 322756 116758 322808 116764
rect 320192 4134 320496 4162
rect 318890 4111 318946 4120
rect 318798 4040 318854 4049
rect 318798 3975 318854 3984
rect 319258 3768 319314 3777
rect 319258 3703 319314 3712
rect 319272 480 319300 3703
rect 320468 480 320496 4134
rect 322768 3398 322796 116758
rect 321652 3392 321704 3398
rect 321652 3334 321704 3340
rect 322756 3392 322808 3398
rect 322756 3334 322808 3340
rect 321664 480 321692 3334
rect 322860 480 322888 121751
rect 323582 111208 323638 111217
rect 323582 111143 323584 111152
rect 323636 111143 323638 111152
rect 323584 111114 323636 111120
rect 325620 12102 325648 122046
rect 326988 122052 327040 122058
rect 326988 121994 327040 122000
rect 327092 122046 327842 122074
rect 329852 122046 330234 122074
rect 325698 19136 325754 19145
rect 325698 19071 325754 19080
rect 325712 18873 325740 19071
rect 325698 18864 325754 18873
rect 325698 18799 325754 18808
rect 325608 12096 325660 12102
rect 325608 12038 325660 12044
rect 325238 6080 325294 6089
rect 325238 6015 325294 6024
rect 324044 3392 324096 3398
rect 324044 3334 324096 3340
rect 324056 480 324084 3334
rect 325252 480 325280 6015
rect 327000 3398 327028 121994
rect 327092 8158 327120 122046
rect 328366 121000 328422 121009
rect 328366 120935 328422 120944
rect 327080 8152 327132 8158
rect 327080 8094 327132 8100
rect 328380 3398 328408 120935
rect 329748 120488 329800 120494
rect 329748 120430 329800 120436
rect 328458 111480 328514 111489
rect 328458 111415 328514 111424
rect 328472 111217 328500 111415
rect 328458 111208 328514 111217
rect 328458 111143 328514 111152
rect 329760 3398 329788 120430
rect 329852 7886 329880 122046
rect 330944 121780 330996 121786
rect 330944 121722 330996 121728
rect 330956 121689 330984 121722
rect 330942 121680 330998 121689
rect 330942 121615 330998 121624
rect 332612 118998 332640 122060
rect 335018 122046 335308 122074
rect 332600 118992 332652 118998
rect 332600 118934 332652 118940
rect 331126 84824 331182 84833
rect 331126 84759 331182 84768
rect 329840 7880 329892 7886
rect 329840 7822 329892 7828
rect 331140 3398 331168 84759
rect 333980 14748 334032 14754
rect 333980 14690 334032 14696
rect 332508 13660 332560 13666
rect 332508 13602 332560 13608
rect 332520 3398 332548 13602
rect 333612 4752 333664 4758
rect 333612 4694 333664 4700
rect 332598 3632 332654 3641
rect 332598 3567 332654 3576
rect 326436 3392 326488 3398
rect 326436 3334 326488 3340
rect 326988 3392 327040 3398
rect 326988 3334 327040 3340
rect 327632 3392 327684 3398
rect 327632 3334 327684 3340
rect 328368 3392 328420 3398
rect 328368 3334 328420 3340
rect 328828 3392 328880 3398
rect 328828 3334 328880 3340
rect 329748 3392 329800 3398
rect 329748 3334 329800 3340
rect 330024 3392 330076 3398
rect 330024 3334 330076 3340
rect 331128 3392 331180 3398
rect 331128 3334 331180 3340
rect 331220 3392 331272 3398
rect 331220 3334 331272 3340
rect 332508 3392 332560 3398
rect 332508 3334 332560 3340
rect 326448 480 326476 3334
rect 327644 480 327672 3334
rect 328840 480 328868 3334
rect 330036 480 330064 3334
rect 331232 480 331260 3334
rect 332612 3097 332640 3567
rect 332598 3088 332654 3097
rect 332598 3023 332654 3032
rect 332414 2952 332470 2961
rect 332414 2887 332470 2896
rect 332428 480 332456 2887
rect 333624 480 333652 4694
rect 333992 3346 334020 14690
rect 335280 13598 335308 122046
rect 336660 121786 336688 122159
rect 336648 121780 336700 121786
rect 336648 121722 336700 121728
rect 337396 120902 337424 122060
rect 340892 122046 342194 122074
rect 338120 121848 338172 121854
rect 338118 121816 338120 121825
rect 338172 121816 338174 121825
rect 338118 121751 338174 121760
rect 338120 121712 338172 121718
rect 338120 121654 338172 121660
rect 337384 120896 337436 120902
rect 337384 120838 337436 120844
rect 335360 44872 335412 44878
rect 335360 44814 335412 44820
rect 335268 13592 335320 13598
rect 335268 13534 335320 13540
rect 335372 3754 335400 44814
rect 335910 19136 335966 19145
rect 335910 19071 335966 19080
rect 335924 18873 335952 19071
rect 335910 18864 335966 18873
rect 335910 18799 335966 18808
rect 337108 5160 337160 5166
rect 337108 5102 337160 5108
rect 335372 3726 335768 3754
rect 335358 3632 335414 3641
rect 335358 3567 335414 3576
rect 333992 3318 334756 3346
rect 334728 480 334756 3318
rect 335372 3097 335400 3567
rect 335740 3346 335768 3726
rect 335740 3318 335952 3346
rect 335358 3088 335414 3097
rect 335358 3023 335414 3032
rect 335924 480 335952 3318
rect 337120 480 337148 5102
rect 338132 3346 338160 121654
rect 340788 17536 340840 17542
rect 340788 17478 340840 17484
rect 340696 4072 340748 4078
rect 340696 4014 340748 4020
rect 339500 3392 339552 3398
rect 338132 3318 338344 3346
rect 339500 3334 339552 3340
rect 338316 480 338344 3318
rect 339512 480 339540 3334
rect 340708 480 340736 4014
rect 340800 3398 340828 17478
rect 340892 7954 340920 122046
rect 342996 121848 343048 121854
rect 342994 121816 342996 121825
rect 343048 121816 343050 121825
rect 342994 121751 343050 121760
rect 344572 118794 344600 122060
rect 346412 122046 346978 122074
rect 344560 118788 344612 118794
rect 344560 118730 344612 118736
rect 343546 111208 343602 111217
rect 343730 111208 343786 111217
rect 343602 111166 343730 111194
rect 343546 111143 343602 111152
rect 343730 111143 343786 111152
rect 345018 19136 345074 19145
rect 345018 19071 345074 19080
rect 345032 18873 345060 19071
rect 345018 18864 345074 18873
rect 345018 18799 345074 18808
rect 341892 9716 341944 9722
rect 341892 9658 341944 9664
rect 340880 7948 340932 7954
rect 340880 7890 340932 7896
rect 340788 3392 340840 3398
rect 340788 3334 340840 3340
rect 341904 480 341932 9658
rect 346412 7750 346440 122046
rect 349068 120896 349120 120902
rect 349068 120838 349120 120844
rect 348976 113892 349028 113898
rect 348976 113834 349028 113840
rect 346400 7744 346452 7750
rect 346400 7686 346452 7692
rect 345480 6656 345532 6662
rect 345480 6598 345532 6604
rect 343086 3768 343142 3777
rect 343086 3703 343142 3712
rect 343100 480 343128 3703
rect 344284 3392 344336 3398
rect 344284 3334 344336 3340
rect 344296 480 344324 3334
rect 345492 480 345520 6598
rect 346676 6588 346728 6594
rect 346676 6530 346728 6536
rect 346688 480 346716 6530
rect 348988 4078 349016 113834
rect 347872 4072 347924 4078
rect 347872 4014 347924 4020
rect 348976 4072 349028 4078
rect 348976 4014 349028 4020
rect 347884 480 347912 4014
rect 349080 480 349108 120838
rect 349160 119740 349212 119746
rect 349160 119682 349212 119688
rect 349172 12442 349200 119682
rect 349356 118726 349384 122060
rect 349344 118720 349396 118726
rect 349344 118662 349396 118668
rect 351932 104990 351960 122182
rect 355966 122159 356022 122168
rect 354154 122046 354628 122074
rect 352564 119740 352616 119746
rect 352564 119682 352616 119688
rect 351736 104984 351788 104990
rect 351736 104926 351788 104932
rect 351920 104984 351972 104990
rect 351920 104926 351972 104932
rect 351748 104854 351776 104926
rect 351736 104848 351788 104854
rect 351736 104790 351788 104796
rect 351736 89684 351788 89690
rect 351736 89626 351788 89632
rect 351748 80170 351776 89626
rect 351736 80164 351788 80170
rect 351736 80106 351788 80112
rect 351736 80028 351788 80034
rect 351736 79970 351788 79976
rect 351748 70394 351776 79970
rect 351656 70366 351776 70394
rect 351656 70258 351684 70366
rect 351656 70230 351776 70258
rect 351748 51082 351776 70230
rect 351656 51066 351776 51082
rect 351644 51060 351776 51066
rect 351696 51054 351776 51060
rect 351828 51060 351880 51066
rect 351644 51002 351696 51008
rect 351828 51002 351880 51008
rect 351656 50971 351684 51002
rect 351840 48278 351868 51002
rect 351828 48272 351880 48278
rect 351828 48214 351880 48220
rect 351736 38684 351788 38690
rect 351736 38626 351788 38632
rect 351748 31890 351776 38626
rect 351736 31884 351788 31890
rect 351736 31826 351788 31832
rect 351736 31748 351788 31754
rect 351736 31690 351788 31696
rect 351748 22114 351776 31690
rect 351748 22086 351868 22114
rect 351840 19310 351868 22086
rect 351828 19304 351880 19310
rect 351828 19246 351880 19252
rect 351920 14612 351972 14618
rect 351920 14554 351972 14560
rect 351932 12442 351960 14554
rect 349160 12436 349212 12442
rect 349160 12378 349212 12384
rect 350264 12436 350316 12442
rect 350264 12378 350316 12384
rect 351920 12436 351972 12442
rect 351920 12378 351972 12384
rect 352472 12436 352524 12442
rect 352472 12378 352524 12384
rect 350276 480 350304 12378
rect 351736 9784 351788 9790
rect 351736 9726 351788 9732
rect 351748 9654 351776 9726
rect 351736 9648 351788 9654
rect 351736 9590 351788 9596
rect 352484 4026 352512 12378
rect 352576 4146 352604 119682
rect 353298 111208 353354 111217
rect 353298 111143 353300 111152
rect 353352 111143 353354 111152
rect 353300 111114 353352 111120
rect 354600 10606 354628 122046
rect 355980 121689 356008 122159
rect 355966 121680 356022 121689
rect 355966 121615 356022 121624
rect 356348 119746 356376 122060
rect 357452 122046 358754 122074
rect 361146 122046 361528 122074
rect 356336 119740 356388 119746
rect 356336 119682 356388 119688
rect 355968 118992 356020 118998
rect 355968 118934 356020 118940
rect 355322 19136 355378 19145
rect 355322 19071 355378 19080
rect 355336 18873 355364 19071
rect 355322 18864 355378 18873
rect 355322 18799 355378 18808
rect 354588 10600 354640 10606
rect 354588 10542 354640 10548
rect 353758 8936 353814 8945
rect 353758 8871 353814 8880
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 352484 3998 352604 4026
rect 351368 3936 351420 3942
rect 351368 3878 351420 3884
rect 351380 480 351408 3878
rect 351826 3768 351882 3777
rect 351826 3703 351882 3712
rect 351840 3097 351868 3703
rect 351826 3088 351882 3097
rect 351826 3023 351882 3032
rect 352576 480 352604 3998
rect 353772 480 353800 8871
rect 355980 4146 356008 118934
rect 357348 7744 357400 7750
rect 357348 7686 357400 7692
rect 354956 4140 355008 4146
rect 354956 4082 355008 4088
rect 355968 4140 356020 4146
rect 355968 4082 356020 4088
rect 354968 480 354996 4082
rect 356794 4040 356850 4049
rect 357254 4040 357310 4049
rect 356850 3998 357254 4026
rect 356794 3975 356850 3984
rect 357254 3975 357310 3984
rect 356978 3904 357034 3913
rect 357254 3904 357310 3913
rect 357034 3862 357254 3890
rect 356978 3839 357034 3848
rect 357254 3839 357310 3848
rect 356152 3120 356204 3126
rect 356152 3062 356204 3068
rect 356164 480 356192 3062
rect 357360 480 357388 7686
rect 357452 5302 357480 122046
rect 360200 119060 360252 119066
rect 360200 119002 360252 119008
rect 358820 13388 358872 13394
rect 358820 13330 358872 13336
rect 358544 9172 358596 9178
rect 358544 9114 358596 9120
rect 357440 5296 357492 5302
rect 357440 5238 357492 5244
rect 358556 480 358584 9114
rect 358832 2854 358860 13330
rect 360212 12442 360240 119002
rect 361500 37330 361528 122046
rect 363524 119746 363552 122060
rect 363512 119740 363564 119746
rect 363512 119682 363564 119688
rect 362774 111208 362830 111217
rect 362774 111143 362776 111152
rect 362828 111143 362830 111152
rect 362776 111114 362828 111120
rect 361488 37324 361540 37330
rect 361488 37266 361540 37272
rect 362960 37324 363012 37330
rect 362960 37266 363012 37272
rect 362972 27606 363000 37266
rect 362960 27600 363012 27606
rect 362960 27542 363012 27548
rect 363236 27600 363288 27606
rect 363236 27542 363288 27548
rect 360200 12436 360252 12442
rect 360200 12378 360252 12384
rect 360936 12436 360988 12442
rect 360936 12378 360988 12384
rect 358820 2848 358872 2854
rect 358820 2790 358872 2796
rect 359740 2780 359792 2786
rect 359740 2722 359792 2728
rect 359752 480 359780 2722
rect 360948 480 360976 12378
rect 363248 4842 363276 27542
rect 364338 19136 364394 19145
rect 364338 19071 364394 19080
rect 364352 18873 364380 19071
rect 364338 18864 364394 18873
rect 364338 18799 364394 18808
rect 363248 4814 363368 4842
rect 362132 4684 362184 4690
rect 362132 4626 362184 4632
rect 362144 480 362172 4626
rect 363340 480 363368 4814
rect 365640 4146 365668 122470
rect 376772 122318 376892 122346
rect 376772 122233 376800 122318
rect 375286 122224 375342 122233
rect 375286 122159 375342 122168
rect 376758 122224 376814 122233
rect 376758 122159 376814 122168
rect 365916 119338 365944 122060
rect 367008 122052 367060 122058
rect 367008 121994 367060 122000
rect 365904 119332 365956 119338
rect 365904 119274 365956 119280
rect 365720 14680 365772 14686
rect 365720 14622 365772 14628
rect 365732 7546 365760 14622
rect 365720 7540 365772 7546
rect 365720 7482 365772 7488
rect 366916 7540 366968 7546
rect 366916 7482 366968 7488
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 365628 4140 365680 4146
rect 365628 4082 365680 4088
rect 365720 4140 365772 4146
rect 365720 4082 365772 4088
rect 364536 480 364564 4082
rect 365732 480 365760 4082
rect 366928 480 366956 7482
rect 367020 4146 367048 121994
rect 368308 118726 368336 122060
rect 370714 122046 371188 122074
rect 368296 118720 368348 118726
rect 368296 118662 368348 118668
rect 369952 118720 370004 118726
rect 369952 118662 370004 118668
rect 367100 14544 367152 14550
rect 367100 14486 367152 14492
rect 367112 12442 367140 14486
rect 369964 12510 369992 118662
rect 371160 13394 371188 122046
rect 373092 119338 373120 122060
rect 375300 121689 375328 122159
rect 375286 121680 375342 121689
rect 375286 121615 375342 121624
rect 373080 119332 373132 119338
rect 373080 119274 373132 119280
rect 373908 119332 373960 119338
rect 373908 119274 373960 119280
rect 371330 116784 371386 116793
rect 371330 116719 371386 116728
rect 372528 116748 372580 116754
rect 371344 115954 371372 116719
rect 372528 116690 372580 116696
rect 371252 115926 371372 115954
rect 372540 115954 372568 116690
rect 372540 115926 372660 115954
rect 371148 13388 371200 13394
rect 371148 13330 371200 13336
rect 371252 12510 371280 115926
rect 372632 12510 372660 115926
rect 372712 111240 372764 111246
rect 372710 111208 372712 111217
rect 372764 111208 372766 111217
rect 372710 111143 372766 111152
rect 369952 12504 370004 12510
rect 369952 12446 370004 12452
rect 371240 12504 371292 12510
rect 371240 12446 371292 12452
rect 372620 12504 372672 12510
rect 372620 12446 372672 12452
rect 367100 12436 367152 12442
rect 367100 12378 367152 12384
rect 368020 12436 368072 12442
rect 368020 12378 368072 12384
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 368032 480 368060 12378
rect 370412 12368 370464 12374
rect 370412 12310 370464 12316
rect 371608 12368 371660 12374
rect 371608 12310 371660 12316
rect 372804 12368 372856 12374
rect 372804 12310 372856 12316
rect 369214 10568 369270 10577
rect 369214 10503 369270 10512
rect 369228 480 369256 10503
rect 370424 9654 370452 12310
rect 371620 9654 371648 12310
rect 372816 9654 372844 12310
rect 370412 9648 370464 9654
rect 370412 9590 370464 9596
rect 371608 9648 371660 9654
rect 371608 9590 371660 9596
rect 372804 9648 372856 9654
rect 372804 9590 372856 9596
rect 373920 5302 373948 119274
rect 375484 118930 375512 122060
rect 376864 121990 376892 122318
rect 404372 122318 404492 122346
rect 404372 122233 404400 122318
rect 386142 122224 386198 122233
rect 386142 122159 386198 122168
rect 404358 122224 404414 122233
rect 404358 122159 404414 122168
rect 376852 121984 376904 121990
rect 376852 121926 376904 121932
rect 377876 121582 377904 122060
rect 377864 121576 377916 121582
rect 377864 121518 377916 121524
rect 380268 119338 380296 122060
rect 382660 119610 382688 122060
rect 382648 119604 382700 119610
rect 382648 119546 382700 119552
rect 380256 119332 380308 119338
rect 380256 119274 380308 119280
rect 384948 119060 385000 119066
rect 384948 119002 385000 119008
rect 375472 118924 375524 118930
rect 375472 118866 375524 118872
rect 375286 115424 375342 115433
rect 375286 115359 375342 115368
rect 375196 14544 375248 14550
rect 375196 14486 375248 14492
rect 373908 5296 373960 5302
rect 373908 5238 373960 5244
rect 375208 4146 375236 14486
rect 374000 4140 374052 4146
rect 374000 4082 374052 4088
rect 375196 4140 375248 4146
rect 375196 4082 375248 4088
rect 370412 604 370464 610
rect 370412 546 370464 552
rect 371608 604 371660 610
rect 371608 546 371660 552
rect 372804 604 372856 610
rect 372804 546 372856 552
rect 370424 480 370452 546
rect 371620 480 371648 546
rect 372816 480 372844 546
rect 374012 480 374040 4082
rect 375300 4026 375328 115359
rect 382096 111240 382148 111246
rect 382094 111208 382096 111217
rect 382148 111208 382150 111217
rect 382094 111143 382150 111152
rect 378138 111072 378194 111081
rect 378138 111007 378140 111016
rect 378192 111007 378194 111016
rect 378140 110978 378192 110984
rect 378140 95260 378192 95266
rect 378140 95202 378192 95208
rect 378152 85542 378180 95202
rect 378140 85536 378192 85542
rect 378140 85478 378192 85484
rect 378140 75948 378192 75954
rect 378140 75890 378192 75896
rect 378152 66230 378180 75890
rect 378140 66224 378192 66230
rect 378140 66166 378192 66172
rect 378140 56636 378192 56642
rect 378140 56578 378192 56584
rect 378152 46918 378180 56578
rect 378140 46912 378192 46918
rect 378140 46854 378192 46860
rect 378140 37324 378192 37330
rect 378140 37266 378192 37272
rect 378152 27606 378180 37266
rect 378140 27600 378192 27606
rect 378140 27542 378192 27548
rect 378782 19136 378838 19145
rect 378782 19071 378838 19080
rect 383658 19136 383714 19145
rect 383658 19071 383714 19080
rect 378796 18873 378824 19071
rect 383672 18873 383700 19071
rect 378782 18864 378838 18873
rect 378782 18799 378838 18808
rect 383658 18864 383714 18873
rect 383658 18799 383714 18808
rect 378140 18012 378192 18018
rect 378140 17954 378192 17960
rect 377680 13184 377732 13190
rect 377680 13126 377732 13132
rect 377692 12322 377720 13126
rect 378152 12510 378180 17954
rect 378140 12504 378192 12510
rect 378140 12446 378192 12452
rect 377600 12294 377720 12322
rect 378784 12368 378836 12374
rect 378784 12310 378836 12316
rect 377600 9654 377628 12294
rect 378796 9654 378824 12310
rect 383568 10464 383620 10470
rect 383568 10406 383620 10412
rect 377588 9648 377640 9654
rect 377588 9590 377640 9596
rect 378784 9648 378836 9654
rect 378784 9590 378836 9596
rect 382372 6792 382424 6798
rect 382372 6734 382424 6740
rect 376392 6724 376444 6730
rect 376392 6666 376444 6672
rect 375208 3998 375328 4026
rect 375208 480 375236 3998
rect 376404 480 376432 6666
rect 379980 4616 380032 4622
rect 379980 4558 380032 4564
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 378784 604 378836 610
rect 378784 546 378836 552
rect 377600 480 377628 546
rect 378796 480 378824 546
rect 379992 480 380020 4558
rect 381176 4140 381228 4146
rect 381176 4082 381228 4088
rect 381188 480 381216 4082
rect 382384 480 382412 6734
rect 383580 480 383608 10406
rect 384960 2854 384988 119002
rect 385052 4690 385080 122060
rect 386156 121990 386184 122159
rect 400128 122120 400180 122126
rect 386432 122046 387458 122074
rect 386144 121984 386196 121990
rect 386144 121926 386196 121932
rect 386432 13530 386460 122046
rect 389836 120057 389864 122060
rect 392228 121106 392256 122060
rect 393964 121984 394016 121990
rect 393964 121926 394016 121932
rect 392216 121100 392268 121106
rect 392216 121042 392268 121048
rect 393228 120420 393280 120426
rect 393228 120362 393280 120368
rect 389638 120048 389694 120057
rect 389638 119983 389694 119992
rect 389822 120048 389878 120057
rect 389822 119983 389878 119992
rect 389652 118697 389680 119983
rect 391848 119604 391900 119610
rect 391848 119546 391900 119552
rect 389638 118688 389694 118697
rect 389638 118623 389694 118632
rect 386510 111208 386566 111217
rect 386510 111143 386566 111152
rect 386524 110945 386552 111143
rect 386510 110936 386566 110945
rect 386510 110871 386566 110880
rect 386420 13524 386472 13530
rect 386420 13466 386472 13472
rect 387062 6896 387118 6905
rect 387062 6831 387118 6840
rect 385040 4684 385092 4690
rect 385040 4626 385092 4632
rect 385868 3936 385920 3942
rect 385868 3878 385920 3884
rect 384672 2848 384724 2854
rect 384672 2790 384724 2796
rect 384948 2848 385000 2854
rect 384948 2790 385000 2796
rect 384684 480 384712 2790
rect 385880 480 385908 3878
rect 387076 480 387104 6831
rect 390650 6760 390706 6769
rect 390650 6695 390706 6704
rect 389454 6624 389510 6633
rect 389454 6559 389510 6568
rect 387800 4956 387852 4962
rect 387800 4898 387852 4904
rect 387812 3126 387840 4898
rect 388260 3392 388312 3398
rect 388260 3334 388312 3340
rect 387800 3120 387852 3126
rect 387800 3062 387852 3068
rect 388272 480 388300 3334
rect 389468 480 389496 6559
rect 390664 480 390692 6695
rect 391860 480 391888 119546
rect 393240 12578 393268 120362
rect 393320 115184 393372 115190
rect 393320 115126 393372 115132
rect 393228 12572 393280 12578
rect 393228 12514 393280 12520
rect 393044 9716 393096 9722
rect 393044 9658 393096 9664
rect 393056 480 393084 9658
rect 393332 3738 393360 115126
rect 393976 8106 394004 121926
rect 394620 115190 394648 122060
rect 396184 122046 397026 122074
rect 400128 122062 400180 122068
rect 396080 119128 396132 119134
rect 396080 119070 396132 119076
rect 394608 115184 394660 115190
rect 394608 115126 394660 115132
rect 393884 8078 394004 8106
rect 393884 3738 393912 8078
rect 395436 6860 395488 6866
rect 395436 6802 395488 6808
rect 394240 5364 394292 5370
rect 394240 5306 394292 5312
rect 393320 3732 393372 3738
rect 393320 3674 393372 3680
rect 393872 3732 393924 3738
rect 393872 3674 393924 3680
rect 394252 480 394280 5306
rect 394606 4176 394662 4185
rect 394606 4111 394662 4120
rect 394620 3777 394648 4111
rect 394606 3768 394662 3777
rect 394606 3703 394662 3712
rect 395448 480 395476 6802
rect 396092 610 396120 119070
rect 396184 7682 396212 122046
rect 399404 121650 399432 122060
rect 399392 121644 399444 121650
rect 399392 121586 399444 121592
rect 398748 118244 398800 118250
rect 398748 118186 398800 118192
rect 396172 7676 396224 7682
rect 396172 7618 396224 7624
rect 398760 3670 398788 118186
rect 400140 3670 400168 122062
rect 401612 120358 401640 122060
rect 402992 122046 404018 122074
rect 401600 120352 401652 120358
rect 401600 120294 401652 120300
rect 402244 119128 402296 119134
rect 402244 119070 402296 119076
rect 401508 116748 401560 116754
rect 401508 116690 401560 116696
rect 400220 8220 400272 8226
rect 400220 8162 400272 8168
rect 397828 3664 397880 3670
rect 397828 3606 397880 3612
rect 398748 3664 398800 3670
rect 398748 3606 398800 3612
rect 399024 3664 399076 3670
rect 399024 3606 399076 3612
rect 400128 3664 400180 3670
rect 400128 3606 400180 3612
rect 396080 604 396132 610
rect 396080 546 396132 552
rect 396632 604 396684 610
rect 396632 546 396684 552
rect 396644 480 396672 546
rect 397840 480 397868 3606
rect 399036 480 399064 3606
rect 400232 480 400260 8162
rect 400862 3768 400918 3777
rect 400862 3703 400918 3712
rect 400876 3097 400904 3703
rect 400862 3088 400918 3097
rect 400862 3023 400918 3032
rect 401520 626 401548 116690
rect 401690 111208 401746 111217
rect 401690 111143 401746 111152
rect 401704 110673 401732 111143
rect 401690 110664 401746 110673
rect 401690 110599 401746 110608
rect 401600 16040 401652 16046
rect 401600 15982 401652 15988
rect 401612 7682 401640 15982
rect 401600 7676 401652 7682
rect 401600 7618 401652 7624
rect 402256 3126 402284 119070
rect 402992 7750 403020 122046
rect 404464 121990 404492 122318
rect 413926 122224 413982 122233
rect 413926 122159 413982 122168
rect 415490 122224 415546 122233
rect 424966 122224 425022 122233
rect 415546 122182 415808 122210
rect 415490 122159 415546 122168
rect 405752 122046 406410 122074
rect 408512 122046 408802 122074
rect 404452 121984 404504 121990
rect 404452 121926 404504 121932
rect 405752 14550 405780 122046
rect 407028 118924 407080 118930
rect 407028 118866 407080 118872
rect 405740 14544 405792 14550
rect 405740 14486 405792 14492
rect 404912 10396 404964 10402
rect 404912 10338 404964 10344
rect 402980 7744 403032 7750
rect 402980 7686 403032 7692
rect 402520 7676 402572 7682
rect 402520 7618 402572 7624
rect 402244 3120 402296 3126
rect 402244 3062 402296 3068
rect 401336 598 401548 626
rect 401336 480 401364 598
rect 402532 480 402560 7618
rect 403714 6624 403770 6633
rect 403714 6559 403770 6568
rect 403728 480 403756 6559
rect 404924 480 404952 10338
rect 405648 4208 405700 4214
rect 405648 4150 405700 4156
rect 405660 3777 405688 4150
rect 405646 3768 405702 3777
rect 405646 3703 405702 3712
rect 407040 3670 407068 118866
rect 408512 8022 408540 122046
rect 408500 8016 408552 8022
rect 408500 7958 408552 7964
rect 407302 6760 407358 6769
rect 407302 6695 407358 6704
rect 406108 3664 406160 3670
rect 406108 3606 406160 3612
rect 407028 3664 407080 3670
rect 407028 3606 407080 3612
rect 406120 480 406148 3606
rect 407316 480 407344 6695
rect 409696 6452 409748 6458
rect 409696 6394 409748 6400
rect 410892 6452 410944 6458
rect 410892 6394 410944 6400
rect 408500 4684 408552 4690
rect 408500 4626 408552 4632
rect 408512 480 408540 4626
rect 409708 480 409736 6394
rect 410904 480 410932 6394
rect 411180 3126 411208 122060
rect 413572 118318 413600 122060
rect 413940 121990 413968 122159
rect 415780 121990 415808 122182
rect 424966 122159 425022 122168
rect 426438 122224 426494 122233
rect 426438 122159 426494 122168
rect 413928 121984 413980 121990
rect 413928 121926 413980 121932
rect 415768 121984 415820 121990
rect 415768 121926 415820 121932
rect 413560 118312 413612 118318
rect 413560 118254 413612 118260
rect 413928 118312 413980 118318
rect 413928 118254 413980 118260
rect 411260 111240 411312 111246
rect 411258 111208 411260 111217
rect 411312 111208 411314 111217
rect 411258 111143 411314 111152
rect 412546 19136 412602 19145
rect 412546 19071 412602 19080
rect 412560 18873 412588 19071
rect 412546 18864 412602 18873
rect 412546 18799 412602 18808
rect 412640 14476 412692 14482
rect 412640 14418 412692 14424
rect 412088 3664 412140 3670
rect 412088 3606 412140 3612
rect 411168 3120 411220 3126
rect 411168 3062 411220 3068
rect 412100 480 412128 3606
rect 412652 610 412680 14418
rect 413940 9246 413968 118254
rect 415964 116142 415992 122060
rect 418172 122046 418370 122074
rect 419644 122046 420762 122074
rect 416780 119196 416832 119202
rect 416780 119138 416832 119144
rect 415492 116136 415544 116142
rect 415492 116078 415544 116084
rect 415952 116136 416004 116142
rect 415952 116078 416004 116084
rect 413928 9240 413980 9246
rect 413928 9182 413980 9188
rect 414478 6488 414534 6497
rect 414478 6423 414534 6432
rect 413836 4208 413888 4214
rect 413836 4150 413888 4156
rect 414020 4208 414072 4214
rect 414020 4150 414072 4156
rect 413848 3890 413876 4150
rect 414032 3890 414060 4150
rect 413848 3862 414060 3890
rect 412640 604 412692 610
rect 412640 546 412692 552
rect 413284 604 413336 610
rect 413284 546 413336 552
rect 413296 480 413324 546
rect 414492 480 414520 6423
rect 415504 3670 415532 116078
rect 415676 5364 415728 5370
rect 415676 5306 415728 5312
rect 415492 3664 415544 3670
rect 415492 3606 415544 3612
rect 415688 480 415716 5306
rect 416792 626 416820 119138
rect 417976 6384 418028 6390
rect 417976 6326 418028 6332
rect 416792 598 416912 626
rect 416884 480 416912 598
rect 417988 480 418016 6326
rect 418172 5506 418200 122046
rect 419446 121680 419502 121689
rect 419446 121615 419502 121624
rect 418160 5500 418212 5506
rect 418160 5442 418212 5448
rect 419460 626 419488 121615
rect 419540 118788 419592 118794
rect 419540 118730 419592 118736
rect 419552 7682 419580 118730
rect 419540 7676 419592 7682
rect 419540 7618 419592 7624
rect 419644 4622 419672 122046
rect 423140 118930 423168 122060
rect 424980 121990 425008 122159
rect 424968 121984 425020 121990
rect 424968 121926 425020 121932
rect 425532 119474 425560 122060
rect 425520 119468 425572 119474
rect 425520 119410 425572 119416
rect 423128 118924 423180 118930
rect 423128 118866 423180 118872
rect 422208 118312 422260 118318
rect 422208 118254 422260 118260
rect 420736 111240 420788 111246
rect 420734 111208 420736 111217
rect 420788 111208 420790 111217
rect 420734 111143 420790 111152
rect 420368 7676 420420 7682
rect 420368 7618 420420 7624
rect 419632 4616 419684 4622
rect 419632 4558 419684 4564
rect 419184 598 419488 626
rect 419184 480 419212 598
rect 420380 480 420408 7618
rect 422220 3126 422248 118254
rect 425610 35184 425666 35193
rect 425610 35119 425666 35128
rect 425624 29034 425652 35119
rect 425612 29028 425664 29034
rect 425612 28970 425664 28976
rect 422298 19136 422354 19145
rect 422298 19071 422354 19080
rect 422312 18873 422340 19071
rect 422298 18864 422354 18873
rect 422298 18799 422354 18808
rect 426452 12442 426480 122159
rect 427924 121242 427952 122060
rect 427912 121236 427964 121242
rect 427912 121178 427964 121184
rect 430316 119950 430344 122060
rect 432722 122046 433288 122074
rect 431868 121236 431920 121242
rect 431868 121178 431920 121184
rect 430304 119944 430356 119950
rect 430304 119886 430356 119892
rect 430578 111208 430634 111217
rect 430578 111143 430580 111152
rect 430632 111143 430634 111152
rect 430580 111114 430632 111120
rect 427820 29028 427872 29034
rect 427820 28970 427872 28976
rect 427832 19310 427860 28970
rect 427636 19304 427688 19310
rect 427636 19246 427688 19252
rect 427820 19304 427872 19310
rect 427820 19246 427872 19252
rect 426440 12436 426492 12442
rect 426440 12378 426492 12384
rect 427544 12436 427596 12442
rect 427544 12378 427596 12384
rect 422758 6488 422814 6497
rect 422758 6423 422814 6432
rect 421564 3120 421616 3126
rect 421564 3062 421616 3068
rect 422208 3120 422260 3126
rect 422208 3062 422260 3068
rect 421576 480 421604 3062
rect 422772 480 422800 6423
rect 423956 6384 424008 6390
rect 423956 6326 424008 6332
rect 423968 480 423996 6326
rect 426348 4888 426400 4894
rect 426348 4830 426400 4836
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 424980 3754 425008 4150
rect 424980 3726 425100 3754
rect 425072 2961 425100 3726
rect 425150 3632 425206 3641
rect 425150 3567 425206 3576
rect 425058 2952 425114 2961
rect 425058 2887 425114 2896
rect 425164 480 425192 3567
rect 426360 480 426388 4830
rect 427556 480 427584 12378
rect 427648 9761 427676 19246
rect 429936 12096 429988 12102
rect 429936 12038 429988 12044
rect 427634 9752 427690 9761
rect 427634 9687 427690 9696
rect 427818 9752 427874 9761
rect 427818 9687 427874 9696
rect 427832 9654 427860 9687
rect 427820 9648 427872 9654
rect 427820 9590 427872 9596
rect 428740 604 428792 610
rect 428740 546 428792 552
rect 428752 480 428780 546
rect 429948 480 429976 12038
rect 431880 3670 431908 121178
rect 432050 19136 432106 19145
rect 432050 19071 432106 19080
rect 432064 18873 432092 19071
rect 432050 18864 432106 18873
rect 432050 18799 432106 18808
rect 432328 6112 432380 6118
rect 432328 6054 432380 6060
rect 431132 3664 431184 3670
rect 431132 3606 431184 3612
rect 431868 3664 431920 3670
rect 431868 3606 431920 3612
rect 431144 480 431172 3606
rect 432340 480 432368 6054
rect 433260 4894 433288 122046
rect 435100 118862 435128 122060
rect 437492 119950 437520 122060
rect 438872 122046 439898 122074
rect 442290 122046 442948 122074
rect 437480 119944 437532 119950
rect 437480 119886 437532 119892
rect 438768 119944 438820 119950
rect 438768 119886 438820 119892
rect 433340 118856 433392 118862
rect 433340 118798 433392 118804
rect 435088 118856 435140 118862
rect 435088 118798 435140 118804
rect 436008 118856 436060 118862
rect 436008 118798 436060 118804
rect 433352 7682 433380 118798
rect 435822 77208 435878 77217
rect 435822 77143 435878 77152
rect 435836 67697 435864 77143
rect 435822 67688 435878 67697
rect 435822 67623 435878 67632
rect 433522 10432 433578 10441
rect 433522 10367 433578 10376
rect 433340 7676 433392 7682
rect 433340 7618 433392 7624
rect 433248 4888 433300 4894
rect 433248 4830 433300 4836
rect 433536 480 433564 10367
rect 436020 9178 436048 118798
rect 436100 96756 436152 96762
rect 436100 96698 436152 96704
rect 436112 96626 436140 96698
rect 436100 96620 436152 96626
rect 436100 96562 436152 96568
rect 436284 96620 436336 96626
rect 436284 96562 436336 96568
rect 436296 87009 436324 96562
rect 436098 87000 436154 87009
rect 436098 86935 436100 86944
rect 436152 86935 436154 86944
rect 436282 87000 436338 87009
rect 436282 86935 436338 86944
rect 436100 86906 436152 86912
rect 436100 77308 436152 77314
rect 436100 77250 436152 77256
rect 436112 77217 436140 77250
rect 436098 77208 436154 77217
rect 436098 77143 436154 77152
rect 436098 67688 436154 67697
rect 436098 67623 436154 67632
rect 436112 67590 436140 67623
rect 436100 67584 436152 67590
rect 436100 67526 436152 67532
rect 436100 57996 436152 58002
rect 436100 57938 436152 57944
rect 436112 57866 436140 57938
rect 436100 57860 436152 57866
rect 436100 57802 436152 57808
rect 436100 48340 436152 48346
rect 436100 48282 436152 48288
rect 436112 38842 436140 48282
rect 436112 38814 436232 38842
rect 436204 38706 436232 38814
rect 436112 38678 436232 38706
rect 436112 38622 436140 38678
rect 436100 38616 436152 38622
rect 436100 38558 436152 38564
rect 436100 29096 436152 29102
rect 436100 29038 436152 29044
rect 436112 28966 436140 29038
rect 436100 28960 436152 28966
rect 436100 28902 436152 28908
rect 436192 28960 436244 28966
rect 436192 28902 436244 28908
rect 436204 19394 436232 28902
rect 436112 19366 436232 19394
rect 436112 19310 436140 19366
rect 436100 19304 436152 19310
rect 436100 19246 436152 19252
rect 437478 11792 437534 11801
rect 437478 11727 437534 11736
rect 436100 9784 436152 9790
rect 436100 9726 436152 9732
rect 436112 9654 436140 9726
rect 436100 9648 436152 9654
rect 436100 9590 436152 9596
rect 436008 9172 436060 9178
rect 436008 9114 436060 9120
rect 434628 7676 434680 7682
rect 434628 7618 434680 7624
rect 434640 480 434668 7618
rect 435822 3632 435878 3641
rect 435822 3567 435878 3576
rect 435836 480 435864 3567
rect 437492 610 437520 11727
rect 438780 10402 438808 119886
rect 438768 10396 438820 10402
rect 438768 10338 438820 10344
rect 438872 7818 438900 122046
rect 440148 121984 440200 121990
rect 440148 121926 440200 121932
rect 440160 111314 440188 121926
rect 441712 119332 441764 119338
rect 441712 119274 441764 119280
rect 440148 111308 440200 111314
rect 440148 111250 440200 111256
rect 440146 111208 440202 111217
rect 440068 111178 440146 111194
rect 440056 111172 440146 111178
rect 440108 111166 440146 111172
rect 440146 111143 440202 111152
rect 440056 111114 440108 111120
rect 440148 111104 440200 111110
rect 440148 111046 440200 111052
rect 438860 7812 438912 7818
rect 438860 7754 438912 7760
rect 440160 3670 440188 111046
rect 441618 19136 441674 19145
rect 441618 19071 441674 19080
rect 441632 18873 441660 19071
rect 441618 18864 441674 18873
rect 441618 18799 441674 18808
rect 439412 3664 439464 3670
rect 439412 3606 439464 3612
rect 440148 3664 440200 3670
rect 440148 3606 440200 3612
rect 437020 604 437072 610
rect 437020 546 437072 552
rect 437480 604 437532 610
rect 437480 546 437532 552
rect 438216 604 438268 610
rect 438216 546 438268 552
rect 437032 480 437060 546
rect 438228 480 438256 546
rect 439424 480 439452 3606
rect 440608 3120 440660 3126
rect 440608 3062 440660 3068
rect 440620 480 440648 3062
rect 441724 626 441752 119274
rect 442920 5506 442948 122046
rect 444392 122046 444682 122074
rect 442908 5500 442960 5506
rect 442908 5442 442960 5448
rect 444392 4758 444420 122046
rect 445852 121508 445904 121514
rect 445852 121450 445904 121456
rect 445864 115938 445892 121450
rect 447060 119066 447088 122060
rect 449268 119270 449296 122060
rect 449256 119264 449308 119270
rect 449256 119206 449308 119212
rect 451660 119134 451688 122060
rect 454052 121378 454080 122060
rect 455432 122046 456458 122074
rect 458850 122046 459508 122074
rect 454040 121372 454092 121378
rect 454040 121314 454092 121320
rect 451648 119128 451700 119134
rect 451648 119070 451700 119076
rect 447048 119060 447100 119066
rect 447048 119002 447100 119008
rect 451280 116612 451332 116618
rect 451280 116554 451332 116560
rect 445852 115932 445904 115938
rect 445852 115874 445904 115880
rect 444470 111208 444526 111217
rect 444470 111143 444526 111152
rect 444484 110945 444512 111143
rect 444470 110936 444526 110945
rect 444470 110871 444526 110880
rect 445852 106344 445904 106350
rect 445852 106286 445904 106292
rect 445864 96626 445892 106286
rect 445852 96620 445904 96626
rect 445852 96562 445904 96568
rect 445852 87032 445904 87038
rect 445852 86974 445904 86980
rect 444472 83496 444524 83502
rect 444472 83438 444524 83444
rect 444380 4752 444432 4758
rect 444380 4694 444432 4700
rect 442262 3768 442318 3777
rect 442262 3703 442318 3712
rect 442276 2961 442304 3703
rect 444196 3664 444248 3670
rect 444196 3606 444248 3612
rect 442998 3088 443054 3097
rect 442998 3023 443054 3032
rect 442262 2952 442318 2961
rect 442262 2887 442318 2896
rect 441724 598 441844 626
rect 441816 480 441844 598
rect 443012 480 443040 3023
rect 444208 480 444236 3606
rect 444484 610 444512 83438
rect 445864 77178 445892 86974
rect 445852 77172 445904 77178
rect 445852 77114 445904 77120
rect 445852 67652 445904 67658
rect 445852 67594 445904 67600
rect 445864 57934 445892 67594
rect 445852 57928 445904 57934
rect 445852 57870 445904 57876
rect 445852 48340 445904 48346
rect 445852 48282 445904 48288
rect 445864 38622 445892 48282
rect 445852 38616 445904 38622
rect 445852 38558 445904 38564
rect 445852 29028 445904 29034
rect 445852 28970 445904 28976
rect 445864 19310 445892 28970
rect 445852 19304 445904 19310
rect 445852 19246 445904 19252
rect 447138 19136 447194 19145
rect 447138 19071 447194 19080
rect 447152 18873 447180 19071
rect 447138 18864 447194 18873
rect 447138 18799 447194 18808
rect 448518 18728 448574 18737
rect 448518 18663 448574 18672
rect 445760 10940 445812 10946
rect 445760 10882 445812 10888
rect 445772 5438 445800 10882
rect 445852 9716 445904 9722
rect 445852 9658 445904 9664
rect 445760 5432 445812 5438
rect 445760 5374 445812 5380
rect 445864 3210 445892 9658
rect 445772 3182 445892 3210
rect 445772 610 445800 3182
rect 447784 3120 447836 3126
rect 447784 3062 447836 3068
rect 444472 604 444524 610
rect 444472 546 444524 552
rect 445392 604 445444 610
rect 445392 546 445444 552
rect 445760 604 445812 610
rect 445760 546 445812 552
rect 446588 604 446640 610
rect 446588 546 446640 552
rect 445404 480 445432 546
rect 446600 480 446628 546
rect 447796 480 447824 3062
rect 448532 610 448560 18663
rect 450176 3052 450228 3058
rect 450176 2994 450228 3000
rect 448520 604 448572 610
rect 448520 546 448572 552
rect 448980 604 449032 610
rect 448980 546 449032 552
rect 448992 480 449020 546
rect 450188 480 450216 2994
rect 451292 2990 451320 116554
rect 454040 113824 454092 113830
rect 454040 113766 454092 113772
rect 453946 39264 454002 39273
rect 453946 39199 454002 39208
rect 452660 17196 452712 17202
rect 452660 17138 452712 17144
rect 452672 10946 452700 17138
rect 452660 10940 452712 10946
rect 452660 10882 452712 10888
rect 451372 6044 451424 6050
rect 451372 5986 451424 5992
rect 451280 2984 451332 2990
rect 451280 2926 451332 2932
rect 451384 2802 451412 5986
rect 451462 3768 451518 3777
rect 451462 3703 451518 3712
rect 451476 2825 451504 3703
rect 452476 2984 452528 2990
rect 452476 2926 452528 2932
rect 451292 2774 451412 2802
rect 451462 2816 451518 2825
rect 451292 480 451320 2774
rect 451462 2751 451518 2760
rect 452488 480 452516 2926
rect 453960 610 453988 39199
rect 454052 610 454080 113766
rect 454684 27600 454736 27606
rect 454684 27542 454736 27548
rect 454696 17202 454724 27542
rect 454684 17196 454736 17202
rect 454684 17138 454736 17144
rect 455432 4690 455460 122046
rect 456708 121372 456760 121378
rect 456708 121314 456760 121320
rect 455420 4684 455472 4690
rect 455420 4626 455472 4632
rect 456720 2990 456748 121314
rect 458178 115152 458234 115161
rect 458178 115087 458234 115096
rect 457444 36372 457496 36378
rect 457444 36314 457496 36320
rect 457456 27606 457484 36314
rect 457444 27600 457496 27606
rect 457444 27542 457496 27548
rect 457260 8084 457312 8090
rect 457260 8026 457312 8032
rect 456064 2984 456116 2990
rect 456064 2926 456116 2932
rect 456708 2984 456760 2990
rect 456708 2926 456760 2932
rect 453672 604 453724 610
rect 453672 546 453724 552
rect 453948 604 454000 610
rect 453948 546 454000 552
rect 454040 604 454092 610
rect 454040 546 454092 552
rect 454868 604 454920 610
rect 454868 546 454920 552
rect 453684 480 453712 546
rect 454880 480 454908 546
rect 456076 480 456104 2926
rect 457272 480 457300 8026
rect 458192 626 458220 115087
rect 458272 12436 458324 12442
rect 458272 12378 458324 12384
rect 458284 5234 458312 12378
rect 459480 7682 459508 122046
rect 461228 119950 461256 122060
rect 461216 119944 461268 119950
rect 461216 119886 461268 119892
rect 463620 119474 463648 122060
rect 466012 121310 466040 122060
rect 467852 122046 468418 122074
rect 470612 122046 470810 122074
rect 466000 121304 466052 121310
rect 466000 121246 466052 121252
rect 463608 119468 463660 119474
rect 463608 119410 463660 119416
rect 467748 119332 467800 119338
rect 467748 119274 467800 119280
rect 459650 111208 459706 111217
rect 459650 111143 459706 111152
rect 459664 110673 459692 111143
rect 459650 110664 459706 110673
rect 459650 110599 459706 110608
rect 467104 68944 467156 68950
rect 467104 68886 467156 68892
rect 467116 57662 467144 68886
rect 465724 57656 465776 57662
rect 465724 57598 465776 57604
rect 467104 57656 467156 57662
rect 467104 57598 467156 57604
rect 465736 39370 465764 57598
rect 467104 53712 467156 53718
rect 467104 53654 467156 53660
rect 459560 39364 459612 39370
rect 459560 39306 459612 39312
rect 465724 39364 465776 39370
rect 465724 39306 465776 39312
rect 459572 36378 459600 39306
rect 459560 36372 459612 36378
rect 459560 36314 459612 36320
rect 467116 19242 467144 53654
rect 463700 19236 463752 19242
rect 463700 19178 463752 19184
rect 467104 19236 467156 19242
rect 467104 19178 467156 19184
rect 462594 18864 462650 18873
rect 462594 18799 462650 18808
rect 462608 18465 462636 18799
rect 462594 18456 462650 18465
rect 462594 18391 462650 18400
rect 463712 15230 463740 19178
rect 461860 15224 461912 15230
rect 461860 15166 461912 15172
rect 463700 15224 463752 15230
rect 463700 15166 463752 15172
rect 461872 12510 461900 15166
rect 461860 12504 461912 12510
rect 461860 12446 461912 12452
rect 462044 12028 462096 12034
rect 462044 11970 462096 11976
rect 459468 7676 459520 7682
rect 459468 7618 459520 7624
rect 458272 5228 458324 5234
rect 458272 5170 458324 5176
rect 460846 3360 460902 3369
rect 460846 3295 460902 3304
rect 459650 2952 459706 2961
rect 459650 2887 459706 2896
rect 458192 598 458496 626
rect 458468 480 458496 598
rect 459664 480 459692 2887
rect 460860 480 460888 3295
rect 462056 480 462084 11970
rect 465630 6896 465686 6905
rect 465630 6831 465686 6840
rect 463238 3768 463294 3777
rect 463238 3703 463294 3712
rect 463698 3768 463754 3777
rect 463698 3703 463754 3712
rect 463252 480 463280 3703
rect 463712 2825 463740 3703
rect 464434 3360 464490 3369
rect 464434 3295 464490 3304
rect 463698 2816 463754 2825
rect 463698 2751 463754 2760
rect 464448 480 464476 3295
rect 465644 480 465672 6831
rect 467760 2990 467788 119274
rect 467852 10538 467880 122046
rect 469128 121916 469180 121922
rect 469128 121858 469180 121864
rect 467840 10532 467892 10538
rect 467840 10474 467892 10480
rect 467932 5500 467984 5506
rect 467932 5442 467984 5448
rect 466828 2984 466880 2990
rect 466828 2926 466880 2932
rect 467748 2984 467800 2990
rect 467748 2926 467800 2932
rect 466840 480 466868 2926
rect 467944 480 467972 5442
rect 469140 480 469168 121858
rect 469218 111480 469274 111489
rect 469218 111415 469274 111424
rect 469232 111217 469260 111415
rect 469218 111208 469274 111217
rect 469218 111143 469274 111152
rect 470612 13326 470640 122046
rect 473188 119610 473216 122060
rect 474752 122046 475594 122074
rect 477512 122046 477986 122074
rect 473176 119604 473228 119610
rect 473176 119546 473228 119552
rect 471244 119468 471296 119474
rect 471244 119410 471296 119416
rect 470692 77172 470744 77178
rect 470692 77114 470744 77120
rect 470704 69086 470732 77114
rect 470692 69080 470744 69086
rect 470692 69022 470744 69028
rect 470600 13320 470652 13326
rect 470600 13262 470652 13268
rect 469312 7200 469364 7206
rect 469312 7142 469364 7148
rect 469220 5568 469272 5574
rect 469220 5510 469272 5516
rect 469232 5098 469260 5510
rect 469220 5092 469272 5098
rect 469220 5034 469272 5040
rect 469324 5030 469352 7142
rect 470322 6080 470378 6089
rect 470322 6015 470378 6024
rect 469312 5024 469364 5030
rect 469312 4966 469364 4972
rect 470336 480 470364 6015
rect 471256 5794 471284 119410
rect 473360 119400 473412 119406
rect 473360 119342 473412 119348
rect 472348 81456 472400 81462
rect 472348 81398 472400 81404
rect 472360 77178 472388 81398
rect 472348 77172 472400 77178
rect 472348 77114 472400 77120
rect 471980 57928 472032 57934
rect 471980 57870 472032 57876
rect 471992 53854 472020 57870
rect 471980 53848 472032 53854
rect 471980 53790 472032 53796
rect 471336 16652 471388 16658
rect 471336 16594 471388 16600
rect 471164 5766 471284 5794
rect 470598 3768 470654 3777
rect 470598 3703 470654 3712
rect 470612 2825 470640 3703
rect 471164 2922 471192 5766
rect 471244 5704 471296 5710
rect 471244 5646 471296 5652
rect 471256 4962 471284 5646
rect 471348 5574 471376 16594
rect 471612 11008 471664 11014
rect 471612 10950 471664 10956
rect 471624 7206 471652 10950
rect 471612 7200 471664 7206
rect 471612 7142 471664 7148
rect 472716 6316 472768 6322
rect 472716 6258 472768 6264
rect 471336 5568 471388 5574
rect 471336 5510 471388 5516
rect 471244 4956 471296 4962
rect 471244 4898 471296 4904
rect 471520 2984 471572 2990
rect 471520 2926 471572 2932
rect 471152 2916 471204 2922
rect 471152 2858 471204 2864
rect 470598 2816 470654 2825
rect 470598 2751 470654 2760
rect 471532 480 471560 2926
rect 472728 480 472756 6258
rect 473372 610 473400 119342
rect 474004 91112 474056 91118
rect 474004 91054 474056 91060
rect 474016 81462 474044 91054
rect 474004 81456 474056 81462
rect 474004 81398 474056 81404
rect 474752 14754 474780 122046
rect 476764 119468 476816 119474
rect 476764 119410 476816 119416
rect 475384 98456 475436 98462
rect 475384 98398 475436 98404
rect 475396 91118 475424 98398
rect 475384 91112 475436 91118
rect 475384 91054 475436 91060
rect 476028 62076 476080 62082
rect 476028 62018 476080 62024
rect 476040 58002 476068 62018
rect 476028 57996 476080 58002
rect 476028 57938 476080 57944
rect 474832 19304 474884 19310
rect 474832 19246 474884 19252
rect 474844 16658 474872 19246
rect 475016 18352 475068 18358
rect 475016 18294 475068 18300
rect 474832 16652 474884 16658
rect 474832 16594 474884 16600
rect 474740 14748 474792 14754
rect 474740 14690 474792 14696
rect 475028 11082 475056 18294
rect 475016 11076 475068 11082
rect 475016 11018 475068 11024
rect 476304 5296 476356 5302
rect 476304 5238 476356 5244
rect 475108 4888 475160 4894
rect 475108 4830 475160 4836
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 473924 480 473952 546
rect 475120 480 475148 4830
rect 476316 480 476344 5238
rect 476776 3194 476804 119410
rect 476856 38616 476908 38622
rect 476856 38558 476908 38564
rect 476868 18358 476896 38558
rect 476856 18352 476908 18358
rect 476856 18294 476908 18300
rect 477512 11898 477540 122046
rect 480168 121780 480220 121786
rect 480168 121722 480220 121728
rect 479524 119604 479576 119610
rect 479524 119546 479576 119552
rect 478786 111208 478842 111217
rect 478970 111208 479026 111217
rect 478842 111166 478970 111194
rect 478786 111143 478842 111152
rect 478970 111143 479026 111152
rect 478880 64864 478932 64870
rect 478880 64806 478932 64812
rect 478892 62150 478920 64806
rect 478880 62144 478932 62150
rect 478880 62086 478932 62092
rect 478880 24880 478932 24886
rect 478880 24822 478932 24828
rect 478892 19446 478920 24822
rect 478880 19440 478932 19446
rect 478880 19382 478932 19388
rect 478142 19136 478198 19145
rect 478142 19071 478198 19080
rect 478156 18465 478184 19071
rect 478142 18456 478198 18465
rect 478142 18391 478198 18400
rect 477500 11892 477552 11898
rect 477500 11834 477552 11840
rect 478052 7404 478104 7410
rect 478052 7346 478104 7352
rect 478064 5710 478092 7346
rect 478052 5704 478104 5710
rect 478052 5646 478104 5652
rect 478694 3768 478750 3777
rect 478694 3703 478750 3712
rect 476764 3188 476816 3194
rect 476764 3130 476816 3136
rect 477500 3188 477552 3194
rect 477500 3130 477552 3136
rect 477512 480 477540 3130
rect 478708 480 478736 3703
rect 479536 3262 479564 119546
rect 479616 107500 479668 107506
rect 479616 107442 479668 107448
rect 479628 98462 479656 107442
rect 479616 98456 479668 98462
rect 479616 98398 479668 98404
rect 479616 46980 479668 46986
rect 479616 46922 479668 46928
rect 479628 38622 479656 46922
rect 479616 38616 479668 38622
rect 479616 38558 479668 38564
rect 479524 3256 479576 3262
rect 479524 3198 479576 3204
rect 480180 626 480208 121722
rect 480364 119338 480392 122060
rect 481652 122046 482770 122074
rect 484412 122046 485162 122074
rect 480352 119332 480404 119338
rect 480352 119274 480404 119280
rect 481364 109812 481416 109818
rect 481364 109754 481416 109760
rect 481376 107506 481404 109754
rect 481364 107500 481416 107506
rect 481364 107442 481416 107448
rect 481272 53848 481324 53854
rect 481272 53790 481324 53796
rect 481284 46986 481312 53790
rect 481272 46980 481324 46986
rect 481272 46922 481324 46928
rect 480260 28960 480312 28966
rect 480260 28902 480312 28908
rect 480272 24886 480300 28902
rect 480260 24880 480312 24886
rect 480260 24822 480312 24828
rect 481652 5166 481680 122046
rect 484308 121848 484360 121854
rect 484308 121790 484360 121796
rect 481732 111852 481784 111858
rect 481732 111794 481784 111800
rect 481744 109818 481772 111794
rect 481732 109812 481784 109818
rect 481732 109754 481784 109760
rect 482560 71800 482612 71806
rect 482560 71742 482612 71748
rect 482572 64938 482600 71742
rect 482560 64932 482612 64938
rect 482560 64874 482612 64880
rect 482284 62144 482336 62150
rect 482284 62086 482336 62092
rect 482296 53854 482324 62086
rect 482284 53848 482336 53854
rect 482284 53790 482336 53796
rect 484216 36916 484268 36922
rect 484216 36858 484268 36864
rect 484228 29034 484256 36858
rect 484216 29028 484268 29034
rect 484216 28970 484268 28976
rect 481730 17232 481786 17241
rect 481730 17167 481786 17176
rect 481640 5160 481692 5166
rect 481640 5102 481692 5108
rect 481088 2848 481140 2854
rect 481088 2790 481140 2796
rect 479904 598 480208 626
rect 479904 480 479932 598
rect 481100 480 481128 2790
rect 481744 2666 481772 17167
rect 482836 12504 482888 12510
rect 482836 12446 482888 12452
rect 482848 7410 482876 12446
rect 482836 7404 482888 7410
rect 482836 7346 482888 7352
rect 482374 3768 482430 3777
rect 482374 3703 482430 3712
rect 482388 2825 482416 3703
rect 484320 3262 484348 121790
rect 484412 7614 484440 122046
rect 487068 119332 487120 119338
rect 487068 119274 487120 119280
rect 486148 81456 486200 81462
rect 486148 81398 486200 81404
rect 486160 79218 486188 81398
rect 485044 79212 485096 79218
rect 485044 79154 485096 79160
rect 486148 79212 486200 79218
rect 486148 79154 486200 79160
rect 485056 71806 485084 79154
rect 485044 71800 485096 71806
rect 485044 71742 485096 71748
rect 486148 40180 486200 40186
rect 486148 40122 486200 40128
rect 486160 36922 486188 40122
rect 486148 36916 486200 36922
rect 486148 36858 486200 36864
rect 485686 19136 485742 19145
rect 485686 19071 485742 19080
rect 485700 18737 485728 19071
rect 485686 18728 485742 18737
rect 485686 18663 485742 18672
rect 484400 7608 484452 7614
rect 484400 7550 484452 7556
rect 487080 3262 487108 119274
rect 487540 119270 487568 122060
rect 488448 121304 488500 121310
rect 488448 121246 488500 121252
rect 487528 119264 487580 119270
rect 487528 119206 487580 119212
rect 487528 114164 487580 114170
rect 487528 114106 487580 114112
rect 487540 111858 487568 114106
rect 487528 111852 487580 111858
rect 487528 111794 487580 111800
rect 487160 86760 487212 86766
rect 487160 86702 487212 86708
rect 487172 81462 487200 86702
rect 487160 81456 487212 81462
rect 487160 81398 487212 81404
rect 487160 64932 487212 64938
rect 487160 64874 487212 64880
rect 487172 62150 487200 64874
rect 487160 62144 487212 62150
rect 487160 62086 487212 62092
rect 487896 47388 487948 47394
rect 487896 47330 487948 47336
rect 487908 40186 487936 47330
rect 487896 40180 487948 40186
rect 487896 40122 487948 40128
rect 487804 40044 487856 40050
rect 487804 39986 487856 39992
rect 487816 12510 487844 39986
rect 487804 12504 487856 12510
rect 487804 12446 487856 12452
rect 483480 3256 483532 3262
rect 483480 3198 483532 3204
rect 484308 3256 484360 3262
rect 484308 3198 484360 3204
rect 485780 3256 485832 3262
rect 485780 3198 485832 3204
rect 487068 3256 487120 3262
rect 487068 3198 487120 3204
rect 482374 2816 482430 2825
rect 482374 2751 482430 2760
rect 481744 2638 482324 2666
rect 482296 480 482324 2638
rect 483492 480 483520 3198
rect 484584 2916 484636 2922
rect 484584 2858 484636 2864
rect 484596 480 484624 2858
rect 485792 480 485820 3198
rect 486974 2816 487030 2825
rect 486974 2751 487030 2760
rect 486988 480 487016 2751
rect 488460 626 488488 121246
rect 489932 119678 489960 122060
rect 492324 121718 492352 122060
rect 491300 121712 491352 121718
rect 491300 121654 491352 121660
rect 492312 121712 492364 121718
rect 492312 121654 492364 121660
rect 493324 121712 493376 121718
rect 493324 121654 493376 121660
rect 489920 119672 489972 119678
rect 489920 119614 489972 119620
rect 491208 119672 491260 119678
rect 491208 119614 491260 119620
rect 490564 117156 490616 117162
rect 490564 117098 490616 117104
rect 488538 111344 488594 111353
rect 488538 111279 488594 111288
rect 488552 111217 488580 111279
rect 488538 111208 488594 111217
rect 488538 111143 488594 111152
rect 490576 103154 490604 117098
rect 489184 103148 489236 103154
rect 489184 103090 489236 103096
rect 490564 103148 490616 103154
rect 490564 103090 490616 103096
rect 489196 86766 489224 103090
rect 489184 86760 489236 86766
rect 489184 86702 489236 86708
rect 491024 69012 491076 69018
rect 491024 68954 491076 68960
rect 491036 64938 491064 68954
rect 491024 64932 491076 64938
rect 491024 64874 491076 64880
rect 490288 53916 490340 53922
rect 490288 53858 490340 53864
rect 490300 53786 490328 53858
rect 488540 53780 488592 53786
rect 488540 53722 488592 53728
rect 490288 53780 490340 53786
rect 490288 53722 490340 53728
rect 488552 47394 488580 53722
rect 488540 47388 488592 47394
rect 488540 47330 488592 47336
rect 488540 47048 488592 47054
rect 488540 46990 488592 46996
rect 488552 40050 488580 46990
rect 488540 40044 488592 40050
rect 488540 39986 488592 39992
rect 491220 10470 491248 119614
rect 491208 10464 491260 10470
rect 491208 10406 491260 10412
rect 491312 5370 491340 121654
rect 492680 119400 492732 119406
rect 492680 119342 492732 119348
rect 492312 117360 492364 117366
rect 492312 117302 492364 117308
rect 492324 114170 492352 117302
rect 492312 114164 492364 114170
rect 492312 114106 492364 114112
rect 491944 62144 491996 62150
rect 491944 62086 491996 62092
rect 491956 53922 491984 62086
rect 491944 53916 491996 53922
rect 491944 53858 491996 53864
rect 491484 49836 491536 49842
rect 491484 49778 491536 49784
rect 491496 47054 491524 49778
rect 491484 47048 491536 47054
rect 491484 46990 491536 46996
rect 491392 10328 491444 10334
rect 491392 10270 491444 10276
rect 491300 5364 491352 5370
rect 491300 5306 491352 5312
rect 489368 2916 489420 2922
rect 489368 2858 489420 2864
rect 488184 598 488488 626
rect 488184 480 488212 598
rect 489380 480 489408 2858
rect 490562 2816 490618 2825
rect 490562 2751 490618 2760
rect 490576 480 490604 2751
rect 491404 2258 491432 10270
rect 491404 2230 491708 2258
rect 491680 626 491708 2230
rect 491680 598 491800 626
rect 492692 610 492720 119342
rect 492772 73228 492824 73234
rect 492772 73170 492824 73176
rect 492784 69086 492812 73170
rect 492772 69080 492824 69086
rect 492772 69022 492824 69028
rect 493336 3330 493364 121654
rect 494532 121446 494560 122060
rect 496084 121508 496136 121514
rect 496084 121450 496136 121456
rect 494520 121440 494572 121446
rect 494520 121382 494572 121388
rect 496096 121145 496124 121450
rect 496082 121136 496138 121145
rect 496082 121071 496138 121080
rect 496924 120086 496952 122060
rect 499316 121718 499344 122060
rect 498476 121712 498528 121718
rect 498212 121660 498476 121666
rect 498212 121654 498528 121660
rect 499304 121712 499356 121718
rect 499304 121654 499356 121660
rect 498212 121638 498516 121654
rect 496912 120080 496964 120086
rect 496912 120022 496964 120028
rect 495440 119808 495492 119814
rect 495440 119750 495492 119756
rect 493506 117192 493562 117201
rect 493506 117127 493508 117136
rect 493560 117127 493562 117136
rect 493508 117098 493560 117104
rect 494060 76628 494112 76634
rect 494060 76570 494112 76576
rect 494072 73234 494100 76570
rect 494704 74520 494756 74526
rect 494704 74462 494756 74468
rect 494060 73228 494112 73234
rect 494060 73170 494112 73176
rect 494244 66972 494296 66978
rect 494244 66914 494296 66920
rect 494256 62150 494284 66914
rect 494244 62144 494296 62150
rect 494244 62086 494296 62092
rect 494716 57526 494744 74462
rect 493600 57520 493652 57526
rect 493600 57462 493652 57468
rect 494704 57520 494756 57526
rect 494704 57462 494756 57468
rect 493612 49842 493640 57462
rect 493600 49836 493652 49842
rect 493600 49778 493652 49784
rect 495348 11824 495400 11830
rect 495348 11766 495400 11772
rect 494704 4276 494756 4282
rect 494704 4218 494756 4224
rect 494716 4049 494744 4218
rect 495072 4208 495124 4214
rect 495072 4150 495124 4156
rect 494702 4040 494758 4049
rect 494702 3975 494758 3984
rect 495084 3777 495112 4150
rect 495070 3768 495126 3777
rect 495070 3703 495126 3712
rect 493324 3324 493376 3330
rect 493324 3266 493376 3272
rect 494152 3324 494204 3330
rect 494152 3266 494204 3272
rect 491772 480 491800 598
rect 492680 604 492732 610
rect 492680 546 492732 552
rect 492956 604 493008 610
rect 492956 546 493008 552
rect 492968 480 492996 546
rect 494164 480 494192 3266
rect 495360 480 495388 11766
rect 495452 610 495480 119750
rect 496726 118960 496782 118969
rect 496726 118895 496782 118904
rect 496740 117366 496768 118895
rect 496728 117360 496780 117366
rect 496728 117302 496780 117308
rect 497464 99884 497516 99890
rect 497464 99826 497516 99832
rect 497476 78742 497504 99826
rect 497556 84516 497608 84522
rect 497556 84458 497608 84464
rect 495992 78736 496044 78742
rect 495992 78678 496044 78684
rect 497464 78736 497516 78742
rect 497464 78678 497516 78684
rect 496004 76634 496032 78678
rect 495992 76628 496044 76634
rect 495992 76570 496044 76576
rect 497568 74594 497596 84458
rect 497556 74588 497608 74594
rect 497556 74530 497608 74536
rect 496728 73160 496780 73166
rect 496728 73102 496780 73108
rect 496740 66978 496768 73102
rect 496728 66972 496780 66978
rect 496728 66914 496780 66920
rect 498212 13462 498240 121638
rect 499396 121440 499448 121446
rect 499210 121408 499266 121417
rect 499394 121408 499396 121417
rect 499448 121408 499450 121417
rect 499266 121366 499344 121394
rect 499210 121343 499266 121352
rect 499316 121281 499344 121366
rect 499854 121408 499910 121417
rect 499394 121343 499450 121352
rect 499776 121366 499854 121394
rect 499776 121310 499804 121366
rect 499854 121343 499910 121352
rect 499764 121304 499816 121310
rect 499118 121272 499174 121281
rect 499118 121207 499174 121216
rect 499302 121272 499358 121281
rect 499764 121246 499816 121252
rect 499302 121207 499358 121216
rect 499948 121236 500000 121242
rect 498382 121000 498438 121009
rect 498382 120935 498438 120944
rect 498566 121000 498622 121009
rect 498566 120935 498622 120944
rect 498396 120601 498424 120935
rect 498382 120592 498438 120601
rect 498382 120527 498438 120536
rect 498580 116793 498608 120935
rect 498936 120692 498988 120698
rect 498936 120634 498988 120640
rect 498948 120601 498976 120634
rect 498934 120592 498990 120601
rect 498934 120527 498990 120536
rect 499132 120465 499160 121207
rect 499948 121178 500000 121184
rect 499960 120737 499988 121178
rect 500040 121100 500092 121106
rect 500040 121042 500092 121048
rect 499946 120728 500002 120737
rect 499946 120663 500002 120672
rect 499118 120456 499174 120465
rect 499118 120391 499174 120400
rect 500052 120329 500080 121042
rect 500038 120320 500094 120329
rect 500038 120255 500094 120264
rect 500224 118380 500276 118386
rect 500224 118322 500276 118328
rect 500132 117836 500184 117842
rect 500132 117778 500184 117784
rect 498566 116784 498622 116793
rect 498566 116719 498622 116728
rect 500144 113393 500172 117778
rect 500130 113384 500186 113393
rect 500130 113319 500186 113328
rect 500130 109712 500186 109721
rect 500130 109647 500186 109656
rect 500144 96801 500172 109647
rect 500130 96792 500186 96801
rect 500130 96727 500186 96736
rect 499946 95160 500002 95169
rect 499946 95095 500002 95104
rect 499960 73166 499988 95095
rect 500236 93906 500264 118322
rect 500328 118017 500356 122567
rect 500406 121000 500462 121009
rect 500406 120935 500462 120944
rect 500314 118008 500370 118017
rect 500314 117943 500370 117952
rect 500316 114708 500368 114714
rect 500316 114650 500368 114656
rect 500328 99890 500356 114650
rect 500420 114617 500448 120935
rect 501524 119338 501552 124578
rect 501616 123593 501644 126103
rect 501602 123584 501658 123593
rect 501602 123519 501658 123528
rect 501604 123480 501656 123486
rect 501602 123448 501604 123457
rect 501656 123448 501658 123457
rect 501602 123383 501658 123392
rect 501604 123344 501656 123350
rect 501604 123286 501656 123292
rect 501512 119332 501564 119338
rect 501512 119274 501564 119280
rect 500868 119196 500920 119202
rect 500868 119138 500920 119144
rect 500406 114608 500462 114617
rect 500406 114543 500462 114552
rect 500774 104680 500830 104689
rect 500774 104615 500830 104624
rect 500316 99884 500368 99890
rect 500316 99826 500368 99832
rect 500316 98048 500368 98054
rect 500316 97990 500368 97996
rect 500224 93900 500276 93906
rect 500224 93842 500276 93848
rect 500328 84522 500356 97990
rect 500590 92848 500646 92857
rect 500590 92783 500646 92792
rect 500604 91769 500632 92783
rect 500682 92712 500738 92721
rect 500682 92647 500738 92656
rect 500590 91760 500646 91769
rect 500590 91695 500646 91704
rect 500316 84516 500368 84522
rect 500316 84458 500368 84464
rect 500224 77308 500276 77314
rect 500224 77250 500276 77256
rect 499948 73160 500000 73166
rect 499948 73102 500000 73108
rect 500040 73160 500092 73166
rect 500040 73102 500092 73108
rect 499394 72992 499450 73001
rect 499394 72927 499450 72936
rect 498382 67552 498438 67561
rect 498382 67487 498438 67496
rect 498396 62801 498424 67487
rect 498382 62792 498438 62801
rect 498382 62727 498438 62736
rect 498382 57760 498438 57769
rect 498382 57695 498438 57704
rect 498396 48385 498424 57695
rect 499408 55457 499436 72927
rect 500052 56817 500080 73102
rect 500038 56808 500094 56817
rect 500038 56743 500094 56752
rect 499394 55448 499450 55457
rect 499394 55383 499450 55392
rect 500236 53802 500264 77250
rect 500406 77208 500462 77217
rect 500406 77143 500462 77152
rect 500420 68377 500448 77143
rect 500696 73166 500724 92647
rect 500788 87009 500816 104615
rect 500774 87000 500830 87009
rect 500774 86935 500830 86944
rect 500684 73160 500736 73166
rect 500684 73102 500736 73108
rect 500776 73160 500828 73166
rect 500776 73102 500828 73108
rect 500406 68368 500462 68377
rect 500406 68303 500462 68312
rect 500498 56536 500554 56545
rect 500498 56471 500554 56480
rect 500236 53774 500356 53802
rect 499946 49056 500002 49065
rect 499946 48991 500002 49000
rect 498382 48376 498438 48385
rect 498382 48311 498438 48320
rect 499960 38865 499988 48991
rect 500328 39114 500356 53774
rect 500406 49056 500462 49065
rect 500406 48991 500462 49000
rect 500420 39273 500448 48991
rect 500512 48929 500540 56471
rect 500498 48920 500554 48929
rect 500498 48855 500554 48864
rect 500788 44198 500816 73102
rect 500684 44192 500736 44198
rect 500684 44134 500736 44140
rect 500776 44192 500828 44198
rect 500776 44134 500828 44140
rect 500406 39264 500462 39273
rect 500406 39199 500462 39208
rect 500236 39086 500356 39114
rect 499946 38856 500002 38865
rect 499946 38791 500002 38800
rect 498290 34368 498346 34377
rect 498290 34303 498346 34312
rect 498304 25129 498332 34303
rect 498290 25120 498346 25129
rect 498290 25055 498346 25064
rect 498474 15328 498530 15337
rect 498474 15263 498530 15272
rect 498200 13456 498252 13462
rect 498200 13398 498252 13404
rect 498488 9761 498516 15263
rect 500236 15201 500264 39086
rect 500590 37224 500646 37233
rect 500590 37159 500646 37168
rect 500604 29753 500632 37159
rect 500590 29744 500646 29753
rect 500590 29679 500646 29688
rect 499946 15192 500002 15201
rect 499946 15127 500002 15136
rect 500222 15192 500278 15201
rect 500222 15127 500278 15136
rect 498474 9752 498530 9761
rect 498474 9687 498530 9696
rect 497740 6316 497792 6322
rect 497740 6258 497792 6264
rect 495624 4276 495676 4282
rect 495624 4218 495676 4224
rect 495532 4208 495584 4214
rect 495532 4150 495584 4156
rect 495544 3913 495572 4150
rect 495636 4049 495664 4218
rect 495622 4040 495678 4049
rect 495622 3975 495678 3984
rect 495530 3904 495586 3913
rect 495530 3839 495586 3848
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 6258
rect 499960 5574 499988 15127
rect 500696 7274 500724 44134
rect 500040 7268 500092 7274
rect 500040 7210 500092 7216
rect 500684 7268 500736 7274
rect 500684 7210 500736 7216
rect 499948 5568 500000 5574
rect 499948 5510 500000 5516
rect 498936 3868 498988 3874
rect 498936 3810 498988 3816
rect 498948 480 498976 3810
rect 500052 3641 500080 7210
rect 500132 5568 500184 5574
rect 500132 5510 500184 5516
rect 500144 4350 500172 5510
rect 500132 4344 500184 4350
rect 500132 4286 500184 4292
rect 500880 4146 500908 119138
rect 501236 102128 501288 102134
rect 501236 102070 501288 102076
rect 501248 98054 501276 102070
rect 501236 98048 501288 98054
rect 501236 97990 501288 97996
rect 501236 9240 501288 9246
rect 501236 9182 501288 9188
rect 500132 4140 500184 4146
rect 500132 4082 500184 4088
rect 500868 4140 500920 4146
rect 500868 4082 500920 4088
rect 500038 3632 500094 3641
rect 500038 3567 500094 3576
rect 500144 480 500172 4082
rect 501248 480 501276 9182
rect 501616 4146 501644 123286
rect 501604 4140 501656 4146
rect 501604 4082 501656 4088
rect 501708 3874 501736 133146
rect 501800 124642 501828 457127
rect 501892 158846 501920 580926
rect 501984 499526 502012 582762
rect 502064 582208 502116 582214
rect 502064 582150 502116 582156
rect 502076 581058 502104 582150
rect 502064 581052 502116 581058
rect 502064 580994 502116 581000
rect 502062 573744 502118 573753
rect 502062 573679 502118 573688
rect 502076 572257 502104 573679
rect 502062 572248 502118 572257
rect 502062 572183 502118 572192
rect 502062 557152 502118 557161
rect 502062 557087 502118 557096
rect 502076 547913 502104 557087
rect 502062 547904 502118 547913
rect 502062 547839 502118 547848
rect 502062 500576 502118 500585
rect 502062 500511 502118 500520
rect 501972 499520 502024 499526
rect 501972 499462 502024 499468
rect 502076 493377 502104 500511
rect 502062 493368 502118 493377
rect 502062 493303 502118 493312
rect 502154 464400 502210 464409
rect 502154 464335 502210 464344
rect 502168 454889 502196 464335
rect 502154 454880 502210 454889
rect 502154 454815 502210 454824
rect 502062 454744 502118 454753
rect 502062 454679 502118 454688
rect 502076 449041 502104 454679
rect 502062 449032 502118 449041
rect 502062 448967 502118 448976
rect 501970 442504 502026 442513
rect 501970 442439 502026 442448
rect 501984 439793 502012 442439
rect 501970 439784 502026 439793
rect 501970 439719 502026 439728
rect 502154 427816 502210 427825
rect 502154 427751 502210 427760
rect 502062 423464 502118 423473
rect 502062 423399 502118 423408
rect 502076 414089 502104 423399
rect 502168 418305 502196 427751
rect 502154 418296 502210 418305
rect 502154 418231 502210 418240
rect 502062 414080 502118 414089
rect 502062 414015 502118 414024
rect 502062 413808 502118 413817
rect 502062 413743 502118 413752
rect 501970 411496 502026 411505
rect 501970 411431 502026 411440
rect 501984 410145 502012 411431
rect 501970 410136 502026 410145
rect 501970 410071 502026 410080
rect 501970 405784 502026 405793
rect 501970 405719 502026 405728
rect 501984 400761 502012 405719
rect 502076 405657 502104 413743
rect 502062 405648 502118 405657
rect 502062 405583 502118 405592
rect 502062 403744 502118 403753
rect 502062 403679 502118 403688
rect 501970 400752 502026 400761
rect 501970 400687 502026 400696
rect 502076 398721 502104 403679
rect 502062 398712 502118 398721
rect 502062 398647 502118 398656
rect 502246 394632 502302 394641
rect 502246 394567 502302 394576
rect 502260 387161 502288 394567
rect 502246 387152 502302 387161
rect 502246 387087 502302 387096
rect 501970 351656 502026 351665
rect 501970 351591 502026 351600
rect 501984 346361 502012 351591
rect 502062 350568 502118 350577
rect 502062 350503 502118 350512
rect 502076 346497 502104 350503
rect 502062 346488 502118 346497
rect 502062 346423 502118 346432
rect 501970 346352 502026 346361
rect 501970 346287 502026 346296
rect 502154 344992 502210 345001
rect 502154 344927 502210 344936
rect 502168 338881 502196 344927
rect 502154 338872 502210 338881
rect 502154 338807 502210 338816
rect 502062 337512 502118 337521
rect 502062 337447 502118 337456
rect 501970 325680 502026 325689
rect 501970 325615 502026 325624
rect 501984 315897 502012 325615
rect 501970 315888 502026 315897
rect 501970 315823 502026 315832
rect 501970 308544 502026 308553
rect 501970 308479 502026 308488
rect 501984 290465 502012 308479
rect 501970 290456 502026 290465
rect 501970 290391 502026 290400
rect 501970 290320 502026 290329
rect 501970 290255 501972 290264
rect 502024 290255 502026 290264
rect 501972 290226 502024 290232
rect 501970 290184 502026 290193
rect 501970 290119 502026 290128
rect 501984 282441 502012 290119
rect 501970 282432 502026 282441
rect 501970 282367 502026 282376
rect 501970 282296 502026 282305
rect 501970 282231 501972 282240
rect 502024 282231 502026 282240
rect 501972 282202 502024 282208
rect 501970 281480 502026 281489
rect 501970 281415 502026 281424
rect 501984 278458 502012 281415
rect 501972 278452 502024 278458
rect 501972 278394 502024 278400
rect 501972 278316 502024 278322
rect 501972 278258 502024 278264
rect 501984 275097 502012 278258
rect 501970 275088 502026 275097
rect 501970 275023 502026 275032
rect 501970 273184 502026 273193
rect 501970 273119 502026 273128
rect 501984 272814 502012 273119
rect 501972 272808 502024 272814
rect 501972 272750 502024 272756
rect 501972 272672 502024 272678
rect 501970 272640 501972 272649
rect 502024 272640 502026 272649
rect 501970 272575 502026 272584
rect 501972 272536 502024 272542
rect 501970 272504 501972 272513
rect 502024 272504 502026 272513
rect 501970 272439 502026 272448
rect 501972 272400 502024 272406
rect 501970 272368 501972 272377
rect 502024 272368 502026 272377
rect 501970 272303 502026 272312
rect 501972 270904 502024 270910
rect 501970 270872 501972 270881
rect 502024 270872 502026 270881
rect 501970 270807 502026 270816
rect 501970 270464 502026 270473
rect 501970 270399 501972 270408
rect 502024 270399 502026 270408
rect 501972 270370 502024 270376
rect 501970 268288 502026 268297
rect 501970 268223 502026 268232
rect 501984 267170 502012 268223
rect 501972 267164 502024 267170
rect 501972 267106 502024 267112
rect 501970 267064 502026 267073
rect 501970 266999 501972 267008
rect 502024 266999 502026 267008
rect 501972 266970 502024 266976
rect 501970 263528 502026 263537
rect 501970 263463 502026 263472
rect 501880 158840 501932 158846
rect 501880 158782 501932 158788
rect 501880 158704 501932 158710
rect 501880 158646 501932 158652
rect 501892 155582 501920 158646
rect 501880 155576 501932 155582
rect 501880 155518 501932 155524
rect 501880 155440 501932 155446
rect 501880 155382 501932 155388
rect 501892 155281 501920 155382
rect 501878 155272 501934 155281
rect 501878 155207 501934 155216
rect 501880 155168 501932 155174
rect 501880 155110 501932 155116
rect 501892 141710 501920 155110
rect 501880 141704 501932 141710
rect 501880 141646 501932 141652
rect 501878 140584 501934 140593
rect 501878 140519 501880 140528
rect 501932 140519 501934 140528
rect 501880 140490 501932 140496
rect 501878 140448 501934 140457
rect 501878 140383 501880 140392
rect 501932 140383 501934 140392
rect 501880 140354 501932 140360
rect 501878 140312 501934 140321
rect 501878 140247 501880 140256
rect 501932 140247 501934 140256
rect 501880 140218 501932 140224
rect 501878 140176 501934 140185
rect 501878 140111 501880 140120
rect 501932 140111 501934 140120
rect 501880 140082 501932 140088
rect 501878 140040 501934 140049
rect 501878 139975 501880 139984
rect 501932 139975 501934 139984
rect 501880 139946 501932 139952
rect 501878 138816 501934 138825
rect 501878 138751 501934 138760
rect 501892 138106 501920 138751
rect 501880 138100 501932 138106
rect 501880 138042 501932 138048
rect 501878 137864 501934 137873
rect 501878 137799 501880 137808
rect 501932 137799 501934 137808
rect 501880 137770 501932 137776
rect 501880 137080 501932 137086
rect 501878 137048 501880 137057
rect 501932 137048 501934 137057
rect 501878 136983 501934 136992
rect 501880 136944 501932 136950
rect 501880 136886 501932 136892
rect 501892 136785 501920 136886
rect 501878 136776 501934 136785
rect 501878 136711 501934 136720
rect 501880 135516 501932 135522
rect 501880 135458 501932 135464
rect 501892 127362 501920 135458
rect 501880 127356 501932 127362
rect 501880 127298 501932 127304
rect 501880 127220 501932 127226
rect 501880 127162 501932 127168
rect 501788 124636 501840 124642
rect 501788 124578 501840 124584
rect 501788 123888 501840 123894
rect 501788 123830 501840 123836
rect 501800 121242 501828 123830
rect 501788 121236 501840 121242
rect 501788 121178 501840 121184
rect 501892 120737 501920 127162
rect 501878 120728 501934 120737
rect 501878 120663 501934 120672
rect 501984 13666 502012 263463
rect 502076 124953 502104 337447
rect 502154 320376 502210 320385
rect 502154 320311 502210 320320
rect 502168 209370 502196 320311
rect 502246 290048 502302 290057
rect 502246 289983 502302 289992
rect 502260 278322 502288 289983
rect 502248 278316 502300 278322
rect 502248 278258 502300 278264
rect 502246 278216 502302 278225
rect 502246 278151 502302 278160
rect 502260 277846 502288 278151
rect 502248 277840 502300 277846
rect 502248 277782 502300 277788
rect 502248 277636 502300 277642
rect 502248 277578 502300 277584
rect 502156 209364 502208 209370
rect 502156 209306 502208 209312
rect 502154 209264 502210 209273
rect 502154 209199 502210 209208
rect 502168 198121 502196 209199
rect 502154 198112 502210 198121
rect 502154 198047 502210 198056
rect 502156 197736 502208 197742
rect 502156 197678 502208 197684
rect 502168 141846 502196 197678
rect 502156 141840 502208 141846
rect 502156 141782 502208 141788
rect 502156 141704 502208 141710
rect 502156 141646 502208 141652
rect 502168 127362 502196 141646
rect 502156 127356 502208 127362
rect 502156 127298 502208 127304
rect 502156 127152 502208 127158
rect 502156 127094 502208 127100
rect 502062 124944 502118 124953
rect 502062 124879 502118 124888
rect 502168 123865 502196 127094
rect 502154 123856 502210 123865
rect 502154 123791 502210 123800
rect 502156 123752 502208 123758
rect 502154 123720 502156 123729
rect 502208 123720 502210 123729
rect 502154 123655 502210 123664
rect 502062 122768 502118 122777
rect 502062 122703 502118 122712
rect 502076 121009 502104 122703
rect 502062 121000 502118 121009
rect 502062 120935 502118 120944
rect 502064 118584 502116 118590
rect 502064 118526 502116 118532
rect 502076 118289 502104 118526
rect 502062 118280 502118 118289
rect 502062 118215 502118 118224
rect 501972 13660 502024 13666
rect 501972 13602 502024 13608
rect 501696 3868 501748 3874
rect 501696 3810 501748 3816
rect 502260 3806 502288 277578
rect 502352 155242 502380 583782
rect 502430 415576 502486 415585
rect 502430 415511 502486 415520
rect 502340 155236 502392 155242
rect 502340 155178 502392 155184
rect 502340 155100 502392 155106
rect 502340 155042 502392 155048
rect 502352 148986 502380 155042
rect 502340 148980 502392 148986
rect 502340 148922 502392 148928
rect 502338 148880 502394 148889
rect 502338 148815 502340 148824
rect 502392 148815 502394 148824
rect 502340 148786 502392 148792
rect 502338 147520 502394 147529
rect 502338 147455 502340 147464
rect 502392 147455 502394 147464
rect 502340 147426 502392 147432
rect 502340 147280 502392 147286
rect 502338 147248 502340 147257
rect 502392 147248 502394 147257
rect 502338 147183 502394 147192
rect 502338 146976 502394 146985
rect 502338 146911 502394 146920
rect 502352 138417 502380 146911
rect 502338 138408 502394 138417
rect 502338 138343 502394 138352
rect 502340 138304 502392 138310
rect 502338 138272 502340 138281
rect 502392 138272 502394 138281
rect 502338 138207 502394 138216
rect 502340 137488 502392 137494
rect 502338 137456 502340 137465
rect 502392 137456 502394 137465
rect 502338 137391 502394 137400
rect 502338 137320 502394 137329
rect 502338 137255 502394 137264
rect 502352 113898 502380 137255
rect 502340 113892 502392 113898
rect 502340 113834 502392 113840
rect 502444 6458 502472 415511
rect 502536 316849 502564 700606
rect 504456 700392 504508 700398
rect 504456 700334 504508 700340
rect 502616 667956 502668 667962
rect 502616 667898 502668 667904
rect 502628 401441 502656 667898
rect 502984 583500 503036 583506
rect 502984 583442 503036 583448
rect 502706 582856 502762 582865
rect 502706 582791 502762 582800
rect 502720 575521 502748 582791
rect 502706 575512 502762 575521
rect 502706 575447 502762 575456
rect 502890 433256 502946 433265
rect 502890 433191 502946 433200
rect 502904 425105 502932 433191
rect 502890 425096 502946 425105
rect 502890 425031 502946 425040
rect 502614 401432 502670 401441
rect 502614 401367 502670 401376
rect 502614 397896 502670 397905
rect 502614 397831 502670 397840
rect 502522 316840 502578 316849
rect 502522 316775 502578 316784
rect 502522 302968 502578 302977
rect 502522 302903 502578 302912
rect 502432 6452 502484 6458
rect 502432 6394 502484 6400
rect 502432 6248 502484 6254
rect 502432 6190 502484 6196
rect 502248 3800 502300 3806
rect 502248 3742 502300 3748
rect 502444 480 502472 6190
rect 502536 4146 502564 302903
rect 502628 124778 502656 397831
rect 502706 383752 502762 383761
rect 502706 383687 502762 383696
rect 502616 124772 502668 124778
rect 502616 124714 502668 124720
rect 502614 124672 502670 124681
rect 502614 124607 502670 124616
rect 502628 122233 502656 124607
rect 502614 122224 502670 122233
rect 502614 122159 502670 122168
rect 502720 115462 502748 383687
rect 502798 359272 502854 359281
rect 502798 359207 502854 359216
rect 502812 121310 502840 359207
rect 502890 327448 502946 327457
rect 502890 327383 502946 327392
rect 502904 121378 502932 327383
rect 502996 166734 503024 583442
rect 503352 583296 503404 583302
rect 503352 583238 503404 583244
rect 503076 583228 503128 583234
rect 503076 583170 503128 583176
rect 503088 192642 503116 583170
rect 503260 582888 503312 582894
rect 503260 582830 503312 582836
rect 503168 582684 503220 582690
rect 503168 582626 503220 582632
rect 503180 393310 503208 582626
rect 503272 440230 503300 582830
rect 503364 534070 503392 583238
rect 504364 581392 504416 581398
rect 504364 581334 504416 581340
rect 503902 580408 503958 580417
rect 503902 580343 503958 580352
rect 503718 579728 503774 579737
rect 503718 579663 503774 579672
rect 503732 574161 503760 579663
rect 503718 574152 503774 574161
rect 503718 574087 503774 574096
rect 503810 567080 503866 567089
rect 503810 567015 503866 567024
rect 503824 565894 503852 567015
rect 503812 565888 503864 565894
rect 503812 565830 503864 565836
rect 503916 565706 503944 580343
rect 503732 565678 503944 565706
rect 503352 534064 503404 534070
rect 503352 534006 503404 534012
rect 503732 514758 503760 565678
rect 503810 563544 503866 563553
rect 503810 563479 503866 563488
rect 503824 563106 503852 563479
rect 503812 563100 503864 563106
rect 503812 563042 503864 563048
rect 503810 521112 503866 521121
rect 503810 521047 503866 521056
rect 503720 514752 503772 514758
rect 503720 514694 503772 514700
rect 503720 505164 503772 505170
rect 503720 505106 503772 505112
rect 503732 475794 503760 505106
rect 503720 475788 503772 475794
rect 503720 475730 503772 475736
rect 503534 471880 503590 471889
rect 503534 471815 503590 471824
rect 503548 470626 503576 471815
rect 503536 470620 503588 470626
rect 503536 470562 503588 470568
rect 503720 461440 503772 461446
rect 503720 461382 503772 461388
rect 503732 456482 503760 461382
rect 503720 456476 503772 456482
rect 503720 456418 503772 456424
rect 503720 447160 503772 447166
rect 503720 447102 503772 447108
rect 503260 440224 503312 440230
rect 503260 440166 503312 440172
rect 503732 437442 503760 447102
rect 503720 437436 503772 437442
rect 503720 437378 503772 437384
rect 503720 427848 503772 427854
rect 503720 427790 503772 427796
rect 503258 419112 503314 419121
rect 503258 419047 503314 419056
rect 503272 418266 503300 419047
rect 503260 418260 503312 418266
rect 503260 418202 503312 418208
rect 503732 418130 503760 427790
rect 503720 418124 503772 418130
rect 503720 418066 503772 418072
rect 503720 408536 503772 408542
rect 503720 408478 503772 408484
rect 503168 393304 503220 393310
rect 503168 393246 503220 393252
rect 503442 341592 503498 341601
rect 503442 341527 503498 341536
rect 503456 340950 503484 341527
rect 503444 340944 503496 340950
rect 503444 340886 503496 340892
rect 503166 299432 503222 299441
rect 503166 299367 503222 299376
rect 503076 192636 503128 192642
rect 503076 192578 503128 192584
rect 503074 192536 503130 192545
rect 503074 192471 503130 192480
rect 503088 189825 503116 192471
rect 503074 189816 503130 189825
rect 503074 189751 503130 189760
rect 503076 189712 503128 189718
rect 503076 189654 503128 189660
rect 503088 186697 503116 189654
rect 503074 186688 503130 186697
rect 503074 186623 503130 186632
rect 503074 186552 503130 186561
rect 503074 186487 503130 186496
rect 503088 181830 503116 186487
rect 503076 181824 503128 181830
rect 503076 181766 503128 181772
rect 503074 180160 503130 180169
rect 503074 180095 503130 180104
rect 503088 173097 503116 180095
rect 503074 173088 503130 173097
rect 503074 173023 503130 173032
rect 503076 172984 503128 172990
rect 503076 172926 503128 172932
rect 502984 166728 503036 166734
rect 502984 166670 503036 166676
rect 502982 166424 503038 166433
rect 502982 166359 502984 166368
rect 503036 166359 503038 166368
rect 502984 166330 503036 166336
rect 502984 165640 503036 165646
rect 502984 165582 503036 165588
rect 502996 165481 503024 165582
rect 502982 165472 503038 165481
rect 502982 165407 503038 165416
rect 502982 165064 503038 165073
rect 502982 164999 503038 165008
rect 502996 164966 503024 164999
rect 502984 164960 503036 164966
rect 502984 164902 503036 164908
rect 502982 163840 503038 163849
rect 502982 163775 502984 163784
rect 503036 163775 503038 163784
rect 502984 163746 503036 163752
rect 502982 162888 503038 162897
rect 502982 162823 502984 162832
rect 503036 162823 503038 162832
rect 502984 162794 503036 162800
rect 502982 162480 503038 162489
rect 502982 162415 502984 162424
rect 503036 162415 503038 162424
rect 502984 162386 503036 162392
rect 502982 162344 503038 162353
rect 502982 162279 503038 162288
rect 502996 162178 503024 162279
rect 502984 162172 503036 162178
rect 502984 162114 503036 162120
rect 502982 162072 503038 162081
rect 502982 162007 503038 162016
rect 502892 121372 502944 121378
rect 502892 121314 502944 121320
rect 502800 121304 502852 121310
rect 502800 121246 502852 121252
rect 502996 116754 503024 162007
rect 502984 116748 503036 116754
rect 502984 116690 503036 116696
rect 502708 115456 502760 115462
rect 502708 115398 502760 115404
rect 502524 4140 502576 4146
rect 502524 4082 502576 4088
rect 503088 3194 503116 172926
rect 503180 122058 503208 299367
rect 503258 271144 503314 271153
rect 503258 271079 503314 271088
rect 503168 122052 503220 122058
rect 503168 121994 503220 122000
rect 503272 118250 503300 271079
rect 503442 270600 503498 270609
rect 503442 270535 503498 270544
rect 503350 270328 503406 270337
rect 503350 270263 503406 270272
rect 503364 259570 503392 270263
rect 503456 260137 503484 270535
rect 503628 267164 503680 267170
rect 503628 267106 503680 267112
rect 503534 262440 503590 262449
rect 503534 262375 503590 262384
rect 503442 260128 503498 260137
rect 503442 260063 503498 260072
rect 503548 259593 503576 262375
rect 503640 260273 503668 267106
rect 503626 260264 503682 260273
rect 503626 260199 503682 260208
rect 503534 259584 503590 259593
rect 503364 259542 503484 259570
rect 503350 259448 503406 259457
rect 503350 259383 503406 259392
rect 503364 255377 503392 259383
rect 503456 256737 503484 259542
rect 503534 259519 503590 259528
rect 503534 258768 503590 258777
rect 503534 258703 503590 258712
rect 503442 256728 503498 256737
rect 503442 256663 503498 256672
rect 503548 256193 503576 258703
rect 503534 256184 503590 256193
rect 503534 256119 503590 256128
rect 503350 255368 503406 255377
rect 503350 255303 503406 255312
rect 503626 255096 503682 255105
rect 503626 255031 503682 255040
rect 503534 254960 503590 254969
rect 503534 254895 503590 254904
rect 503352 254652 503404 254658
rect 503352 254594 503404 254600
rect 503364 254561 503392 254594
rect 503350 254552 503406 254561
rect 503350 254487 503406 254496
rect 503350 254144 503406 254153
rect 503350 254079 503406 254088
rect 503364 242146 503392 254079
rect 503444 253224 503496 253230
rect 503442 253192 503444 253201
rect 503496 253192 503498 253201
rect 503442 253127 503498 253136
rect 503442 253056 503498 253065
rect 503442 252991 503444 253000
rect 503496 252991 503498 253000
rect 503444 252962 503496 252968
rect 503442 246664 503498 246673
rect 503442 246599 503498 246608
rect 503456 245342 503484 246599
rect 503444 245336 503496 245342
rect 503444 245278 503496 245284
rect 503444 245200 503496 245206
rect 503444 245142 503496 245148
rect 503352 242140 503404 242146
rect 503352 242082 503404 242088
rect 503456 242026 503484 245142
rect 503548 244225 503576 254895
rect 503534 244216 503590 244225
rect 503534 244151 503590 244160
rect 503534 243128 503590 243137
rect 503534 243063 503590 243072
rect 503364 241998 503484 242026
rect 503364 229129 503392 241998
rect 503444 241936 503496 241942
rect 503444 241878 503496 241884
rect 503456 241505 503484 241878
rect 503442 241496 503498 241505
rect 503548 241482 503576 243063
rect 503640 241602 503668 255031
rect 503628 241596 503680 241602
rect 503628 241538 503680 241544
rect 503548 241454 503668 241482
rect 503442 241431 503498 241440
rect 503442 239592 503498 239601
rect 503442 239527 503498 239536
rect 503456 238882 503484 239527
rect 503444 238876 503496 238882
rect 503444 238818 503496 238824
rect 503442 238096 503498 238105
rect 503442 238031 503498 238040
rect 503350 229120 503406 229129
rect 503350 229055 503406 229064
rect 503350 228984 503406 228993
rect 503350 228919 503406 228928
rect 503260 118244 503312 118250
rect 503260 118186 503312 118192
rect 503364 118182 503392 228919
rect 503456 225554 503484 238031
rect 503534 237688 503590 237697
rect 503534 237623 503590 237632
rect 503548 235793 503576 237623
rect 503534 235784 503590 235793
rect 503534 235719 503590 235728
rect 503534 235512 503590 235521
rect 503534 235447 503590 235456
rect 503548 233646 503576 235447
rect 503640 235278 503668 241454
rect 503628 235272 503680 235278
rect 503628 235214 503680 235220
rect 503536 233640 503588 233646
rect 503536 233582 503588 233588
rect 503534 233200 503590 233209
rect 503534 233135 503590 233144
rect 503444 225548 503496 225554
rect 503444 225490 503496 225496
rect 503442 225448 503498 225457
rect 503442 225383 503498 225392
rect 503456 225010 503484 225383
rect 503444 225004 503496 225010
rect 503444 224946 503496 224952
rect 503442 224904 503498 224913
rect 503442 224839 503498 224848
rect 503456 222057 503484 224839
rect 503442 222048 503498 222057
rect 503442 221983 503498 221992
rect 503442 221912 503498 221921
rect 503442 221847 503444 221856
rect 503496 221847 503498 221856
rect 503444 221818 503496 221824
rect 503442 221504 503498 221513
rect 503442 221439 503498 221448
rect 503456 211857 503484 221439
rect 503548 220130 503576 233135
rect 503628 227452 503680 227458
rect 503628 227394 503680 227400
rect 503640 226545 503668 227394
rect 503626 226536 503682 226545
rect 503626 226471 503682 226480
rect 503626 225176 503682 225185
rect 503626 225111 503682 225120
rect 503640 221542 503668 225111
rect 503628 221536 503680 221542
rect 503628 221478 503680 221484
rect 503628 221264 503680 221270
rect 503628 221206 503680 221212
rect 503640 220425 503668 221206
rect 503626 220416 503682 220425
rect 503626 220351 503682 220360
rect 503626 220280 503682 220289
rect 503626 220215 503628 220224
rect 503680 220215 503682 220224
rect 503628 220186 503680 220192
rect 503548 220102 503668 220130
rect 503536 220040 503588 220046
rect 503536 219982 503588 219988
rect 503548 219881 503576 219982
rect 503534 219872 503590 219881
rect 503534 219807 503590 219816
rect 503536 219700 503588 219706
rect 503536 219642 503588 219648
rect 503548 215937 503576 219642
rect 503640 216073 503668 220102
rect 503626 216064 503682 216073
rect 503626 215999 503682 216008
rect 503534 215928 503590 215937
rect 503534 215863 503590 215872
rect 503534 215792 503590 215801
rect 503534 215727 503590 215736
rect 503442 211848 503498 211857
rect 503442 211783 503498 211792
rect 503442 211304 503498 211313
rect 503442 211239 503498 211248
rect 503456 121922 503484 211239
rect 503548 205034 503576 215727
rect 503628 210792 503680 210798
rect 503626 210760 503628 210769
rect 503680 210760 503682 210769
rect 503626 210695 503682 210704
rect 503626 207768 503682 207777
rect 503626 207703 503682 207712
rect 503640 207058 503668 207703
rect 503628 207052 503680 207058
rect 503628 206994 503680 207000
rect 503548 205006 503668 205034
rect 503534 204912 503590 204921
rect 503534 204847 503536 204856
rect 503588 204847 503590 204856
rect 503536 204818 503588 204824
rect 503534 204096 503590 204105
rect 503534 204031 503590 204040
rect 503548 197441 503576 204031
rect 503640 199510 503668 205006
rect 503628 199504 503680 199510
rect 503628 199446 503680 199452
rect 503628 199368 503680 199374
rect 503626 199336 503628 199345
rect 503680 199336 503682 199345
rect 503626 199271 503682 199280
rect 503534 197432 503590 197441
rect 503534 197367 503590 197376
rect 503626 196888 503682 196897
rect 503626 196823 503682 196832
rect 503536 196240 503588 196246
rect 503534 196208 503536 196217
rect 503588 196208 503590 196217
rect 503534 196143 503590 196152
rect 503534 194440 503590 194449
rect 503534 194375 503536 194384
rect 503588 194375 503590 194384
rect 503536 194346 503588 194352
rect 503534 193624 503590 193633
rect 503534 193559 503590 193568
rect 503444 121916 503496 121922
rect 503444 121858 503496 121864
rect 503548 118318 503576 193559
rect 503640 186998 503668 196823
rect 503628 186992 503680 186998
rect 503628 186934 503680 186940
rect 503626 186824 503682 186833
rect 503626 186759 503682 186768
rect 503640 173233 503668 186759
rect 503626 173224 503682 173233
rect 503626 173159 503682 173168
rect 503626 173088 503682 173097
rect 503626 173023 503682 173032
rect 503640 169250 503668 173023
rect 503628 169244 503680 169250
rect 503628 169186 503680 169192
rect 503626 169144 503682 169153
rect 503626 169079 503682 169088
rect 503640 160750 503668 169079
rect 503628 160744 503680 160750
rect 503628 160686 503680 160692
rect 503628 158840 503680 158846
rect 503628 158782 503680 158788
rect 503640 132530 503668 158782
rect 503732 148034 503760 408478
rect 503824 185881 503852 521047
rect 503904 514752 503956 514758
rect 503904 514694 503956 514700
rect 503916 505170 503944 514694
rect 503904 505164 503956 505170
rect 503904 505106 503956 505112
rect 504178 500168 504234 500177
rect 504178 500103 504234 500112
rect 503902 482488 503958 482497
rect 503902 482423 503958 482432
rect 503810 185872 503866 185881
rect 503810 185807 503866 185816
rect 503810 183560 503866 183569
rect 503810 183495 503866 183504
rect 503824 180305 503852 183495
rect 503810 180296 503866 180305
rect 503810 180231 503866 180240
rect 503812 180192 503864 180198
rect 503810 180160 503812 180169
rect 503864 180160 503866 180169
rect 503810 180095 503866 180104
rect 503810 179480 503866 179489
rect 503810 179415 503866 179424
rect 503720 148028 503772 148034
rect 503720 147970 503772 147976
rect 503718 147928 503774 147937
rect 503718 147863 503774 147872
rect 503732 147694 503760 147863
rect 503720 147688 503772 147694
rect 503720 147630 503772 147636
rect 503720 147008 503772 147014
rect 503720 146950 503772 146956
rect 503732 137329 503760 146950
rect 503718 137320 503774 137329
rect 503718 137255 503774 137264
rect 503720 136332 503772 136338
rect 503720 136274 503772 136280
rect 503732 135017 503760 136274
rect 503718 135008 503774 135017
rect 503718 134943 503774 134952
rect 503720 133952 503772 133958
rect 503718 133920 503720 133929
rect 503772 133920 503774 133929
rect 503718 133855 503774 133864
rect 503718 133784 503774 133793
rect 503718 133719 503774 133728
rect 503628 132524 503680 132530
rect 503628 132466 503680 132472
rect 503732 131102 503760 133719
rect 503720 131096 503772 131102
rect 503720 131038 503772 131044
rect 503718 130656 503774 130665
rect 503718 130591 503720 130600
rect 503772 130591 503774 130600
rect 503720 130562 503772 130568
rect 503626 130248 503682 130257
rect 503626 130183 503682 130192
rect 503640 127838 503668 130183
rect 503720 130008 503772 130014
rect 503720 129950 503772 129956
rect 503628 127832 503680 127838
rect 503628 127774 503680 127780
rect 503628 127696 503680 127702
rect 503628 127638 503680 127644
rect 503640 124953 503668 127638
rect 503626 124944 503682 124953
rect 503626 124879 503682 124888
rect 503628 124840 503680 124846
rect 503628 124782 503680 124788
rect 503640 121417 503668 124782
rect 503732 124001 503760 129950
rect 503718 123992 503774 124001
rect 503718 123927 503774 123936
rect 503824 122602 503852 179415
rect 503916 165889 503944 482423
rect 504088 475788 504140 475794
rect 504088 475730 504140 475736
rect 504100 461446 504128 475730
rect 504088 461440 504140 461446
rect 504088 461382 504140 461388
rect 504088 456476 504140 456482
rect 504088 456418 504140 456424
rect 504100 447166 504128 456418
rect 504088 447160 504140 447166
rect 504088 447102 504140 447108
rect 503994 440328 504050 440337
rect 503994 440263 504050 440272
rect 503902 165880 503958 165889
rect 503902 165815 503958 165824
rect 503902 165608 503958 165617
rect 503902 165543 503904 165552
rect 503956 165543 503958 165552
rect 503904 165514 503956 165520
rect 503902 163704 503958 163713
rect 503902 163639 503958 163648
rect 503916 161809 503944 163639
rect 503902 161800 503958 161809
rect 503902 161735 503958 161744
rect 503904 160744 503956 160750
rect 503904 160686 503956 160692
rect 503812 122596 503864 122602
rect 503812 122538 503864 122544
rect 503626 121408 503682 121417
rect 503626 121343 503682 121352
rect 503536 118312 503588 118318
rect 503536 118254 503588 118260
rect 503352 118176 503404 118182
rect 503352 118118 503404 118124
rect 503720 79688 503772 79694
rect 503720 79630 503772 79636
rect 503732 75970 503760 79630
rect 503640 75942 503760 75970
rect 503640 73234 503668 75942
rect 503628 73228 503680 73234
rect 503628 73170 503680 73176
rect 503916 17338 503944 160686
rect 504008 157457 504036 440263
rect 504086 436792 504142 436801
rect 504086 436727 504142 436736
rect 504100 158817 504128 436727
rect 504192 388385 504220 500103
rect 504272 437436 504324 437442
rect 504272 437378 504324 437384
rect 504284 427854 504312 437378
rect 504272 427848 504324 427854
rect 504272 427790 504324 427796
rect 504272 418124 504324 418130
rect 504272 418066 504324 418072
rect 504284 408542 504312 418066
rect 504272 408536 504324 408542
rect 504272 408478 504324 408484
rect 504178 388376 504234 388385
rect 504178 388311 504234 388320
rect 504270 380216 504326 380225
rect 504270 380151 504326 380160
rect 504178 376952 504234 376961
rect 504178 376887 504234 376896
rect 504192 376786 504220 376887
rect 504180 376780 504232 376786
rect 504180 376722 504232 376728
rect 504178 373416 504234 373425
rect 504178 373351 504234 373360
rect 504192 372638 504220 373351
rect 504180 372632 504232 372638
rect 504180 372574 504232 372580
rect 504178 352200 504234 352209
rect 504178 352135 504234 352144
rect 504192 351966 504220 352135
rect 504180 351960 504232 351966
rect 504180 351902 504232 351908
rect 504178 345128 504234 345137
rect 504178 345063 504234 345072
rect 504192 277642 504220 345063
rect 504180 277636 504232 277642
rect 504180 277578 504232 277584
rect 504180 274712 504232 274718
rect 504178 274680 504180 274689
rect 504232 274680 504234 274689
rect 504178 274615 504234 274624
rect 504180 274576 504232 274582
rect 504180 274518 504232 274524
rect 504086 158808 504142 158817
rect 504086 158743 504142 158752
rect 504086 158536 504142 158545
rect 504086 158471 504142 158480
rect 503994 157448 504050 157457
rect 503994 157383 504050 157392
rect 504100 155088 504128 158471
rect 504008 155060 504128 155088
rect 504008 116113 504036 155060
rect 504086 155000 504142 155009
rect 504086 154935 504142 154944
rect 504100 148646 504128 154935
rect 504088 148640 504140 148646
rect 504088 148582 504140 148588
rect 504088 146192 504140 146198
rect 504086 146160 504088 146169
rect 504140 146160 504142 146169
rect 504086 146095 504142 146104
rect 504086 146024 504142 146033
rect 504086 145959 504088 145968
rect 504140 145959 504142 145968
rect 504088 145930 504140 145936
rect 504086 145888 504142 145897
rect 504086 145823 504142 145832
rect 504100 144498 504128 145823
rect 504088 144492 504140 144498
rect 504088 144434 504140 144440
rect 504086 144392 504142 144401
rect 504086 144327 504142 144336
rect 503994 116104 504050 116113
rect 503994 116039 504050 116048
rect 503994 87680 504050 87689
rect 503994 87615 504050 87624
rect 504008 77353 504036 87615
rect 503994 77344 504050 77353
rect 503994 77279 504050 77288
rect 503994 49056 504050 49065
rect 503994 48991 504050 49000
rect 504008 38865 504036 48991
rect 503994 38856 504050 38865
rect 503994 38791 504050 38800
rect 503904 17332 503956 17338
rect 503904 17274 503956 17280
rect 504100 15910 504128 144327
rect 504192 17474 504220 274518
rect 504284 118114 504312 380151
rect 504376 148782 504404 581334
rect 504468 534177 504496 700334
rect 507124 638988 507176 638994
rect 507124 638930 507176 638936
rect 506480 584860 506532 584866
rect 506480 584802 506532 584808
rect 505284 584452 505336 584458
rect 505284 584394 505336 584400
rect 504914 582040 504970 582049
rect 504914 581975 504970 581984
rect 504928 581233 504956 581975
rect 505006 581632 505062 581641
rect 505006 581567 505062 581576
rect 505190 581632 505246 581641
rect 505190 581567 505246 581576
rect 504914 581224 504970 581233
rect 504914 581159 504970 581168
rect 505020 581097 505048 581567
rect 505100 581528 505152 581534
rect 505100 581470 505152 581476
rect 505006 581088 505062 581097
rect 505006 581023 505062 581032
rect 504916 556300 504968 556306
rect 504916 556242 504968 556248
rect 504928 556209 504956 556242
rect 504914 556200 504970 556209
rect 504914 556135 504970 556144
rect 504822 552120 504878 552129
rect 504822 552055 504824 552064
rect 504876 552055 504878 552064
rect 504824 552026 504876 552032
rect 505006 549400 505062 549409
rect 505006 549335 505008 549344
rect 505060 549335 505062 549344
rect 505008 549306 505060 549312
rect 504454 534168 504510 534177
rect 504454 534103 504510 534112
rect 505006 528184 505062 528193
rect 505006 528119 505062 528128
rect 505020 527202 505048 528119
rect 505008 527196 505060 527202
rect 505008 527138 505060 527144
rect 504454 524648 504510 524657
rect 504454 524583 504510 524592
rect 504468 510610 504496 524583
rect 504456 510604 504508 510610
rect 504456 510546 504508 510552
rect 504454 496632 504510 496641
rect 504454 496567 504510 496576
rect 504468 485858 504496 496567
rect 505008 492720 505060 492726
rect 505006 492688 505008 492697
rect 505060 492688 505062 492697
rect 505006 492623 505062 492632
rect 504456 485852 504508 485858
rect 504456 485794 504508 485800
rect 505006 478952 505062 478961
rect 505006 478887 505008 478896
rect 505060 478887 505062 478896
rect 505008 478858 505060 478864
rect 504546 454200 504602 454209
rect 504546 454135 504602 454144
rect 504560 454102 504588 454135
rect 504548 454096 504600 454102
rect 504548 454038 504600 454044
rect 504638 426184 504694 426193
rect 504638 426119 504694 426128
rect 504546 390824 504602 390833
rect 504546 390759 504602 390768
rect 504560 390590 504588 390759
rect 504548 390584 504600 390590
rect 504548 390526 504600 390532
rect 504548 369912 504600 369918
rect 504546 369880 504548 369889
rect 504600 369880 504602 369889
rect 504546 369815 504602 369824
rect 504548 362840 504600 362846
rect 504546 362808 504548 362817
rect 504600 362808 504602 362817
rect 504546 362743 504602 362752
rect 504546 347576 504602 347585
rect 504546 347511 504602 347520
rect 504560 338881 504588 347511
rect 504546 338872 504602 338881
rect 504546 338807 504602 338816
rect 504546 334520 504602 334529
rect 504546 334455 504602 334464
rect 504454 330984 504510 330993
rect 504454 330919 504510 330928
rect 504468 329866 504496 330919
rect 504456 329860 504508 329866
rect 504456 329802 504508 329808
rect 504456 324284 504508 324290
rect 504456 324226 504508 324232
rect 504468 323921 504496 324226
rect 504454 323912 504510 323921
rect 504454 323847 504510 323856
rect 504454 310040 504510 310049
rect 504454 309975 504510 309984
rect 504468 309194 504496 309975
rect 504456 309188 504508 309194
rect 504456 309130 504508 309136
rect 504454 306504 504510 306513
rect 504454 306439 504510 306448
rect 504468 306406 504496 306439
rect 504456 306400 504508 306406
rect 504456 306342 504508 306348
rect 504456 296676 504508 296682
rect 504456 296618 504508 296624
rect 504468 295905 504496 296618
rect 504454 295896 504510 295905
rect 504454 295831 504510 295840
rect 504454 288824 504510 288833
rect 504454 288759 504510 288768
rect 504364 148776 504416 148782
rect 504364 148718 504416 148724
rect 504364 148640 504416 148646
rect 504364 148582 504416 148588
rect 504376 122738 504404 148582
rect 504364 122732 504416 122738
rect 504364 122674 504416 122680
rect 504272 118108 504324 118114
rect 504272 118050 504324 118056
rect 504468 86290 504496 288759
rect 504560 149054 504588 334455
rect 504652 246537 504680 426119
rect 505006 404968 505062 404977
rect 505006 404903 505062 404912
rect 505020 402830 505048 404903
rect 505008 402824 505060 402830
rect 505008 402766 505060 402772
rect 504822 348664 504878 348673
rect 504822 348599 504878 348608
rect 504730 307184 504786 307193
rect 504730 307119 504786 307128
rect 504744 297401 504772 307119
rect 504730 297392 504786 297401
rect 504730 297327 504786 297336
rect 504730 281752 504786 281761
rect 504730 281687 504786 281696
rect 504744 274582 504772 281687
rect 504732 274576 504784 274582
rect 504732 274518 504784 274524
rect 504730 271824 504786 271833
rect 504730 271759 504786 271768
rect 504744 267073 504772 271759
rect 504730 267064 504786 267073
rect 504730 266999 504786 267008
rect 504730 257000 504786 257009
rect 504730 256935 504786 256944
rect 504638 246528 504694 246537
rect 504638 246463 504694 246472
rect 504640 246424 504692 246430
rect 504640 246366 504692 246372
rect 504652 244769 504680 246366
rect 504638 244760 504694 244769
rect 504638 244695 504694 244704
rect 504638 236056 504694 236065
rect 504638 235991 504640 236000
rect 504692 235991 504694 236000
rect 504640 235962 504692 235968
rect 504640 235272 504692 235278
rect 504640 235214 504692 235220
rect 504548 149048 504600 149054
rect 504548 148990 504600 148996
rect 504548 148776 504600 148782
rect 504548 148718 504600 148724
rect 504560 147665 504588 148718
rect 504546 147656 504602 147665
rect 504546 147591 504602 147600
rect 504548 147416 504600 147422
rect 504548 147358 504600 147364
rect 504560 143993 504588 147358
rect 504546 143984 504602 143993
rect 504546 143919 504602 143928
rect 504548 143676 504600 143682
rect 504548 143618 504600 143624
rect 504560 143585 504588 143618
rect 504546 143576 504602 143585
rect 504546 143511 504602 143520
rect 504546 143440 504602 143449
rect 504546 143375 504548 143384
rect 504600 143375 504602 143384
rect 504548 143346 504600 143352
rect 504546 140856 504602 140865
rect 504546 140791 504602 140800
rect 504560 118386 504588 140791
rect 504548 118380 504600 118386
rect 504548 118322 504600 118328
rect 504546 118280 504602 118289
rect 504546 118215 504602 118224
rect 504560 106049 504588 118215
rect 504652 115326 504680 235214
rect 504640 115320 504692 115326
rect 504640 115262 504692 115268
rect 504546 106040 504602 106049
rect 504546 105975 504602 105984
rect 504456 86284 504508 86290
rect 504456 86226 504508 86232
rect 504744 82142 504772 256935
rect 504836 207874 504864 348599
rect 505006 292360 505062 292369
rect 505006 292295 505062 292304
rect 504914 260536 504970 260545
rect 504914 260471 504970 260480
rect 504824 207868 504876 207874
rect 504824 207810 504876 207816
rect 504822 197160 504878 197169
rect 504822 197095 504878 197104
rect 504836 196042 504864 197095
rect 504824 196036 504876 196042
rect 504824 195978 504876 195984
rect 504822 183016 504878 183025
rect 504822 182951 504878 182960
rect 504836 182238 504864 182951
rect 504824 182232 504876 182238
rect 504824 182174 504876 182180
rect 504824 181824 504876 181830
rect 504824 181766 504876 181772
rect 504732 82136 504784 82142
rect 504732 82078 504784 82084
rect 504270 80200 504326 80209
rect 504270 80135 504326 80144
rect 504284 77353 504312 80135
rect 504270 77344 504326 77353
rect 504270 77279 504326 77288
rect 504454 49056 504510 49065
rect 504454 48991 504510 49000
rect 504468 38729 504496 48991
rect 504454 38720 504510 38729
rect 504454 38655 504510 38664
rect 504180 17468 504232 17474
rect 504180 17410 504232 17416
rect 504836 17406 504864 181766
rect 504928 115394 504956 260471
rect 505020 172990 505048 292295
rect 505008 172984 505060 172990
rect 505008 172926 505060 172932
rect 505006 172680 505062 172689
rect 505006 172615 505062 172624
rect 505020 116686 505048 172615
rect 505008 116680 505060 116686
rect 505008 116622 505060 116628
rect 504916 115388 504968 115394
rect 504916 115330 504968 115336
rect 504824 17400 504876 17406
rect 504824 17342 504876 17348
rect 504088 15904 504140 15910
rect 504088 15846 504140 15852
rect 503628 4140 503680 4146
rect 503628 4082 503680 4088
rect 503076 3188 503128 3194
rect 503076 3130 503128 3136
rect 503640 480 503668 4082
rect 504824 3596 504876 3602
rect 504824 3538 504876 3544
rect 504836 480 504864 3538
rect 505112 3398 505140 581470
rect 505204 581097 505232 581567
rect 505190 581088 505246 581097
rect 505190 581023 505246 581032
rect 505190 489560 505246 489569
rect 505190 489495 505246 489504
rect 505204 17542 505232 489495
rect 505296 122534 505324 584394
rect 505376 584248 505428 584254
rect 505376 584190 505428 584196
rect 505284 122528 505336 122534
rect 505284 122470 505336 122476
rect 505388 121854 505416 584190
rect 505836 583772 505888 583778
rect 505836 583714 505888 583720
rect 505744 462392 505796 462398
rect 505744 462334 505796 462340
rect 505558 429720 505614 429729
rect 505558 429655 505614 429664
rect 505468 418260 505520 418266
rect 505468 418202 505520 418208
rect 505376 121848 505428 121854
rect 505376 121790 505428 121796
rect 505192 17536 505244 17542
rect 505192 17478 505244 17484
rect 505480 15978 505508 418202
rect 505572 37942 505600 429655
rect 505650 412040 505706 412049
rect 505650 411975 505706 411984
rect 505664 109750 505692 411975
rect 505756 120970 505784 462334
rect 505848 322930 505876 583714
rect 505928 402824 505980 402830
rect 505928 402766 505980 402772
rect 505940 358170 505968 402766
rect 506018 366344 506074 366353
rect 506018 366279 506074 366288
rect 506032 358306 506060 366279
rect 506032 358278 506152 358306
rect 505940 358142 506060 358170
rect 505928 358080 505980 358086
rect 505928 358022 505980 358028
rect 505940 339726 505968 358022
rect 505928 339720 505980 339726
rect 505928 339662 505980 339668
rect 505836 322924 505888 322930
rect 505836 322866 505888 322872
rect 506032 321858 506060 358142
rect 506124 358086 506152 358278
rect 506112 358080 506164 358086
rect 506112 358022 506164 358028
rect 506204 339720 506256 339726
rect 506204 339662 506256 339668
rect 506216 331242 506244 339662
rect 506216 331214 506336 331242
rect 505848 321830 506060 321858
rect 505848 254862 505876 321830
rect 506308 318850 506336 331214
rect 506020 318844 506072 318850
rect 506020 318786 506072 318792
rect 506296 318844 506348 318850
rect 506296 318786 506348 318792
rect 506032 311930 506060 318786
rect 506032 311902 506152 311930
rect 506124 277914 506152 311902
rect 506112 277908 506164 277914
rect 506112 277850 506164 277856
rect 506296 264852 506348 264858
rect 506296 264794 506348 264800
rect 505836 254856 505888 254862
rect 505836 254798 505888 254804
rect 505834 253464 505890 253473
rect 505834 253399 505890 253408
rect 505848 224670 505876 253399
rect 506204 251320 506256 251326
rect 506204 251262 506256 251268
rect 506112 251252 506164 251258
rect 506112 251194 506164 251200
rect 505928 249824 505980 249830
rect 505928 249766 505980 249772
rect 505836 224664 505888 224670
rect 505836 224606 505888 224612
rect 505940 224126 505968 249766
rect 506018 232520 506074 232529
rect 506018 232455 506074 232464
rect 505928 224120 505980 224126
rect 505928 224062 505980 224068
rect 505928 214396 505980 214402
rect 505928 214338 505980 214344
rect 505836 212356 505888 212362
rect 505836 212298 505888 212304
rect 505848 203998 505876 212298
rect 505836 203992 505888 203998
rect 505836 203934 505888 203940
rect 505940 199646 505968 214338
rect 505928 199640 505980 199646
rect 505928 199582 505980 199588
rect 505928 190800 505980 190806
rect 505928 190742 505980 190748
rect 505834 178256 505890 178265
rect 505834 178191 505836 178200
rect 505888 178191 505890 178200
rect 505836 178162 505888 178168
rect 505836 170060 505888 170066
rect 505836 170002 505888 170008
rect 505848 162994 505876 170002
rect 505836 162988 505888 162994
rect 505836 162930 505888 162936
rect 505834 152688 505890 152697
rect 505834 152623 505890 152632
rect 505848 152590 505876 152623
rect 505836 152584 505888 152590
rect 505836 152526 505888 152532
rect 505834 152144 505890 152153
rect 505834 152079 505836 152088
rect 505888 152079 505890 152088
rect 505836 152050 505888 152056
rect 505836 151904 505888 151910
rect 505834 151872 505836 151881
rect 505888 151872 505890 151881
rect 505834 151807 505890 151816
rect 505836 151292 505888 151298
rect 505836 151234 505888 151240
rect 505848 143682 505876 151234
rect 505836 143676 505888 143682
rect 505836 143618 505888 143624
rect 505834 143440 505890 143449
rect 505834 143375 505890 143384
rect 505848 139913 505876 143375
rect 505834 139904 505890 139913
rect 505834 139839 505890 139848
rect 505836 131844 505888 131850
rect 505836 131786 505888 131792
rect 505848 126478 505876 131786
rect 505836 126472 505888 126478
rect 505836 126414 505888 126420
rect 505744 120964 505796 120970
rect 505744 120906 505796 120912
rect 505836 113212 505888 113218
rect 505836 113154 505888 113160
rect 505848 109886 505876 113154
rect 505940 112470 505968 190742
rect 505928 112464 505980 112470
rect 505928 112406 505980 112412
rect 505836 109880 505888 109886
rect 505836 109822 505888 109828
rect 505652 109744 505704 109750
rect 505652 109686 505704 109692
rect 505744 106344 505796 106350
rect 505744 106286 505796 106292
rect 505756 79694 505784 106286
rect 506032 80170 506060 232455
rect 506124 121038 506152 251194
rect 506216 218006 506244 251262
rect 506308 249830 506336 264794
rect 506296 249824 506348 249830
rect 506296 249766 506348 249772
rect 506296 224664 506348 224670
rect 506296 224606 506348 224612
rect 506204 218000 506256 218006
rect 506204 217942 506256 217948
rect 506308 212362 506336 224606
rect 506388 224120 506440 224126
rect 506388 224062 506440 224068
rect 506400 214402 506428 224062
rect 506388 214396 506440 214402
rect 506388 214338 506440 214344
rect 506296 212356 506348 212362
rect 506296 212298 506348 212304
rect 506296 212220 506348 212226
rect 506296 212162 506348 212168
rect 506204 204332 506256 204338
rect 506204 204274 506256 204280
rect 506112 121032 506164 121038
rect 506112 120974 506164 120980
rect 506216 120834 506244 204274
rect 506308 155378 506336 212162
rect 506388 203992 506440 203998
rect 506388 203934 506440 203940
rect 506400 170066 506428 203934
rect 506388 170060 506440 170066
rect 506388 170002 506440 170008
rect 506388 166728 506440 166734
rect 506388 166670 506440 166676
rect 506296 155372 506348 155378
rect 506296 155314 506348 155320
rect 506400 155258 506428 166670
rect 506308 155230 506428 155258
rect 506308 140690 506336 155230
rect 506388 155168 506440 155174
rect 506388 155110 506440 155116
rect 506296 140684 506348 140690
rect 506296 140626 506348 140632
rect 506400 132025 506428 155110
rect 506386 132016 506442 132025
rect 506386 131951 506442 131960
rect 506388 131844 506440 131850
rect 506388 131786 506440 131792
rect 506296 126472 506348 126478
rect 506296 126414 506348 126420
rect 506204 120828 506256 120834
rect 506204 120770 506256 120776
rect 506308 113218 506336 126414
rect 506296 113212 506348 113218
rect 506296 113154 506348 113160
rect 506112 109880 506164 109886
rect 506112 109822 506164 109828
rect 506020 80164 506072 80170
rect 506020 80106 506072 80112
rect 506020 80028 506072 80034
rect 506020 79970 506072 79976
rect 505744 79688 505796 79694
rect 505744 79630 505796 79636
rect 505928 78056 505980 78062
rect 505928 77998 505980 78004
rect 505940 63578 505968 77998
rect 505836 63572 505888 63578
rect 505836 63514 505888 63520
rect 505928 63572 505980 63578
rect 505928 63514 505980 63520
rect 505848 60790 505876 63514
rect 505836 60784 505888 60790
rect 505836 60726 505888 60732
rect 505928 60648 505980 60654
rect 505928 60590 505980 60596
rect 505940 46918 505968 60590
rect 505928 46912 505980 46918
rect 505928 46854 505980 46860
rect 505928 41268 505980 41274
rect 505928 41210 505980 41216
rect 505940 38622 505968 41210
rect 505836 38616 505888 38622
rect 505836 38558 505888 38564
rect 505928 38616 505980 38622
rect 505928 38558 505980 38564
rect 505560 37936 505612 37942
rect 505560 37878 505612 37884
rect 505848 29714 505876 38558
rect 505836 29708 505888 29714
rect 505836 29650 505888 29656
rect 505744 19236 505796 19242
rect 505744 19178 505796 19184
rect 505468 15972 505520 15978
rect 505468 15914 505520 15920
rect 505756 6118 505784 19178
rect 506032 17270 506060 79970
rect 506124 78062 506152 109822
rect 506112 78056 506164 78062
rect 506112 77998 506164 78004
rect 506020 17264 506072 17270
rect 506020 17206 506072 17212
rect 506020 11960 506072 11966
rect 506020 11902 506072 11908
rect 505744 6112 505796 6118
rect 505744 6054 505796 6060
rect 505100 3392 505152 3398
rect 505100 3334 505152 3340
rect 506032 480 506060 11902
rect 506400 2990 506428 131786
rect 506492 3942 506520 584802
rect 506572 584792 506624 584798
rect 506572 584734 506624 584740
rect 506584 4010 506612 584734
rect 506662 580952 506718 580961
rect 506662 580887 506718 580896
rect 506676 120630 506704 580887
rect 507030 434616 507086 434625
rect 507030 434551 507086 434560
rect 507044 425241 507072 434551
rect 507030 425232 507086 425241
rect 507030 425167 507086 425176
rect 507030 405648 507086 405657
rect 507030 405583 507086 405592
rect 507044 396137 507072 405583
rect 507030 396128 507086 396137
rect 507030 396063 507086 396072
rect 507030 394632 507086 394641
rect 507030 394567 507086 394576
rect 507044 387161 507072 394567
rect 507030 387152 507086 387161
rect 507030 387087 507086 387096
rect 506846 328400 506902 328409
rect 506846 328335 506902 328344
rect 506860 323649 506888 328335
rect 506846 323640 506902 323649
rect 506846 323575 506902 323584
rect 506756 309188 506808 309194
rect 506756 309130 506808 309136
rect 506768 122466 506796 309130
rect 507032 307148 507084 307154
rect 507032 307090 507084 307096
rect 507044 297401 507072 307090
rect 507030 297392 507086 297401
rect 507030 297327 507086 297336
rect 507030 280800 507086 280809
rect 507030 280735 507086 280744
rect 507044 270745 507072 280735
rect 507030 270736 507086 270745
rect 507030 270671 507086 270680
rect 507030 242176 507086 242185
rect 507030 242111 507086 242120
rect 507044 235385 507072 242111
rect 507030 235376 507086 235385
rect 507030 235311 507086 235320
rect 506938 218376 506994 218385
rect 506938 218311 506994 218320
rect 506846 190088 506902 190097
rect 506846 190023 506902 190032
rect 506756 122460 506808 122466
rect 506756 122402 506808 122408
rect 506860 121650 506888 190023
rect 506952 122194 506980 218311
rect 507030 204232 507086 204241
rect 507030 204167 507086 204176
rect 507044 122670 507072 204167
rect 507032 122664 507084 122670
rect 507032 122606 507084 122612
rect 506940 122188 506992 122194
rect 506940 122130 506992 122136
rect 506848 121644 506900 121650
rect 506848 121586 506900 121592
rect 507136 120698 507164 638930
rect 507216 592068 507268 592074
rect 507216 592010 507268 592016
rect 507228 121582 507256 592010
rect 508044 584996 508096 585002
rect 508044 584938 508096 584944
rect 507952 584724 508004 584730
rect 507952 584666 508004 584672
rect 507858 584080 507914 584089
rect 507858 584015 507914 584024
rect 507676 583092 507728 583098
rect 507676 583034 507728 583040
rect 507492 582480 507544 582486
rect 507492 582422 507544 582428
rect 507308 579692 507360 579698
rect 507308 579634 507360 579640
rect 507320 121718 507348 579634
rect 507400 552084 507452 552090
rect 507400 552026 507452 552032
rect 507412 124166 507440 552026
rect 507504 229090 507532 582422
rect 507584 368552 507636 368558
rect 507584 368494 507636 368500
rect 507492 229084 507544 229090
rect 507492 229026 507544 229032
rect 507492 157616 507544 157622
rect 507492 157558 507544 157564
rect 507400 124160 507452 124166
rect 507400 124102 507452 124108
rect 507308 121712 507360 121718
rect 507308 121654 507360 121660
rect 507216 121576 507268 121582
rect 507216 121518 507268 121524
rect 507308 121508 507360 121514
rect 507308 121450 507360 121456
rect 507124 120692 507176 120698
rect 507124 120634 507176 120640
rect 506664 120624 506716 120630
rect 506664 120566 506716 120572
rect 506662 119368 506718 119377
rect 506662 119303 506718 119312
rect 506572 4004 506624 4010
rect 506572 3946 506624 3952
rect 506480 3936 506532 3942
rect 506480 3878 506532 3884
rect 506388 2984 506440 2990
rect 506388 2926 506440 2932
rect 506676 610 506704 119303
rect 507320 114714 507348 121450
rect 507504 120057 507532 157558
rect 507596 120601 507624 368494
rect 507688 346390 507716 583034
rect 507768 376780 507820 376786
rect 507768 376722 507820 376728
rect 507676 346384 507728 346390
rect 507676 346326 507728 346332
rect 507674 319560 507730 319569
rect 507674 319495 507730 319504
rect 507688 318889 507716 319495
rect 507674 318880 507730 318889
rect 507674 318815 507730 318824
rect 507674 316024 507730 316033
rect 507674 315959 507730 315968
rect 507688 307154 507716 315959
rect 507676 307148 507728 307154
rect 507676 307090 507728 307096
rect 507674 249928 507730 249937
rect 507674 249863 507730 249872
rect 507582 120592 507638 120601
rect 507582 120527 507638 120536
rect 507490 120048 507546 120057
rect 507490 119983 507546 119992
rect 507308 114708 507360 114714
rect 507308 114650 507360 114656
rect 506940 111852 506992 111858
rect 506940 111794 506992 111800
rect 506952 102202 506980 111794
rect 506940 102196 506992 102202
rect 506940 102138 506992 102144
rect 507688 4146 507716 249863
rect 507780 158710 507808 376722
rect 507768 158704 507820 158710
rect 507768 158646 507820 158652
rect 507766 158128 507822 158137
rect 507766 158063 507822 158072
rect 507780 143857 507808 158063
rect 507766 143848 507822 143857
rect 507766 143783 507822 143792
rect 507768 140684 507820 140690
rect 507768 140626 507820 140632
rect 507780 6730 507808 140626
rect 507768 6724 507820 6730
rect 507768 6666 507820 6672
rect 507676 4140 507728 4146
rect 507676 4082 507728 4088
rect 507872 2825 507900 584015
rect 507964 3194 507992 584666
rect 507952 3188 508004 3194
rect 507952 3130 508004 3136
rect 508056 3126 508084 584938
rect 508148 119950 508176 700742
rect 508412 700460 508464 700466
rect 508412 700402 508464 700408
rect 508320 584656 508372 584662
rect 508320 584598 508372 584604
rect 508228 581800 508280 581806
rect 508228 581742 508280 581748
rect 508136 119944 508188 119950
rect 508136 119886 508188 119892
rect 508136 111444 508188 111450
rect 508136 111386 508188 111392
rect 508148 106350 508176 111386
rect 508136 106344 508188 106350
rect 508136 106286 508188 106292
rect 508044 3120 508096 3126
rect 508044 3062 508096 3068
rect 508240 2854 508268 581742
rect 508332 6050 508360 584598
rect 508424 121553 508452 700402
rect 508780 685908 508832 685914
rect 508780 685850 508832 685856
rect 508502 580680 508558 580689
rect 508502 580615 508558 580624
rect 508410 121544 508466 121553
rect 508410 121479 508466 121488
rect 508516 120358 508544 580615
rect 508596 549364 508648 549370
rect 508596 549306 508648 549312
rect 508608 121009 508636 549306
rect 508688 390584 508740 390590
rect 508688 390526 508740 390532
rect 508594 121000 508650 121009
rect 508594 120935 508650 120944
rect 508504 120352 508556 120358
rect 508504 120294 508556 120300
rect 508700 8294 508728 390526
rect 508792 362846 508820 685850
rect 509884 585132 509936 585138
rect 509884 585074 509936 585080
rect 509238 584216 509294 584225
rect 509238 584151 509294 584160
rect 508780 362840 508832 362846
rect 508780 362782 508832 362788
rect 508780 351960 508832 351966
rect 508780 351902 508832 351908
rect 508792 122262 508820 351902
rect 509056 277840 509108 277846
rect 509056 277782 509108 277788
rect 508872 236020 508924 236026
rect 508872 235962 508924 235968
rect 508780 122256 508832 122262
rect 508780 122198 508832 122204
rect 508884 119785 508912 235962
rect 508964 221876 509016 221882
rect 508964 221818 509016 221824
rect 508870 119776 508926 119785
rect 508870 119711 508926 119720
rect 508976 109002 509004 221818
rect 509068 218006 509096 277782
rect 509056 218000 509108 218006
rect 509056 217942 509108 217948
rect 509054 214840 509110 214849
rect 509054 214775 509110 214784
rect 509068 122330 509096 214775
rect 509148 196036 509200 196042
rect 509148 195978 509200 195984
rect 509056 122324 509108 122330
rect 509056 122266 509108 122272
rect 509160 119542 509188 195978
rect 509148 119536 509200 119542
rect 509148 119478 509200 119484
rect 508964 108996 509016 109002
rect 508964 108938 509016 108944
rect 508688 8288 508740 8294
rect 508688 8230 508740 8236
rect 508320 6044 508372 6050
rect 508320 5986 508372 5992
rect 508412 4140 508464 4146
rect 508412 4082 508464 4088
rect 508228 2848 508280 2854
rect 507858 2816 507914 2825
rect 508228 2790 508280 2796
rect 507858 2751 507914 2760
rect 506664 604 506716 610
rect 506664 546 506716 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 4082
rect 509252 3058 509280 584151
rect 509792 583976 509844 583982
rect 509792 583918 509844 583924
rect 509424 583908 509476 583914
rect 509424 583850 509476 583856
rect 509332 582140 509384 582146
rect 509332 582082 509384 582088
rect 509344 4078 509372 582082
rect 509436 6390 509464 583850
rect 509516 583432 509568 583438
rect 509516 583374 509568 583380
rect 509528 6662 509556 583374
rect 509700 583160 509752 583166
rect 509700 583102 509752 583108
rect 509608 582072 509660 582078
rect 509608 582014 509660 582020
rect 509620 118998 509648 582014
rect 509712 120562 509740 583102
rect 509804 121825 509832 583918
rect 509896 122126 509924 585074
rect 511356 585064 511408 585070
rect 511356 585006 511408 585012
rect 511264 584928 511316 584934
rect 511264 584870 511316 584876
rect 511172 584588 511224 584594
rect 511172 584530 511224 584536
rect 510804 584384 510856 584390
rect 510804 584326 510856 584332
rect 510068 583024 510120 583030
rect 510068 582966 510120 582972
rect 509974 581632 510030 581641
rect 509974 581567 510030 581576
rect 509988 581233 510016 581567
rect 509974 581224 510030 581233
rect 509974 581159 510030 581168
rect 509974 580272 510030 580281
rect 509974 580207 510030 580216
rect 509884 122120 509936 122126
rect 509884 122062 509936 122068
rect 509790 121816 509846 121825
rect 509790 121751 509846 121760
rect 509884 121440 509936 121446
rect 509884 121382 509936 121388
rect 509700 120556 509752 120562
rect 509700 120498 509752 120504
rect 509608 118992 509660 118998
rect 509608 118934 509660 118940
rect 509608 116000 509660 116006
rect 509608 115942 509660 115948
rect 509620 111858 509648 115942
rect 509608 111852 509660 111858
rect 509608 111794 509660 111800
rect 509896 111450 509924 121382
rect 509988 119610 510016 580207
rect 510080 171086 510108 582966
rect 510712 582344 510764 582350
rect 510712 582286 510764 582292
rect 510620 581868 510672 581874
rect 510620 581810 510672 581816
rect 510160 527196 510212 527202
rect 510160 527138 510212 527144
rect 510068 171080 510120 171086
rect 510068 171022 510120 171028
rect 510172 122806 510200 527138
rect 510252 492720 510304 492726
rect 510252 492662 510304 492668
rect 510160 122800 510212 122806
rect 510160 122742 510212 122748
rect 509976 119604 510028 119610
rect 509976 119546 510028 119552
rect 510264 119105 510292 492662
rect 510344 454096 510396 454102
rect 510344 454038 510396 454044
rect 510356 119474 510384 454038
rect 510434 246392 510490 246401
rect 510434 246327 510490 246336
rect 510448 120426 510476 246327
rect 510528 192636 510580 192642
rect 510528 192578 510580 192584
rect 510540 121514 510568 192578
rect 510528 121508 510580 121514
rect 510528 121450 510580 121456
rect 510436 120420 510488 120426
rect 510436 120362 510488 120368
rect 510344 119468 510396 119474
rect 510344 119410 510396 119416
rect 510250 119096 510306 119105
rect 510250 119031 510306 119040
rect 509884 111444 509936 111450
rect 509884 111386 509936 111392
rect 509608 11756 509660 11762
rect 509608 11698 509660 11704
rect 509516 6656 509568 6662
rect 509516 6598 509568 6604
rect 509424 6384 509476 6390
rect 509424 6326 509476 6332
rect 509332 4072 509384 4078
rect 509332 4014 509384 4020
rect 509240 3052 509292 3058
rect 509240 2994 509292 3000
rect 509620 480 509648 11698
rect 510632 2922 510660 581810
rect 510724 3262 510752 582286
rect 510816 6322 510844 584326
rect 510988 583364 511040 583370
rect 510988 583306 511040 583312
rect 510896 582956 510948 582962
rect 510896 582898 510948 582904
rect 510908 6866 510936 582898
rect 510896 6860 510948 6866
rect 510896 6802 510948 6808
rect 511000 6594 511028 583306
rect 511080 582276 511132 582282
rect 511080 582218 511132 582224
rect 511092 6798 511120 582218
rect 511184 116822 511212 584530
rect 511172 116816 511224 116822
rect 511172 116758 511224 116764
rect 511080 6792 511132 6798
rect 511080 6734 511132 6740
rect 510988 6588 511040 6594
rect 510988 6530 511040 6536
rect 510804 6316 510856 6322
rect 510804 6258 510856 6264
rect 511276 4146 511304 584870
rect 511368 119921 511396 585006
rect 524420 584520 524472 584526
rect 517518 584488 517574 584497
rect 524420 584462 524472 584468
rect 517518 584423 517574 584432
rect 511540 584044 511592 584050
rect 511540 583986 511592 583992
rect 511446 580136 511502 580145
rect 511446 580071 511502 580080
rect 511354 119912 511410 119921
rect 511354 119847 511410 119856
rect 511460 116006 511488 580071
rect 511552 121990 511580 583986
rect 514024 582616 514076 582622
rect 514024 582558 514076 582564
rect 511724 565888 511776 565894
rect 511724 565830 511776 565836
rect 511632 485784 511684 485790
rect 511632 485726 511684 485732
rect 511540 121984 511592 121990
rect 511540 121926 511592 121932
rect 511644 121446 511672 485726
rect 511736 299470 511764 565830
rect 513380 478916 513432 478922
rect 513380 478858 513432 478864
rect 511816 369912 511868 369918
rect 511816 369854 511868 369860
rect 511724 299464 511776 299470
rect 511724 299406 511776 299412
rect 511632 121440 511684 121446
rect 511632 121382 511684 121388
rect 511828 121106 511856 369854
rect 511908 340944 511960 340950
rect 511908 340886 511960 340892
rect 511816 121100 511868 121106
rect 511816 121042 511868 121048
rect 511920 120902 511948 340886
rect 511908 120896 511960 120902
rect 511908 120838 511960 120844
rect 511448 116000 511500 116006
rect 511448 115942 511500 115948
rect 511632 115864 511684 115870
rect 511632 115806 511684 115812
rect 511644 114510 511672 115806
rect 511632 114504 511684 114510
rect 511632 114446 511684 114452
rect 511540 104916 511592 104922
rect 511540 104858 511592 104864
rect 511552 104802 511580 104858
rect 511552 104786 511672 104802
rect 511552 104780 511684 104786
rect 511552 104774 511632 104780
rect 511632 104722 511684 104728
rect 511724 96552 511776 96558
rect 511724 96494 511776 96500
rect 511736 87038 511764 96494
rect 511632 87032 511684 87038
rect 511552 86980 511632 86986
rect 511552 86974 511684 86980
rect 511724 87032 511776 87038
rect 511724 86974 511776 86980
rect 511552 86958 511672 86974
rect 511552 85542 511580 86958
rect 511540 85536 511592 85542
rect 511540 85478 511592 85484
rect 511540 75948 511592 75954
rect 511540 75890 511592 75896
rect 511552 66230 511580 75890
rect 511540 66224 511592 66230
rect 511540 66166 511592 66172
rect 511540 56636 511592 56642
rect 511540 56578 511592 56584
rect 511552 46918 511580 56578
rect 511540 46912 511592 46918
rect 511540 46854 511592 46860
rect 511540 29096 511592 29102
rect 511540 29038 511592 29044
rect 511552 27606 511580 29038
rect 511540 27600 511592 27606
rect 511540 27542 511592 27548
rect 511540 18012 511592 18018
rect 511540 17954 511592 17960
rect 511552 12510 511580 17954
rect 511540 12504 511592 12510
rect 511540 12446 511592 12452
rect 511448 12436 511500 12442
rect 511448 12378 511500 12384
rect 511264 4140 511316 4146
rect 511264 4082 511316 4088
rect 510712 3256 510764 3262
rect 510712 3198 510764 3204
rect 510620 2916 510672 2922
rect 510620 2858 510672 2864
rect 511460 2802 511488 12378
rect 512090 11656 512146 11665
rect 512090 11591 512146 11600
rect 512000 4140 512052 4146
rect 512000 4082 512052 4088
rect 510816 2774 511488 2802
rect 510816 480 510844 2774
rect 512012 480 512040 4082
rect 512104 610 512132 11591
rect 513392 610 513420 478858
rect 514036 416770 514064 582558
rect 514666 545456 514722 545465
rect 514666 545391 514722 545400
rect 514680 545306 514708 545391
rect 514850 545320 514906 545329
rect 514680 545278 514850 545306
rect 514850 545255 514906 545264
rect 514024 416764 514076 416770
rect 514024 416706 514076 416712
rect 514668 181144 514720 181150
rect 514666 181112 514668 181121
rect 514720 181112 514722 181121
rect 514666 181047 514722 181056
rect 514760 118040 514812 118046
rect 514760 117982 514812 117988
rect 514772 610 514800 117982
rect 516784 6180 516836 6186
rect 516784 6122 516836 6128
rect 512092 604 512144 610
rect 512092 546 512144 552
rect 513196 604 513248 610
rect 513196 546 513248 552
rect 513380 604 513432 610
rect 513380 546 513432 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514760 604 514812 610
rect 514760 546 514812 552
rect 515588 604 515640 610
rect 515588 546 515640 552
rect 513208 480 513236 546
rect 514404 480 514432 546
rect 515600 480 515628 546
rect 516796 480 516824 6122
rect 517532 626 517560 584423
rect 520278 584352 520334 584361
rect 520278 584287 520334 584296
rect 519544 485852 519596 485858
rect 519544 485794 519596 485800
rect 519556 296682 519584 485794
rect 519544 296676 519596 296682
rect 519544 296618 519596 296624
rect 519544 225004 519596 225010
rect 519544 224946 519596 224952
rect 519556 64870 519584 224946
rect 519636 119740 519688 119746
rect 519636 119682 519688 119688
rect 519544 64864 519596 64870
rect 519544 64806 519596 64812
rect 519084 9036 519136 9042
rect 519084 8978 519136 8984
rect 517532 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 8978
rect 519648 3670 519676 119682
rect 520292 7614 520320 584287
rect 523038 581360 523094 581369
rect 523038 581295 523094 581304
rect 521568 181144 521620 181150
rect 521566 181112 521568 181121
rect 521620 181112 521622 181121
rect 521566 181047 521622 181056
rect 522304 119876 522356 119882
rect 522304 119818 522356 119824
rect 520280 7608 520332 7614
rect 520280 7550 520332 7556
rect 521476 7608 521528 7614
rect 521476 7550 521528 7556
rect 520280 6520 520332 6526
rect 520280 6462 520332 6468
rect 519636 3664 519688 3670
rect 519636 3606 519688 3612
rect 520292 480 520320 6462
rect 521488 480 521516 7550
rect 522316 3602 522344 119818
rect 523052 12442 523080 581295
rect 524432 570217 524460 584462
rect 524418 570208 524474 570217
rect 524418 570143 524474 570152
rect 524418 570072 524474 570081
rect 524418 570007 524474 570016
rect 524432 568546 524460 570007
rect 524420 568540 524472 568546
rect 524420 568482 524472 568488
rect 524604 550656 524656 550662
rect 524604 550598 524656 550604
rect 524326 545320 524382 545329
rect 524382 545278 524552 545306
rect 524326 545255 524382 545264
rect 524524 545193 524552 545278
rect 524510 545184 524566 545193
rect 524510 545119 524566 545128
rect 524616 543794 524644 550598
rect 524420 543788 524472 543794
rect 524420 543730 524472 543736
rect 524604 543788 524656 543794
rect 524604 543730 524656 543736
rect 524432 471986 524460 543730
rect 524420 471980 524472 471986
rect 524420 471922 524472 471928
rect 524420 462460 524472 462466
rect 524420 462402 524472 462408
rect 524432 452606 524460 462402
rect 524420 452600 524472 452606
rect 524420 452542 524472 452548
rect 524420 443012 524472 443018
rect 524420 442954 524472 442960
rect 524432 433294 524460 442954
rect 524420 433288 524472 433294
rect 524420 433230 524472 433236
rect 524420 423700 524472 423706
rect 524420 423642 524472 423648
rect 524432 413982 524460 423642
rect 524420 413976 524472 413982
rect 524420 413918 524472 413924
rect 524420 404388 524472 404394
rect 524420 404330 524472 404336
rect 524432 394670 524460 404330
rect 524420 394664 524472 394670
rect 524420 394606 524472 394612
rect 524420 385076 524472 385082
rect 524420 385018 524472 385024
rect 524432 375358 524460 385018
rect 524420 375352 524472 375358
rect 524420 375294 524472 375300
rect 524420 365764 524472 365770
rect 524420 365706 524472 365712
rect 524432 356046 524460 365706
rect 524420 356040 524472 356046
rect 524420 355982 524472 355988
rect 524420 346452 524472 346458
rect 524420 346394 524472 346400
rect 524432 336734 524460 346394
rect 524420 336728 524472 336734
rect 524420 336670 524472 336676
rect 524420 327140 524472 327146
rect 524420 327082 524472 327088
rect 524432 317422 524460 327082
rect 524420 317416 524472 317422
rect 524420 317358 524472 317364
rect 524420 307828 524472 307834
rect 524420 307770 524472 307776
rect 524432 298110 524460 307770
rect 524420 298104 524472 298110
rect 524420 298046 524472 298052
rect 524420 288448 524472 288454
rect 524420 288390 524472 288396
rect 524432 278769 524460 288390
rect 524418 278760 524474 278769
rect 524418 278695 524474 278704
rect 524602 278760 524658 278769
rect 524602 278695 524658 278704
rect 524616 269142 524644 278695
rect 524420 269136 524472 269142
rect 524420 269078 524472 269084
rect 524604 269136 524656 269142
rect 524604 269078 524656 269084
rect 524432 259457 524460 269078
rect 524418 259448 524474 259457
rect 524418 259383 524474 259392
rect 524602 259448 524658 259457
rect 524602 259383 524658 259392
rect 524616 249830 524644 259383
rect 524420 249824 524472 249830
rect 524420 249766 524472 249772
rect 524604 249824 524656 249830
rect 524604 249766 524656 249772
rect 524432 241777 524460 249766
rect 524418 241768 524474 241777
rect 524418 241703 524474 241712
rect 524418 241632 524474 241641
rect 524418 241567 524474 241576
rect 524432 240145 524460 241567
rect 524418 240136 524474 240145
rect 524418 240071 524474 240080
rect 524602 240136 524658 240145
rect 524602 240071 524658 240080
rect 524616 230518 524644 240071
rect 524420 230512 524472 230518
rect 524420 230454 524472 230460
rect 524604 230512 524656 230518
rect 524604 230454 524656 230460
rect 524432 220833 524460 230454
rect 524418 220824 524474 220833
rect 524418 220759 524474 220768
rect 524602 220824 524658 220833
rect 524602 220759 524658 220768
rect 524616 211177 524644 220759
rect 524418 211168 524474 211177
rect 524418 211103 524474 211112
rect 524602 211168 524658 211177
rect 524602 211103 524658 211112
rect 524432 201482 524460 211103
rect 524420 201476 524472 201482
rect 524420 201418 524472 201424
rect 524604 201476 524656 201482
rect 524604 201418 524656 201424
rect 524616 191865 524644 201418
rect 524418 191856 524474 191865
rect 524418 191791 524474 191800
rect 524602 191856 524658 191865
rect 524602 191791 524658 191800
rect 524432 182170 524460 191791
rect 524420 182164 524472 182170
rect 524420 182106 524472 182112
rect 524604 182164 524656 182170
rect 524604 182106 524656 182112
rect 524616 172553 524644 182106
rect 524418 172544 524474 172553
rect 524418 172479 524474 172488
rect 524602 172544 524658 172553
rect 524602 172479 524658 172488
rect 524432 162858 524460 172479
rect 527192 165578 527220 703520
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 542358 585032 542414 585041
rect 542358 584967 542414 584976
rect 534080 584112 534132 584118
rect 534080 584054 534132 584060
rect 532700 581664 532752 581670
rect 532700 581606 532752 581612
rect 532712 578241 532740 581606
rect 532698 578232 532754 578241
rect 532698 578167 532754 578176
rect 532882 578232 532938 578241
rect 532882 578167 532938 578176
rect 532896 568614 532924 578167
rect 532700 568608 532752 568614
rect 532422 568576 532478 568585
rect 532422 568511 532478 568520
rect 532698 568576 532700 568585
rect 532884 568608 532936 568614
rect 532752 568576 532754 568585
rect 532884 568550 532936 568556
rect 532698 568511 532754 568520
rect 532436 558958 532464 568511
rect 532424 558952 532476 558958
rect 532424 558894 532476 558900
rect 532516 558952 532568 558958
rect 532516 558894 532568 558900
rect 529204 556232 529256 556238
rect 529204 556174 529256 556180
rect 529216 324290 529244 556174
rect 532528 553314 532556 558894
rect 532516 553308 532568 553314
rect 532516 553250 532568 553256
rect 532884 553308 532936 553314
rect 532884 553250 532936 553256
rect 532896 550610 532924 553250
rect 532896 550582 533016 550610
rect 531962 545456 532018 545465
rect 531962 545391 532018 545400
rect 531976 545222 532004 545391
rect 529940 545216 529992 545222
rect 529938 545184 529940 545193
rect 531964 545216 532016 545222
rect 529992 545184 529994 545193
rect 531964 545158 532016 545164
rect 529938 545119 529994 545128
rect 532988 541006 533016 550582
rect 532700 541000 532752 541006
rect 532700 540942 532752 540948
rect 532976 541000 533028 541006
rect 532976 540942 533028 540948
rect 532712 531321 532740 540942
rect 532698 531312 532754 531321
rect 532698 531247 532754 531256
rect 532882 531312 532938 531321
rect 532882 531247 532938 531256
rect 532896 521694 532924 531247
rect 532700 521688 532752 521694
rect 532700 521630 532752 521636
rect 532884 521688 532936 521694
rect 532884 521630 532936 521636
rect 532712 512009 532740 521630
rect 532698 512000 532754 512009
rect 532698 511935 532754 511944
rect 532882 512000 532938 512009
rect 532882 511935 532938 511944
rect 532896 502382 532924 511935
rect 532700 502376 532752 502382
rect 532700 502318 532752 502324
rect 532884 502376 532936 502382
rect 532884 502318 532936 502324
rect 532712 492658 532740 502318
rect 532700 492652 532752 492658
rect 532700 492594 532752 492600
rect 532884 492652 532936 492658
rect 532884 492594 532936 492600
rect 532896 483041 532924 492594
rect 532698 483032 532754 483041
rect 532698 482967 532754 482976
rect 532882 483032 532938 483041
rect 532882 482967 532938 482976
rect 531964 470620 532016 470626
rect 531964 470562 532016 470568
rect 529204 324284 529256 324290
rect 529204 324226 529256 324232
rect 529938 238912 529994 238921
rect 529938 238847 529940 238856
rect 529992 238847 529994 238856
rect 529940 238818 529992 238824
rect 527180 165572 527232 165578
rect 527180 165514 527232 165520
rect 524420 162852 524472 162858
rect 524420 162794 524472 162800
rect 524420 153264 524472 153270
rect 524420 153206 524472 153212
rect 524432 143546 524460 153206
rect 524420 143540 524472 143546
rect 524420 143482 524472 143488
rect 524420 133952 524472 133958
rect 524420 133894 524472 133900
rect 524432 124098 524460 133894
rect 524420 124092 524472 124098
rect 524420 124034 524472 124040
rect 529938 116648 529994 116657
rect 529938 116583 529994 116592
rect 524420 114572 524472 114578
rect 524420 114514 524472 114520
rect 524432 104854 524460 114514
rect 524420 104848 524472 104854
rect 524420 104790 524472 104796
rect 524420 95260 524472 95266
rect 524420 95202 524472 95208
rect 524432 85542 524460 95202
rect 524420 85536 524472 85542
rect 524420 85478 524472 85484
rect 524420 75948 524472 75954
rect 524420 75890 524472 75896
rect 524432 66230 524460 75890
rect 524420 66224 524472 66230
rect 524420 66166 524472 66172
rect 524420 56636 524472 56642
rect 524420 56578 524472 56584
rect 524432 46918 524460 56578
rect 524420 46912 524472 46918
rect 524420 46854 524472 46860
rect 524420 37324 524472 37330
rect 524420 37266 524472 37272
rect 524432 27606 524460 37266
rect 524420 27600 524472 27606
rect 524420 27542 524472 27548
rect 524420 18012 524472 18018
rect 524420 17954 524472 17960
rect 524432 12510 524460 17954
rect 524420 12504 524472 12510
rect 524420 12446 524472 12452
rect 529952 12442 529980 116583
rect 523040 12436 523092 12442
rect 523040 12378 523092 12384
rect 523868 12436 523920 12442
rect 523868 12378 523920 12384
rect 529940 12436 529992 12442
rect 529940 12378 529992 12384
rect 531044 12436 531096 12442
rect 531044 12378 531096 12384
rect 522672 4820 522724 4826
rect 522672 4762 522724 4768
rect 522304 3596 522356 3602
rect 522304 3538 522356 3544
rect 522684 480 522712 4762
rect 523880 480 523908 12378
rect 525064 12368 525116 12374
rect 525064 12310 525116 12316
rect 527456 12368 527508 12374
rect 527456 12310 527508 12316
rect 525076 9654 525104 12310
rect 527468 9654 527496 12310
rect 525064 9648 525116 9654
rect 525064 9590 525116 9596
rect 527456 9648 527508 9654
rect 527456 9590 527508 9596
rect 525064 9512 525116 9518
rect 525064 9454 525116 9460
rect 527456 9512 527508 9518
rect 527456 9454 527508 9460
rect 525076 480 525104 9454
rect 526260 9172 526312 9178
rect 526260 9114 526312 9120
rect 526272 480 526300 9114
rect 527468 480 527496 9454
rect 529848 7676 529900 7682
rect 529848 7618 529900 7624
rect 528652 3664 528704 3670
rect 528652 3606 528704 3612
rect 528664 480 528692 3606
rect 529860 480 529888 7618
rect 531056 480 531084 12378
rect 531976 3670 532004 470562
rect 532712 183569 532740 482967
rect 532698 183560 532754 183569
rect 532698 183495 532754 183504
rect 532882 183560 532938 183569
rect 532882 183495 532938 183504
rect 532896 172553 532924 183495
rect 533988 181008 534040 181014
rect 533986 180976 533988 180985
rect 534040 180976 534042 180985
rect 533986 180911 534042 180920
rect 532698 172544 532754 172553
rect 532698 172479 532754 172488
rect 532882 172544 532938 172553
rect 532882 172479 532938 172488
rect 532712 162858 532740 172479
rect 532700 162852 532752 162858
rect 532700 162794 532752 162800
rect 532700 153264 532752 153270
rect 532700 153206 532752 153212
rect 532712 143546 532740 153206
rect 532700 143540 532752 143546
rect 532700 143482 532752 143488
rect 532700 133952 532752 133958
rect 532700 133894 532752 133900
rect 532712 124098 532740 133894
rect 532700 124092 532752 124098
rect 532700 124034 532752 124040
rect 532700 114572 532752 114578
rect 532700 114514 532752 114520
rect 532712 104854 532740 114514
rect 532700 104848 532752 104854
rect 532700 104790 532752 104796
rect 532700 95260 532752 95266
rect 532700 95202 532752 95208
rect 532712 85542 532740 95202
rect 532700 85536 532752 85542
rect 532700 85478 532752 85484
rect 532700 75948 532752 75954
rect 532700 75890 532752 75896
rect 532712 66230 532740 75890
rect 532700 66224 532752 66230
rect 532700 66166 532752 66172
rect 532700 56636 532752 56642
rect 532700 56578 532752 56584
rect 532712 46918 532740 56578
rect 532700 46912 532752 46918
rect 532700 46854 532752 46860
rect 532700 37324 532752 37330
rect 532700 37266 532752 37272
rect 532712 27606 532740 37266
rect 532700 27600 532752 27606
rect 532700 27542 532752 27548
rect 534092 12442 534120 584054
rect 536840 556300 536892 556306
rect 536840 556242 536892 556248
rect 535460 181008 535512 181014
rect 535458 180976 535460 180985
rect 535512 180976 535514 180985
rect 535458 180911 535514 180920
rect 534080 12436 534132 12442
rect 534080 12378 534132 12384
rect 534540 12436 534592 12442
rect 534540 12378 534592 12384
rect 533436 9716 533488 9722
rect 533436 9658 533488 9664
rect 531964 3664 532016 3670
rect 531964 3606 532016 3612
rect 532240 3596 532292 3602
rect 532240 3538 532292 3544
rect 532252 480 532280 3538
rect 533448 480 533476 9658
rect 534552 480 534580 12378
rect 536852 7614 536880 556242
rect 540244 372632 540296 372638
rect 540244 372574 540296 372580
rect 538864 329860 538916 329866
rect 538864 329802 538916 329808
rect 536932 117972 536984 117978
rect 536932 117914 536984 117920
rect 536840 7608 536892 7614
rect 536840 7550 536892 7556
rect 535734 6352 535790 6361
rect 535734 6287 535790 6296
rect 535748 480 535776 6287
rect 536944 480 536972 117914
rect 538218 13016 538274 13025
rect 538218 12951 538274 12960
rect 538232 12442 538260 12951
rect 538220 12436 538272 12442
rect 538220 12378 538272 12384
rect 538128 7608 538180 7614
rect 538128 7550 538180 7556
rect 538140 480 538168 7550
rect 538876 3806 538904 329802
rect 539508 239012 539560 239018
rect 539508 238954 539560 238960
rect 539520 238921 539548 238954
rect 539506 238912 539562 238921
rect 539506 238847 539562 238856
rect 540256 41410 540284 372574
rect 540334 119504 540390 119513
rect 540334 119439 540390 119448
rect 540244 41404 540296 41410
rect 540244 41346 540296 41352
rect 539324 12436 539376 12442
rect 539324 12378 539376 12384
rect 538864 3800 538916 3806
rect 538864 3742 538916 3748
rect 539336 480 539364 12378
rect 540348 3670 540376 119439
rect 542372 12442 542400 584967
rect 546498 584624 546554 584633
rect 546498 584559 546554 584568
rect 543740 581936 543792 581942
rect 543740 581878 543792 581884
rect 542360 12436 542412 12442
rect 542360 12378 542412 12384
rect 542912 12436 542964 12442
rect 542912 12378 542964 12384
rect 541716 9716 541768 9722
rect 541716 9658 541768 9664
rect 540520 9104 540572 9110
rect 540520 9046 540572 9052
rect 540336 3664 540388 3670
rect 540336 3606 540388 3612
rect 540532 480 540560 9046
rect 541728 480 541756 9658
rect 542924 480 542952 12378
rect 543752 3482 543780 581878
rect 545120 274712 545172 274718
rect 545120 274654 545172 274660
rect 545132 3482 545160 274654
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 480 546540 584559
rect 556160 584180 556212 584186
rect 556160 584122 556212 584128
rect 554872 581732 554924 581738
rect 554872 581674 554924 581680
rect 549260 239012 549312 239018
rect 549260 238954 549312 238960
rect 546592 10600 546644 10606
rect 546592 10542 546644 10548
rect 546604 3482 546632 10542
rect 548892 3800 548944 3806
rect 548892 3742 548944 3748
rect 546604 3454 547736 3482
rect 547708 480 547736 3454
rect 548904 480 548932 3742
rect 549272 3482 549300 238954
rect 552020 115252 552072 115258
rect 552020 115194 552072 115200
rect 551192 8968 551244 8974
rect 551192 8910 551244 8916
rect 549272 3454 550128 3482
rect 550100 480 550128 3454
rect 551204 480 551232 8910
rect 552032 3482 552060 115194
rect 553398 14512 553454 14521
rect 553398 14447 553454 14456
rect 553412 3482 553440 14447
rect 554780 3528 554832 3534
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 554780 3470 554832 3476
rect 554884 3482 554912 581674
rect 556172 3482 556200 584122
rect 580262 583944 580318 583953
rect 580262 583879 580318 583888
rect 560944 582752 560996 582758
rect 560944 582694 560996 582700
rect 558918 581088 558974 581097
rect 558918 581023 558974 581032
rect 558366 3768 558422 3777
rect 558366 3703 558422 3712
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 3470
rect 554884 3454 556016 3482
rect 556172 3454 557212 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3454
rect 558380 480 558408 3703
rect 558932 3482 558960 581023
rect 560956 276010 560984 582694
rect 579618 582176 579674 582185
rect 579618 582111 579674 582120
rect 569960 581596 570012 581602
rect 569960 581538 570012 581544
rect 564440 306400 564492 306406
rect 564440 306342 564492 306348
rect 560944 276004 560996 276010
rect 560944 275946 560996 275952
rect 563060 147688 563112 147694
rect 563060 147630 563112 147636
rect 560298 15872 560354 15881
rect 560298 15807 560354 15816
rect 560312 3482 560340 15807
rect 561954 6216 562010 6225
rect 561954 6151 562010 6160
rect 558932 3454 559604 3482
rect 560312 3454 560800 3482
rect 559576 480 559604 3454
rect 560772 480 560800 3454
rect 561968 480 561996 6151
rect 563072 2786 563100 147630
rect 563150 116512 563206 116521
rect 563150 116447 563206 116456
rect 563060 2780 563112 2786
rect 563060 2722 563112 2728
rect 563164 480 563192 116447
rect 564452 3482 564480 306342
rect 565820 13116 565872 13122
rect 565820 13058 565872 13064
rect 565832 3482 565860 13058
rect 567844 3732 567896 3738
rect 567844 3674 567896 3680
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 564348 2780 564400 2786
rect 564348 2722 564400 2728
rect 564360 480 564388 2722
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3674
rect 569040 3460 569092 3466
rect 569040 3402 569092 3408
rect 569052 480 569080 3402
rect 569972 3346 570000 581538
rect 574100 563100 574152 563106
rect 574100 563042 574152 563048
rect 572720 207052 572772 207058
rect 572720 206994 572772 207000
rect 571984 182232 572036 182238
rect 571984 182174 572036 182180
rect 571340 119400 571392 119406
rect 571340 119342 571392 119348
rect 571352 3482 571380 119342
rect 571432 10464 571484 10470
rect 571432 10406 571484 10412
rect 571444 3602 571472 10406
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 571352 3454 571472 3482
rect 569972 3318 570276 3346
rect 570248 480 570276 3318
rect 571444 480 571472 3454
rect 571996 2922 572024 182174
rect 572628 3596 572680 3602
rect 572628 3538 572680 3544
rect 571984 2916 572036 2922
rect 571984 2858 572036 2864
rect 572640 480 572668 3538
rect 572732 3346 572760 206994
rect 574112 3346 574140 563042
rect 576860 13252 576912 13258
rect 576860 13194 576912 13200
rect 576216 3460 576268 3466
rect 576216 3402 576268 3408
rect 572732 3318 573864 3346
rect 574112 3318 575060 3346
rect 573836 480 573864 3318
rect 575032 480 575060 3318
rect 576228 480 576256 3402
rect 576872 610 576900 13194
rect 578608 2916 578660 2922
rect 578608 2858 578660 2864
rect 576860 604 576912 610
rect 576860 546 576912 552
rect 577412 604 577464 610
rect 577412 546 577464 552
rect 577424 480 577452 546
rect 578620 480 578648 2858
rect 579632 610 579660 582111
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580172 534064 580224 534070
rect 580172 534006 580224 534012
rect 580184 533905 580212 534006
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580172 510604 580224 510610
rect 580172 510546 580224 510552
rect 580184 510377 580212 510546
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 579988 499520 580040 499526
rect 579988 499462 580040 499468
rect 580000 498681 580028 499462
rect 579986 498672 580042 498681
rect 579986 498607 580042 498616
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 579988 440224 580040 440230
rect 579988 440166 580040 440172
rect 580000 439929 580028 440166
rect 579986 439920 580042 439929
rect 579986 439855 580042 439864
rect 580172 416764 580224 416770
rect 580172 416706 580224 416712
rect 580184 416537 580212 416706
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 579712 393304 579764 393310
rect 579712 393246 579764 393252
rect 579724 393009 579752 393246
rect 579710 393000 579766 393009
rect 579710 392935 579766 392944
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 580172 346384 580224 346390
rect 580172 346326 580224 346332
rect 580184 346089 580212 346326
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 251258 580212 252175
rect 580172 251252 580224 251258
rect 580172 251194 580224 251200
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580184 204338 580212 205255
rect 580172 204332 580224 204338
rect 580172 204274 580224 204280
rect 579710 181928 579766 181937
rect 579710 181863 579766 181872
rect 579724 181121 579752 181863
rect 579710 181112 579766 181121
rect 579710 181047 579766 181056
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 580172 158704 580224 158710
rect 580172 158646 580224 158652
rect 580184 158409 580212 158646
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580276 17649 580304 583879
rect 580540 581460 580592 581466
rect 580540 581402 580592 581408
rect 580356 581324 580408 581330
rect 580356 581266 580408 581272
rect 580368 111489 580396 581266
rect 580448 581256 580500 581262
rect 580448 581198 580500 581204
rect 580460 451761 580488 581198
rect 580446 451752 580502 451761
rect 580446 451687 580502 451696
rect 580446 404832 580502 404841
rect 580446 404767 580502 404776
rect 580460 120766 580488 404767
rect 580552 310865 580580 581402
rect 580630 357912 580686 357921
rect 580630 357847 580686 357856
rect 580538 310856 580594 310865
rect 580538 310791 580594 310800
rect 580644 121174 580672 357847
rect 580632 121168 580684 121174
rect 580632 121110 580684 121116
rect 580448 120760 580500 120766
rect 580448 120702 580500 120708
rect 580354 111480 580410 111489
rect 580354 111415 580410 111424
rect 580262 17640 580318 17649
rect 580262 17575 580318 17584
rect 581092 10396 581144 10402
rect 581092 10338 581144 10344
rect 581104 626 581132 10338
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 579620 604 579672 610
rect 579620 546 579672 552
rect 579804 604 579856 610
rect 579804 546 579856 552
rect 581012 598 581132 626
rect 579816 480 579844 546
rect 581012 480 581040 598
rect 582208 480 582236 3606
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3146 553016 3202 553072
rect 2870 509904 2926 509960
rect 3330 481072 3386 481128
rect 2962 423680 3018 423736
rect 3330 394984 3386 395040
rect 3054 380568 3110 380624
rect 2962 337456 3018 337512
rect 3330 323040 3386 323096
rect 3330 308760 3386 308816
rect 3238 294344 3294 294400
rect 2778 280064 2834 280120
rect 2962 265648 3018 265704
rect 3330 251252 3386 251288
rect 3330 251232 3332 251252
rect 3332 251232 3384 251252
rect 3384 251232 3386 251252
rect 3238 236952 3294 237008
rect 3330 222536 3386 222592
rect 3146 208120 3202 208176
rect 2778 200232 2834 200288
rect 3514 567296 3570 567352
rect 3514 538600 3570 538656
rect 3514 495488 3570 495544
rect 3514 437960 3570 438016
rect 3422 193840 3478 193896
rect 3238 179424 3294 179480
rect 3422 165008 3478 165064
rect 3146 150728 3202 150784
rect 3422 136312 3478 136368
rect 3606 366152 3662 366208
rect 3514 122032 3570 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3422 80008 3478 80064
rect 3422 78920 3478 78976
rect 2778 64540 2780 64560
rect 2780 64540 2832 64560
rect 2832 64540 2834 64560
rect 2778 64504 2834 64540
rect 3422 50088 3478 50144
rect 3146 35844 3148 35864
rect 3148 35844 3200 35864
rect 3200 35844 3202 35864
rect 3146 35808 3202 35844
rect 3422 7112 3478 7168
rect 8758 579672 8814 579728
rect 5262 4800 5318 4856
rect 13634 101360 13690 101416
rect 16026 4936 16082 4992
rect 64694 18536 64750 18592
rect 70306 3984 70362 4040
rect 73618 340992 73674 341048
rect 74446 513712 74502 513768
rect 74354 503104 74410 503160
rect 74170 358672 74226 358728
rect 75090 436192 75146 436248
rect 75642 281152 75698 281208
rect 75458 277616 75514 277672
rect 76838 450336 76894 450392
rect 76746 418512 76802 418568
rect 76470 333940 76526 333976
rect 76470 333920 76472 333940
rect 76472 333920 76524 333940
rect 76524 333920 76526 333940
rect 76654 288224 76710 288280
rect 76010 249600 76066 249656
rect 76562 228384 76618 228440
rect 76378 201864 76434 201920
rect 76378 198056 76434 198112
rect 77574 478352 77630 478408
rect 77574 429120 77630 429176
rect 77666 407904 77722 407960
rect 77574 379888 77630 379944
rect 77574 372816 77630 372872
rect 77574 362208 77630 362264
rect 77574 344528 77630 344584
rect 77574 330384 77630 330440
rect 77666 323584 77722 323640
rect 77574 309440 77630 309496
rect 77574 295432 77630 295488
rect 77574 267008 77630 267064
rect 77482 256672 77538 256728
rect 77390 247832 77446 247888
rect 77390 237632 77446 237688
rect 78126 506640 78182 506696
rect 78034 499568 78090 499624
rect 77942 129648 77998 129704
rect 78678 573552 78734 573608
rect 78678 559408 78734 559464
rect 79966 534656 80022 534712
rect 78678 520784 78734 520840
rect 81346 562944 81402 563000
rect 81162 488960 81218 489016
rect 79874 481888 79930 481944
rect 79690 446800 79746 446856
rect 79414 411440 79470 411496
rect 78770 400832 78826 400888
rect 78770 393760 78826 393816
rect 79138 348064 79194 348120
rect 79046 253136 79102 253192
rect 78954 231920 79010 231976
rect 78862 196560 78918 196616
rect 78770 184592 78826 184648
rect 78770 182688 78826 182744
rect 78678 172080 78734 172136
rect 78678 168544 78734 168600
rect 78678 165008 78734 165064
rect 78678 161472 78734 161528
rect 78770 150864 78826 150920
rect 78770 133184 78826 133240
rect 79322 274080 79378 274136
rect 79230 259936 79286 259992
rect 79138 202952 79194 203008
rect 79506 284688 79562 284744
rect 79414 210704 79470 210760
rect 79598 130464 79654 130520
rect 79598 123256 79654 123312
rect 79782 351600 79838 351656
rect 80978 471280 81034 471336
rect 80886 460672 80942 460728
rect 80794 443264 80850 443320
rect 80702 439728 80758 439784
rect 80610 404368 80666 404424
rect 79966 337456 80022 337512
rect 80518 316512 80574 316568
rect 79966 175616 80022 175672
rect 79966 154400 80022 154456
rect 79874 126112 79930 126168
rect 79966 123120 80022 123176
rect 80426 241440 80482 241496
rect 80426 239400 80482 239456
rect 80334 236952 80390 237008
rect 80334 236136 80390 236192
rect 80334 217776 80390 217832
rect 80150 209072 80206 209128
rect 80242 207712 80298 207768
rect 80150 202680 80206 202736
rect 80150 202000 80206 202056
rect 80334 203632 80390 203688
rect 80426 202952 80482 203008
rect 80242 201592 80298 201648
rect 80150 199552 80206 199608
rect 80150 190304 80206 190360
rect 80334 188400 80390 188456
rect 80334 186224 80390 186280
rect 80242 179968 80298 180024
rect 80242 179832 80298 179888
rect 80150 178336 80206 178392
rect 80150 171400 80206 171456
rect 80242 171128 80298 171184
rect 80150 165552 80206 165608
rect 80150 149640 80206 149696
rect 80242 144084 80298 144120
rect 80242 144064 80244 144084
rect 80244 144064 80296 144084
rect 80296 144064 80298 144084
rect 80242 143792 80298 143848
rect 80150 143112 80206 143168
rect 80150 141888 80206 141944
rect 80150 140256 80206 140312
rect 80150 123392 80206 123448
rect 80426 137264 80482 137320
rect 80426 137164 80428 137184
rect 80428 137164 80480 137184
rect 80480 137164 80482 137184
rect 80426 137128 80482 137164
rect 80426 136856 80482 136912
rect 80426 136720 80482 136776
rect 80426 135904 80482 135960
rect 80058 6840 80114 6896
rect 80334 6840 80390 6896
rect 79046 3712 79102 3768
rect 81070 464208 81126 464264
rect 80978 136720 81034 136776
rect 81254 425584 81310 425640
rect 81438 238992 81494 239048
rect 81438 233708 81494 233744
rect 81438 233688 81440 233708
rect 81440 233688 81492 233708
rect 81492 233688 81494 233708
rect 81438 229472 81494 229528
rect 81438 229236 81440 229256
rect 81440 229236 81492 229256
rect 81492 229236 81494 229256
rect 81438 229200 81494 229236
rect 81438 227876 81440 227896
rect 81440 227876 81492 227896
rect 81492 227876 81494 227896
rect 81438 227840 81494 227876
rect 81438 223352 81494 223408
rect 81622 566480 81678 566536
rect 81530 221312 81586 221368
rect 81530 214240 81586 214296
rect 81530 210432 81586 210488
rect 81438 207984 81494 208040
rect 81530 207168 81586 207224
rect 81530 201864 81586 201920
rect 81530 201220 81532 201240
rect 81532 201220 81584 201240
rect 81584 201220 81586 201240
rect 81530 201184 81586 201220
rect 81530 201048 81586 201104
rect 81438 200096 81494 200152
rect 81530 192228 81586 192264
rect 81530 192208 81532 192228
rect 81532 192208 81584 192228
rect 81584 192208 81586 192228
rect 81530 191820 81586 191856
rect 81530 191800 81532 191820
rect 81532 191800 81584 191820
rect 81584 191800 81586 191820
rect 81530 170720 81586 170776
rect 81530 162172 81586 162208
rect 81530 162152 81532 162172
rect 81532 162152 81584 162172
rect 81584 162152 81586 162172
rect 81530 160792 81586 160848
rect 81530 157292 81532 157312
rect 81532 157292 81584 157312
rect 81584 157292 81586 157312
rect 81530 157256 81586 157292
rect 81530 144064 81586 144120
rect 81530 143928 81586 143984
rect 81806 517248 81862 517304
rect 81714 414976 81770 415032
rect 154118 700712 154174 700768
rect 218978 700576 219034 700632
rect 267646 700440 267702 700496
rect 89166 699760 89222 699816
rect 89534 695408 89590 695464
rect 89534 689288 89590 689344
rect 89534 674736 89590 674792
rect 89534 665216 89590 665272
rect 89534 655424 89590 655480
rect 89534 645904 89590 645960
rect 89534 636112 89590 636168
rect 89534 626592 89590 626648
rect 81990 467200 82046 467256
rect 81898 327392 81954 327448
rect 81898 291216 81954 291272
rect 83554 597488 83610 597544
rect 83738 597488 83794 597544
rect 89442 596128 89498 596184
rect 82634 577632 82690 577688
rect 89350 582800 89406 582856
rect 89074 582256 89130 582312
rect 86314 581712 86370 581768
rect 89718 582020 89720 582040
rect 89720 582020 89772 582040
rect 89772 582020 89774 582040
rect 89718 581984 89774 582020
rect 89810 581848 89866 581904
rect 89074 581576 89130 581632
rect 89810 581576 89866 581632
rect 85210 581440 85266 581496
rect 85486 581440 85542 581496
rect 92110 583752 92166 583808
rect 93674 582256 93730 582312
rect 91926 581848 91982 581904
rect 93398 581984 93454 582040
rect 94226 582392 94282 582448
rect 94134 582256 94190 582312
rect 93766 582120 93822 582176
rect 101310 582392 101366 582448
rect 94226 581712 94282 581768
rect 96894 581712 96950 581768
rect 93766 581440 93822 581496
rect 101586 582256 101642 582312
rect 99470 581440 99526 581496
rect 99838 581440 99894 581496
rect 84934 581304 84990 581360
rect 89258 581304 89314 581360
rect 90454 581304 90510 581360
rect 90914 581304 90970 581360
rect 91742 581304 91798 581360
rect 92662 581304 92718 581360
rect 93214 581304 93270 581360
rect 93398 581304 93454 581360
rect 96894 581304 96950 581360
rect 107658 582392 107714 582448
rect 113270 582392 113326 582448
rect 111062 581576 111118 581632
rect 113270 581440 113326 581496
rect 100022 581304 100078 581360
rect 103426 581340 103428 581360
rect 103428 581340 103480 581360
rect 103480 581340 103482 581360
rect 103426 581304 103482 581340
rect 123482 582256 123538 582312
rect 123758 582276 123814 582312
rect 123758 582256 123760 582276
rect 123760 582256 123812 582276
rect 123812 582256 123814 582276
rect 118606 581984 118662 582040
rect 118514 581576 118570 581632
rect 148782 584840 148838 584896
rect 157246 584840 157302 584896
rect 157430 584840 157486 584896
rect 128358 581984 128414 582040
rect 132498 582392 132554 582448
rect 123482 581440 123538 581496
rect 132958 582256 133014 582312
rect 139214 583752 139270 583808
rect 137926 581984 137982 582040
rect 142802 582256 142858 582312
rect 147678 582256 147734 582312
rect 132590 581440 132646 581496
rect 132958 581440 133014 581496
rect 142802 581440 142858 581496
rect 147678 581984 147734 582040
rect 158350 584704 158406 584760
rect 156326 582392 156382 582448
rect 150990 582276 151046 582312
rect 150990 582256 150992 582276
rect 150992 582256 151044 582276
rect 151044 582256 151046 582276
rect 151174 582256 151230 582312
rect 156602 582256 156658 582312
rect 155866 581984 155922 582040
rect 156326 581984 156382 582040
rect 157154 581984 157210 582040
rect 147862 581576 147918 581632
rect 153934 581576 153990 581632
rect 156602 581576 156658 581632
rect 157062 581440 157118 581496
rect 162490 582276 162546 582312
rect 162490 582256 162492 582276
rect 162492 582256 162544 582276
rect 162544 582256 162546 582276
rect 166814 582256 166870 582312
rect 157522 581440 157578 581496
rect 166998 582256 167054 582312
rect 167090 581984 167146 582040
rect 182178 584704 182234 584760
rect 182270 584432 182326 584488
rect 175094 584296 175150 584352
rect 171598 582256 171654 582312
rect 171782 582256 171838 582312
rect 166998 581576 167054 581632
rect 108946 581304 109002 581360
rect 109130 581304 109186 581360
rect 115202 581304 115258 581360
rect 115846 581304 115902 581360
rect 118698 581304 118754 581360
rect 146942 581304 146998 581360
rect 147862 581304 147918 581360
rect 157246 581304 157302 581360
rect 166906 581304 166962 581360
rect 179878 583888 179934 583944
rect 176566 581984 176622 582040
rect 181442 582256 181498 582312
rect 171782 581440 171838 581496
rect 171966 581440 172022 581496
rect 186870 583888 186926 583944
rect 186318 581984 186374 582040
rect 191746 584860 191802 584896
rect 191746 584840 191748 584860
rect 191748 584840 191800 584860
rect 191800 584840 191802 584860
rect 205638 584976 205694 585032
rect 225142 584976 225198 585032
rect 205546 584840 205602 584896
rect 218150 584840 218206 584896
rect 201222 584024 201278 584080
rect 196438 582392 196494 582448
rect 190826 582256 190882 582312
rect 191654 582120 191710 582176
rect 192022 582120 192078 582176
rect 181442 581440 181498 581496
rect 190826 581440 190882 581496
rect 195886 581984 195942 582040
rect 200762 582256 200818 582312
rect 200670 582120 200726 582176
rect 198002 581612 198004 581632
rect 198004 581612 198056 581632
rect 198056 581612 198058 581632
rect 198002 581576 198058 581612
rect 200854 582120 200910 582176
rect 206006 582528 206062 582584
rect 203338 581984 203394 582040
rect 210330 581984 210386 582040
rect 208306 581848 208362 581904
rect 200762 581440 200818 581496
rect 210422 581848 210478 581904
rect 213182 582800 213238 582856
rect 211158 582256 211214 582312
rect 210422 581440 210478 581496
rect 218058 584704 218114 584760
rect 222750 584024 222806 584080
rect 220082 581848 220138 581904
rect 220910 581984 220966 582040
rect 220726 581848 220782 581904
rect 220082 581440 220138 581496
rect 227718 584840 227774 584896
rect 234526 584704 234582 584760
rect 233238 584432 233294 584488
rect 234526 583752 234582 583808
rect 229374 582120 229430 582176
rect 229466 581984 229522 582040
rect 230110 581848 230166 581904
rect 236458 581984 236514 582040
rect 229466 581440 229522 581496
rect 238758 584724 238814 584760
rect 238758 584704 238760 584724
rect 238760 584704 238812 584724
rect 238812 584704 238814 584724
rect 241702 584160 241758 584216
rect 238758 581984 238814 582040
rect 236458 581440 236514 581496
rect 239034 581848 239090 581904
rect 249246 581848 249302 581904
rect 258446 584160 258502 584216
rect 258354 582120 258410 582176
rect 258170 581984 258226 582040
rect 256238 581848 256294 581904
rect 256330 581576 256386 581632
rect 253386 581440 253442 581496
rect 256238 581440 256294 581496
rect 291750 584568 291806 584624
rect 275006 584432 275062 584488
rect 273166 582120 273222 582176
rect 277398 584296 277454 584352
rect 282918 582256 282974 582312
rect 282550 581848 282606 581904
rect 292486 582256 292542 582312
rect 315670 584568 315726 584624
rect 298926 583752 298982 583808
rect 303710 582936 303766 582992
rect 301318 582664 301374 582720
rect 302238 582256 302294 582312
rect 306286 581984 306342 582040
rect 314658 582936 314714 582992
rect 311806 582256 311862 582312
rect 318062 582800 318118 582856
rect 326434 582120 326490 582176
rect 329838 582120 329894 582176
rect 331954 581712 332010 581768
rect 348790 700304 348846 700360
rect 372618 584704 372674 584760
rect 412914 585656 412970 585712
rect 427542 584840 427598 584896
rect 424966 582120 425022 582176
rect 465630 584704 465686 584760
rect 451462 583752 451518 583808
rect 472806 584704 472862 584760
rect 490194 582256 490250 582312
rect 490378 582256 490434 582312
rect 491850 582120 491906 582176
rect 418158 581712 418214 581768
rect 273166 581576 273222 581632
rect 282918 581576 282974 581632
rect 292486 581576 292542 581632
rect 302238 581576 302294 581632
rect 311806 581576 311862 581632
rect 321558 581576 321614 581632
rect 324778 581576 324834 581632
rect 346858 581576 346914 581632
rect 351642 581576 351698 581632
rect 365258 581576 365314 581632
rect 384854 581576 384910 581632
rect 389730 581576 389786 581632
rect 391754 581576 391810 581632
rect 396998 581576 397054 581632
rect 263506 581440 263562 581496
rect 263690 581440 263746 581496
rect 494610 583888 494666 583944
rect 496726 583888 496782 583944
rect 497554 581984 497610 582040
rect 176566 581304 176622 581360
rect 176750 581304 176806 581360
rect 192022 581304 192078 581360
rect 192206 581304 192262 581360
rect 195886 581304 195942 581360
rect 200670 581304 200726 581360
rect 210330 581304 210386 581360
rect 211158 581304 211214 581360
rect 220726 581304 220782 581360
rect 220910 581304 220966 581360
rect 229374 581304 229430 581360
rect 230110 581304 230166 581360
rect 231950 581304 232006 581360
rect 238758 581304 238814 581360
rect 239034 581304 239090 581360
rect 239678 581304 239734 581360
rect 249246 581304 249302 581360
rect 256330 581304 256386 581360
rect 258170 581304 258226 581360
rect 258354 581304 258410 581360
rect 263506 581304 263562 581360
rect 263690 581304 263746 581360
rect 358726 581304 358782 581360
rect 82634 541456 82690 541512
rect 82358 518744 82414 518800
rect 82358 509496 82414 509552
rect 82542 505688 82598 505744
rect 82358 500792 82414 500848
rect 82542 498072 82598 498128
rect 82358 497120 82414 497176
rect 82542 486104 82598 486160
rect 82358 481208 82414 481264
rect 82542 481072 82598 481128
rect 82542 475768 82598 475824
rect 82450 474136 82506 474192
rect 82358 473592 82414 473648
rect 82634 474272 82690 474328
rect 82542 473456 82598 473512
rect 82542 471008 82598 471064
rect 82450 466112 82506 466168
rect 82542 457952 82598 458008
rect 82634 453328 82690 453384
rect 101586 456456 101642 456512
rect 101494 451832 101550 451888
rect 82542 438912 82598 438968
rect 82542 435376 82598 435432
rect 82542 431160 82598 431216
rect 82542 406408 82598 406464
rect 82542 401512 82598 401568
rect 82358 400152 82414 400208
rect 82266 391176 82322 391232
rect 82082 391040 82138 391096
rect 82450 396752 82506 396808
rect 82450 396072 82506 396128
rect 82634 393080 82690 393136
rect 82542 385736 82598 385792
rect 82082 385600 82138 385656
rect 82358 385600 82414 385656
rect 82450 371864 82506 371920
rect 82358 369008 82414 369064
rect 82542 369008 82598 369064
rect 82450 368056 82506 368112
rect 82634 368872 82690 368928
rect 82634 368736 82690 368792
rect 82450 364792 82506 364848
rect 82358 364656 82414 364712
rect 82358 362888 82414 362944
rect 82358 360168 82414 360224
rect 82634 362752 82690 362808
rect 82634 360032 82690 360088
rect 82450 359352 82506 359408
rect 82634 357992 82690 358048
rect 82082 354592 82138 354648
rect 82542 346976 82598 347032
rect 82174 339632 82230 339688
rect 82358 338952 82414 339008
rect 82174 338000 82230 338056
rect 82174 332152 82230 332208
rect 82634 341672 82690 341728
rect 82542 336912 82598 336968
rect 82542 335008 82598 335064
rect 82358 331200 82414 331256
rect 82634 331200 82690 331256
rect 82542 331064 82598 331120
rect 82174 328072 82230 328128
rect 82634 319504 82690 319560
rect 82450 317328 82506 317384
rect 82450 316240 82506 316296
rect 82634 312432 82690 312488
rect 82450 312296 82506 312352
rect 82450 307400 82506 307456
rect 82634 305360 82690 305416
rect 82174 301824 82230 301880
rect 82082 123528 82138 123584
rect 82542 297744 82598 297800
rect 82358 296792 82414 296848
rect 82266 294752 82322 294808
rect 82358 291216 82414 291272
rect 82634 297472 82690 297528
rect 82634 292032 82690 292088
rect 82542 289040 82598 289096
rect 82634 269592 82690 269648
rect 82450 266192 82506 266248
rect 82634 264016 82690 264072
rect 82450 260208 82506 260264
rect 82542 254768 82598 254824
rect 82542 252728 82598 252784
rect 82358 245520 82414 245576
rect 88706 247968 88762 248024
rect 88430 247696 88486 247752
rect 82542 239400 82598 239456
rect 82450 238312 82506 238368
rect 82450 235068 82506 235104
rect 82450 235048 82452 235068
rect 82452 235048 82504 235068
rect 82504 235048 82506 235068
rect 82450 234912 82506 234968
rect 82634 236952 82690 237008
rect 82634 234776 82690 234832
rect 82634 233416 82690 233472
rect 82634 232620 82690 232656
rect 82634 232600 82636 232620
rect 82636 232600 82688 232620
rect 82688 232600 82690 232620
rect 82542 232328 82598 232384
rect 82634 225664 82690 225720
rect 82634 224304 82690 224360
rect 82634 209344 82690 209400
rect 82634 195200 82690 195256
rect 82634 195084 82690 195120
rect 82634 195064 82636 195084
rect 82636 195064 82688 195084
rect 82688 195064 82690 195084
rect 82634 194948 82690 194984
rect 82634 194928 82636 194948
rect 82636 194928 82688 194948
rect 82688 194928 82690 194948
rect 82634 194812 82690 194848
rect 82634 194792 82636 194812
rect 82636 194792 82688 194812
rect 82688 194792 82690 194812
rect 82634 194656 82690 194712
rect 82634 191140 82690 191176
rect 82634 191120 82636 191140
rect 82636 191120 82688 191140
rect 82688 191120 82690 191140
rect 82634 190848 82690 190904
rect 82542 190732 82598 190768
rect 82542 190712 82544 190732
rect 82544 190712 82596 190732
rect 82596 190712 82598 190732
rect 82542 190476 82544 190496
rect 82544 190476 82596 190496
rect 82596 190476 82598 190496
rect 82542 190440 82598 190476
rect 82542 189216 82598 189272
rect 82634 188672 82690 188728
rect 82634 187312 82690 187368
rect 82634 187040 82690 187096
rect 82634 186940 82636 186960
rect 82636 186940 82688 186960
rect 82688 186940 82690 186960
rect 82634 186904 82690 186940
rect 82634 170212 82636 170232
rect 82636 170212 82688 170232
rect 82688 170212 82690 170232
rect 82634 170176 82690 170212
rect 82634 170076 82636 170096
rect 82636 170076 82688 170096
rect 82688 170076 82690 170096
rect 82634 170040 82690 170076
rect 82634 157392 82690 157448
rect 82634 128968 82690 129024
rect 82634 122848 82690 122904
rect 83002 123800 83058 123856
rect 83094 123664 83150 123720
rect 83370 123800 83426 123856
rect 83186 117952 83242 118008
rect 83554 123800 83610 123856
rect 83646 123256 83702 123312
rect 88706 233008 88762 233064
rect 87878 232736 87934 232792
rect 84566 226752 84622 226808
rect 86130 226752 86186 226808
rect 87326 179832 87382 179888
rect 88706 179832 88762 179888
rect 87326 171536 87382 171592
rect 87602 171536 87658 171592
rect 501786 518064 501842 518120
rect 501786 517248 501842 517304
rect 501786 506912 501842 506968
rect 501786 474816 501842 474872
rect 501786 464208 501842 464264
rect 501786 457136 501842 457192
rect 501694 158888 501750 158944
rect 501602 157428 501604 157448
rect 501604 157428 501656 157448
rect 501656 157428 501658 157448
rect 501602 157392 501658 157428
rect 501694 156576 501750 156632
rect 501510 151836 501566 151872
rect 501510 151816 501512 151836
rect 501512 151816 501564 151836
rect 501564 151816 501566 151836
rect 501694 154708 501696 154728
rect 501696 154708 501748 154728
rect 501748 154708 501750 154728
rect 501694 154672 501750 154708
rect 501694 136312 501750 136368
rect 501602 126112 501658 126168
rect 87510 122576 87566 122632
rect 88982 122576 89038 122632
rect 89258 122576 89314 122632
rect 90638 122576 90694 122632
rect 92294 122576 92350 122632
rect 101034 122576 101090 122632
rect 86866 122304 86922 122360
rect 83830 122168 83886 122224
rect 84106 120672 84162 120728
rect 83186 106256 83242 106312
rect 83278 104760 83334 104816
rect 83278 95240 83334 95296
rect 83278 86808 83334 86864
rect 83278 77288 83334 77344
rect 83278 77016 83334 77072
rect 83278 67632 83334 67688
rect 83278 57840 83334 57896
rect 83278 48320 83334 48376
rect 83278 38528 83334 38584
rect 83278 29144 83334 29200
rect 83278 19080 83334 19136
rect 83278 15816 83334 15872
rect 82726 13912 82782 13968
rect 82634 13776 82690 13832
rect 83922 15952 83978 16008
rect 84290 106936 84346 106992
rect 84290 98640 84346 98696
rect 84382 86264 84438 86320
rect 84382 77968 84438 78024
rect 84382 23296 84438 23352
rect 84382 13776 84438 13832
rect 84382 13640 84438 13696
rect 81438 3848 81494 3904
rect 82634 5344 82690 5400
rect 82542 3440 82598 3496
rect 88982 121760 89038 121816
rect 88430 120672 88486 120728
rect 86038 116864 86094 116920
rect 84382 4120 84438 4176
rect 87142 116728 87198 116784
rect 87326 116728 87382 116784
rect 86590 111152 86646 111208
rect 86590 106936 86646 106992
rect 86038 106392 86094 106448
rect 89258 119992 89314 120048
rect 95330 122168 95386 122224
rect 96710 119312 96766 119368
rect 88246 106256 88302 106312
rect 88430 106256 88486 106312
rect 87142 105848 87198 105904
rect 88246 101496 88302 101552
rect 88154 96464 88210 96520
rect 87970 96328 88026 96384
rect 88154 94560 88210 94616
rect 87970 92656 88026 92712
rect 87142 86264 87198 86320
rect 87142 77968 87198 78024
rect 87602 77968 87658 78024
rect 88246 77968 88302 78024
rect 88246 69128 88302 69184
rect 87602 67632 87658 67688
rect 85762 62736 85818 62792
rect 87510 57840 87566 57896
rect 85762 48456 85818 48512
rect 87510 48320 87566 48376
rect 85854 43424 85910 43480
rect 85854 37440 85910 37496
rect 87510 35264 87566 35320
rect 85854 27512 85910 27568
rect 87510 23432 87566 23488
rect 86406 22752 86462 22808
rect 85946 19216 86002 19272
rect 85854 18128 85910 18184
rect 85946 9832 86002 9888
rect 86222 9424 86278 9480
rect 86130 4664 86186 4720
rect 85578 3440 85634 3496
rect 87786 8064 87842 8120
rect 87786 5752 87842 5808
rect 86406 4120 86462 4176
rect 86222 3168 86278 3224
rect 88522 3848 88578 3904
rect 90730 3848 90786 3904
rect 90914 3848 90970 3904
rect 90730 3440 90786 3496
rect 99102 16088 99158 16144
rect 95146 3576 95202 3632
rect 94502 2896 94558 2952
rect 99378 2760 99434 2816
rect 105358 121080 105414 121136
rect 107566 3032 107622 3088
rect 108762 3032 108818 3088
rect 108946 3032 109002 3088
rect 108946 2760 109002 2816
rect 117778 121488 117834 121544
rect 118422 115912 118478 115968
rect 117318 71712 117374 71768
rect 117502 71712 117558 71768
rect 117502 52400 117558 52456
rect 117686 52400 117742 52456
rect 115754 3732 115810 3768
rect 115754 3712 115756 3732
rect 115756 3712 115808 3732
rect 115808 3712 115810 3732
rect 115938 3712 115994 3768
rect 116858 3732 116914 3768
rect 116858 3712 116860 3732
rect 116860 3712 116912 3732
rect 116912 3712 116914 3732
rect 114742 2896 114798 2952
rect 124218 122576 124274 122632
rect 124218 122168 124274 122224
rect 121366 115776 121422 115832
rect 120078 71712 120134 71768
rect 120262 71712 120318 71768
rect 120262 52400 120318 52456
rect 120446 52400 120502 52456
rect 120078 24792 120134 24848
rect 120354 24792 120410 24848
rect 118698 2760 118754 2816
rect 133786 122576 133842 122632
rect 143538 122576 143594 122632
rect 149058 122576 149114 122632
rect 153106 122612 153108 122632
rect 153108 122612 153160 122632
rect 153160 122612 153162 122632
rect 153106 122576 153162 122612
rect 201314 122576 201370 122632
rect 216586 122576 216642 122632
rect 133786 122168 133842 122224
rect 143538 122168 143594 122224
rect 122010 3440 122066 3496
rect 123022 3440 123078 3496
rect 122010 2896 122066 2952
rect 122930 2760 122986 2816
rect 125414 2896 125470 2952
rect 131210 122032 131266 122088
rect 130014 119584 130070 119640
rect 140686 122032 140742 122088
rect 139582 119720 139638 119776
rect 142158 121624 142214 121680
rect 141974 119448 142030 119504
rect 146390 121760 146446 121816
rect 146206 119584 146262 119640
rect 143446 3576 143502 3632
rect 143446 2896 143502 2952
rect 179418 122440 179474 122496
rect 153106 122168 153162 122224
rect 162858 122168 162914 122224
rect 149058 121896 149114 121952
rect 149058 121760 149114 121816
rect 148046 3440 148102 3496
rect 153198 121896 153254 121952
rect 153106 119720 153162 119776
rect 152922 70352 152978 70408
rect 152830 67632 152886 67688
rect 152922 61376 152978 61432
rect 153014 50904 153070 50960
rect 151726 10240 151782 10296
rect 153106 3576 153162 3632
rect 158718 121352 158774 121408
rect 153106 2896 153162 2952
rect 165526 17312 165582 17368
rect 162122 3712 162178 3768
rect 162766 3576 162822 3632
rect 163502 3712 163558 3768
rect 164698 3712 164754 3768
rect 162122 3440 162178 3496
rect 162858 3440 162914 3496
rect 162858 3304 162914 3360
rect 163318 3304 163374 3360
rect 162766 2896 162822 2952
rect 167090 122304 167146 122360
rect 169666 122304 169722 122360
rect 168286 121488 168342 121544
rect 172426 122168 172482 122224
rect 172610 122168 172666 122224
rect 172518 122052 172574 122088
rect 172518 122032 172520 122052
rect 172520 122032 172572 122052
rect 172572 122032 172574 122052
rect 172794 122052 172850 122088
rect 172794 122032 172796 122052
rect 172796 122032 172848 122052
rect 172848 122032 172850 122052
rect 173898 121760 173954 121816
rect 176658 118768 176714 118824
rect 175370 3440 175426 3496
rect 179326 67768 179382 67824
rect 179326 67632 179382 67688
rect 209686 122440 209742 122496
rect 201406 122304 201462 122360
rect 182086 122168 182142 122224
rect 182362 122168 182418 122224
rect 191746 122168 191802 122224
rect 182454 121216 182510 121272
rect 182086 3576 182142 3632
rect 187238 121216 187294 121272
rect 190458 119176 190514 119232
rect 187698 118904 187754 118960
rect 182086 2896 182142 2952
rect 190366 17448 190422 17504
rect 193218 119040 193274 119096
rect 195426 14592 195482 14648
rect 196622 122032 196678 122088
rect 196622 121760 196678 121816
rect 195426 9696 195482 9752
rect 195610 9696 195666 9752
rect 199934 16224 199990 16280
rect 201498 119856 201554 119912
rect 204166 16360 204222 16416
rect 212262 122304 212318 122360
rect 212446 122304 212502 122360
rect 206926 3712 206982 3768
rect 207478 3712 207534 3768
rect 206926 3440 206982 3496
rect 217966 115232 218022 115288
rect 220266 37304 220322 37360
rect 220450 37304 220506 37360
rect 223578 9832 223634 9888
rect 223578 9662 223634 9718
rect 219346 3712 219402 3768
rect 220082 3712 220138 3768
rect 218150 2896 218206 2952
rect 220082 3440 220138 3496
rect 220266 3440 220322 3496
rect 220266 2896 220322 2952
rect 223578 8200 223634 8256
rect 224222 8064 224278 8120
rect 237102 121896 237158 121952
rect 230110 5752 230166 5808
rect 240046 122168 240102 122224
rect 240322 122168 240378 122224
rect 239862 121624 239918 121680
rect 241518 122168 241574 122224
rect 249798 122168 249854 122224
rect 242806 120672 242862 120728
rect 241518 3576 241574 3632
rect 238390 3032 238446 3088
rect 241518 2760 241574 2816
rect 248326 121896 248382 121952
rect 259366 122168 259422 122224
rect 278686 122168 278742 122224
rect 258078 9696 258134 9752
rect 258262 9696 258318 9752
rect 273166 120808 273222 120864
rect 266082 111152 266138 111208
rect 253846 3032 253902 3088
rect 257434 3712 257490 3768
rect 259826 3712 259882 3768
rect 259366 3576 259422 3632
rect 259366 2760 259422 2816
rect 263414 3848 263470 3904
rect 267002 5208 267058 5264
rect 272614 106120 272670 106176
rect 272890 106120 272946 106176
rect 271510 3984 271566 4040
rect 271694 3984 271750 4040
rect 270498 3712 270554 3768
rect 271510 3032 271566 3088
rect 278686 121760 278742 121816
rect 276018 111172 276074 111208
rect 276018 111152 276020 111172
rect 276020 111152 276072 111172
rect 276072 111152 276074 111172
rect 275282 3984 275338 4040
rect 278870 3984 278926 4040
rect 280066 3032 280122 3088
rect 282458 5072 282514 5128
rect 285494 111172 285550 111208
rect 285494 111152 285496 111172
rect 285496 111152 285548 111172
rect 285548 111152 285550 111172
rect 500130 122576 500186 122632
rect 500314 122576 500370 122632
rect 500498 122576 500554 122632
rect 298006 122168 298062 122224
rect 318614 122168 318670 122224
rect 318798 122168 318854 122224
rect 336646 122168 336702 122224
rect 289542 86944 289598 87000
rect 289726 119856 289782 119912
rect 289726 97008 289782 97064
rect 289726 96620 289782 96656
rect 289726 96600 289728 96620
rect 289728 96600 289780 96620
rect 289780 96600 289782 96620
rect 289726 86944 289782 87000
rect 290738 8880 290794 8936
rect 289726 8200 289782 8256
rect 289910 8200 289966 8256
rect 296626 119176 296682 119232
rect 295338 111188 295340 111208
rect 295340 111188 295392 111208
rect 295392 111188 295394 111208
rect 295338 111152 295394 111188
rect 298006 121624 298062 121680
rect 304906 111152 304962 111208
rect 297914 19080 297970 19136
rect 298006 3576 298062 3632
rect 299110 3168 299166 3224
rect 298006 3032 298062 3088
rect 301410 3168 301466 3224
rect 322846 121760 322902 121816
rect 320638 119992 320694 120048
rect 317326 119040 317382 119096
rect 314658 111172 314714 111208
rect 314658 111152 314660 111172
rect 314660 111152 314712 111172
rect 314712 111152 314714 111172
rect 315946 19080 316002 19136
rect 314566 18944 314622 19000
rect 315946 18808 316002 18864
rect 318062 5888 318118 5944
rect 318890 4120 318946 4176
rect 318798 3984 318854 4040
rect 319258 3712 319314 3768
rect 323582 111172 323638 111208
rect 323582 111152 323584 111172
rect 323584 111152 323636 111172
rect 323636 111152 323638 111172
rect 325698 19080 325754 19136
rect 325698 18808 325754 18864
rect 325238 6024 325294 6080
rect 328366 120944 328422 121000
rect 328458 111424 328514 111480
rect 328458 111152 328514 111208
rect 330942 121624 330998 121680
rect 331126 84768 331182 84824
rect 332598 3576 332654 3632
rect 332598 3032 332654 3088
rect 332414 2896 332470 2952
rect 338118 121796 338120 121816
rect 338120 121796 338172 121816
rect 338172 121796 338174 121816
rect 338118 121760 338174 121796
rect 335910 19080 335966 19136
rect 335910 18808 335966 18864
rect 335358 3576 335414 3632
rect 335358 3032 335414 3088
rect 342994 121796 342996 121816
rect 342996 121796 343048 121816
rect 343048 121796 343050 121816
rect 342994 121760 343050 121796
rect 343546 111152 343602 111208
rect 343730 111152 343786 111208
rect 345018 19080 345074 19136
rect 345018 18808 345074 18864
rect 343086 3712 343142 3768
rect 355966 122168 356022 122224
rect 353298 111172 353354 111208
rect 353298 111152 353300 111172
rect 353300 111152 353352 111172
rect 353352 111152 353354 111172
rect 355966 121624 356022 121680
rect 355322 19080 355378 19136
rect 355322 18808 355378 18864
rect 353758 8880 353814 8936
rect 351826 3712 351882 3768
rect 351826 3032 351882 3088
rect 356794 3984 356850 4040
rect 357254 3984 357310 4040
rect 356978 3848 357034 3904
rect 357254 3848 357310 3904
rect 362774 111172 362830 111208
rect 362774 111152 362776 111172
rect 362776 111152 362828 111172
rect 362828 111152 362830 111172
rect 364338 19080 364394 19136
rect 364338 18808 364394 18864
rect 375286 122168 375342 122224
rect 376758 122168 376814 122224
rect 375286 121624 375342 121680
rect 371330 116728 371386 116784
rect 372710 111188 372712 111208
rect 372712 111188 372764 111208
rect 372764 111188 372766 111208
rect 372710 111152 372766 111188
rect 369214 10512 369270 10568
rect 386142 122168 386198 122224
rect 404358 122168 404414 122224
rect 375286 115368 375342 115424
rect 382094 111188 382096 111208
rect 382096 111188 382148 111208
rect 382148 111188 382150 111208
rect 382094 111152 382150 111188
rect 378138 111036 378194 111072
rect 378138 111016 378140 111036
rect 378140 111016 378192 111036
rect 378192 111016 378194 111036
rect 378782 19080 378838 19136
rect 383658 19080 383714 19136
rect 378782 18808 378838 18864
rect 383658 18808 383714 18864
rect 389638 119992 389694 120048
rect 389822 119992 389878 120048
rect 389638 118632 389694 118688
rect 386510 111152 386566 111208
rect 386510 110880 386566 110936
rect 387062 6840 387118 6896
rect 390650 6704 390706 6760
rect 389454 6568 389510 6624
rect 394606 4120 394662 4176
rect 394606 3712 394662 3768
rect 400862 3712 400918 3768
rect 400862 3032 400918 3088
rect 401690 111152 401746 111208
rect 401690 110608 401746 110664
rect 413926 122168 413982 122224
rect 415490 122168 415546 122224
rect 403714 6568 403770 6624
rect 405646 3712 405702 3768
rect 407302 6704 407358 6760
rect 424966 122168 425022 122224
rect 426438 122168 426494 122224
rect 411258 111188 411260 111208
rect 411260 111188 411312 111208
rect 411312 111188 411314 111208
rect 411258 111152 411314 111188
rect 412546 19080 412602 19136
rect 412546 18808 412602 18864
rect 414478 6432 414534 6488
rect 419446 121624 419502 121680
rect 420734 111188 420736 111208
rect 420736 111188 420788 111208
rect 420788 111188 420790 111208
rect 420734 111152 420790 111188
rect 425610 35128 425666 35184
rect 422298 19080 422354 19136
rect 422298 18808 422354 18864
rect 430578 111172 430634 111208
rect 430578 111152 430580 111172
rect 430580 111152 430632 111172
rect 430632 111152 430634 111172
rect 422758 6432 422814 6488
rect 425150 3576 425206 3632
rect 425058 2896 425114 2952
rect 427634 9696 427690 9752
rect 427818 9696 427874 9752
rect 432050 19080 432106 19136
rect 432050 18808 432106 18864
rect 435822 77152 435878 77208
rect 435822 67632 435878 67688
rect 433522 10376 433578 10432
rect 436098 86964 436154 87000
rect 436098 86944 436100 86964
rect 436100 86944 436152 86964
rect 436152 86944 436154 86964
rect 436282 86944 436338 87000
rect 436098 77152 436154 77208
rect 436098 67632 436154 67688
rect 437478 11736 437534 11792
rect 435822 3576 435878 3632
rect 440146 111152 440202 111208
rect 441618 19080 441674 19136
rect 441618 18808 441674 18864
rect 444470 111152 444526 111208
rect 444470 110880 444526 110936
rect 442262 3712 442318 3768
rect 442998 3032 443054 3088
rect 442262 2896 442318 2952
rect 447138 19080 447194 19136
rect 447138 18808 447194 18864
rect 448518 18672 448574 18728
rect 453946 39208 454002 39264
rect 451462 3712 451518 3768
rect 451462 2760 451518 2816
rect 458178 115096 458234 115152
rect 459650 111152 459706 111208
rect 459650 110608 459706 110664
rect 462594 18808 462650 18864
rect 462594 18400 462650 18456
rect 460846 3304 460902 3360
rect 459650 2896 459706 2952
rect 465630 6840 465686 6896
rect 463238 3712 463294 3768
rect 463698 3712 463754 3768
rect 464434 3304 464490 3360
rect 463698 2760 463754 2816
rect 469218 111424 469274 111480
rect 469218 111152 469274 111208
rect 470322 6024 470378 6080
rect 470598 3712 470654 3768
rect 470598 2760 470654 2816
rect 478786 111152 478842 111208
rect 478970 111152 479026 111208
rect 478142 19080 478198 19136
rect 478142 18400 478198 18456
rect 478694 3712 478750 3768
rect 481730 17176 481786 17232
rect 482374 3712 482430 3768
rect 485686 19080 485742 19136
rect 485686 18672 485742 18728
rect 482374 2760 482430 2816
rect 486974 2760 487030 2816
rect 488538 111288 488594 111344
rect 488538 111152 488594 111208
rect 490562 2760 490618 2816
rect 496082 121080 496138 121136
rect 493506 117156 493562 117192
rect 493506 117136 493508 117156
rect 493508 117136 493560 117156
rect 493560 117136 493562 117156
rect 494702 3984 494758 4040
rect 495070 3712 495126 3768
rect 496726 118904 496782 118960
rect 499210 121352 499266 121408
rect 499394 121388 499396 121408
rect 499396 121388 499448 121408
rect 499448 121388 499450 121408
rect 499394 121352 499450 121388
rect 499854 121352 499910 121408
rect 499118 121216 499174 121272
rect 499302 121216 499358 121272
rect 498382 120944 498438 121000
rect 498566 120944 498622 121000
rect 498382 120536 498438 120592
rect 498934 120536 498990 120592
rect 499946 120672 500002 120728
rect 499118 120400 499174 120456
rect 500038 120264 500094 120320
rect 498566 116728 498622 116784
rect 500130 113328 500186 113384
rect 500130 109656 500186 109712
rect 500130 96736 500186 96792
rect 499946 95104 500002 95160
rect 500406 120944 500462 121000
rect 500314 117952 500370 118008
rect 501602 123528 501658 123584
rect 501602 123428 501604 123448
rect 501604 123428 501656 123448
rect 501656 123428 501658 123448
rect 501602 123392 501658 123428
rect 500406 114552 500462 114608
rect 500774 104624 500830 104680
rect 500590 92792 500646 92848
rect 500682 92656 500738 92712
rect 500590 91704 500646 91760
rect 499394 72936 499450 72992
rect 498382 67496 498438 67552
rect 498382 62736 498438 62792
rect 498382 57704 498438 57760
rect 500038 56752 500094 56808
rect 499394 55392 499450 55448
rect 500406 77152 500462 77208
rect 500774 86944 500830 87000
rect 500406 68312 500462 68368
rect 500498 56480 500554 56536
rect 499946 49000 500002 49056
rect 498382 48320 498438 48376
rect 500406 49000 500462 49056
rect 500498 48864 500554 48920
rect 500406 39208 500462 39264
rect 499946 38800 500002 38856
rect 498290 34312 498346 34368
rect 498290 25064 498346 25120
rect 498474 15272 498530 15328
rect 500590 37168 500646 37224
rect 500590 29688 500646 29744
rect 499946 15136 500002 15192
rect 500222 15136 500278 15192
rect 498474 9696 498530 9752
rect 495622 3984 495678 4040
rect 495530 3848 495586 3904
rect 500038 3576 500094 3632
rect 502062 573688 502118 573744
rect 502062 572192 502118 572248
rect 502062 557096 502118 557152
rect 502062 547848 502118 547904
rect 502062 500520 502118 500576
rect 502062 493312 502118 493368
rect 502154 464344 502210 464400
rect 502154 454824 502210 454880
rect 502062 454688 502118 454744
rect 502062 448976 502118 449032
rect 501970 442448 502026 442504
rect 501970 439728 502026 439784
rect 502154 427760 502210 427816
rect 502062 423408 502118 423464
rect 502154 418240 502210 418296
rect 502062 414024 502118 414080
rect 502062 413752 502118 413808
rect 501970 411440 502026 411496
rect 501970 410080 502026 410136
rect 501970 405728 502026 405784
rect 502062 405592 502118 405648
rect 502062 403688 502118 403744
rect 501970 400696 502026 400752
rect 502062 398656 502118 398712
rect 502246 394576 502302 394632
rect 502246 387096 502302 387152
rect 501970 351600 502026 351656
rect 502062 350512 502118 350568
rect 502062 346432 502118 346488
rect 501970 346296 502026 346352
rect 502154 344936 502210 344992
rect 502154 338816 502210 338872
rect 502062 337456 502118 337512
rect 501970 325624 502026 325680
rect 501970 315832 502026 315888
rect 501970 308488 502026 308544
rect 501970 290400 502026 290456
rect 501970 290284 502026 290320
rect 501970 290264 501972 290284
rect 501972 290264 502024 290284
rect 502024 290264 502026 290284
rect 501970 290128 502026 290184
rect 501970 282376 502026 282432
rect 501970 282260 502026 282296
rect 501970 282240 501972 282260
rect 501972 282240 502024 282260
rect 502024 282240 502026 282260
rect 501970 281424 502026 281480
rect 501970 275032 502026 275088
rect 501970 273128 502026 273184
rect 501970 272620 501972 272640
rect 501972 272620 502024 272640
rect 502024 272620 502026 272640
rect 501970 272584 502026 272620
rect 501970 272484 501972 272504
rect 501972 272484 502024 272504
rect 502024 272484 502026 272504
rect 501970 272448 502026 272484
rect 501970 272348 501972 272368
rect 501972 272348 502024 272368
rect 502024 272348 502026 272368
rect 501970 272312 502026 272348
rect 501970 270852 501972 270872
rect 501972 270852 502024 270872
rect 502024 270852 502026 270872
rect 501970 270816 502026 270852
rect 501970 270428 502026 270464
rect 501970 270408 501972 270428
rect 501972 270408 502024 270428
rect 502024 270408 502026 270428
rect 501970 268232 502026 268288
rect 501970 267028 502026 267064
rect 501970 267008 501972 267028
rect 501972 267008 502024 267028
rect 502024 267008 502026 267028
rect 501970 263472 502026 263528
rect 501878 155216 501934 155272
rect 501878 140548 501934 140584
rect 501878 140528 501880 140548
rect 501880 140528 501932 140548
rect 501932 140528 501934 140548
rect 501878 140412 501934 140448
rect 501878 140392 501880 140412
rect 501880 140392 501932 140412
rect 501932 140392 501934 140412
rect 501878 140276 501934 140312
rect 501878 140256 501880 140276
rect 501880 140256 501932 140276
rect 501932 140256 501934 140276
rect 501878 140140 501934 140176
rect 501878 140120 501880 140140
rect 501880 140120 501932 140140
rect 501932 140120 501934 140140
rect 501878 140004 501934 140040
rect 501878 139984 501880 140004
rect 501880 139984 501932 140004
rect 501932 139984 501934 140004
rect 501878 138760 501934 138816
rect 501878 137828 501934 137864
rect 501878 137808 501880 137828
rect 501880 137808 501932 137828
rect 501932 137808 501934 137828
rect 501878 137028 501880 137048
rect 501880 137028 501932 137048
rect 501932 137028 501934 137048
rect 501878 136992 501934 137028
rect 501878 136720 501934 136776
rect 501878 120672 501934 120728
rect 502154 320320 502210 320376
rect 502246 289992 502302 290048
rect 502246 278160 502302 278216
rect 502154 209208 502210 209264
rect 502154 198056 502210 198112
rect 502062 124888 502118 124944
rect 502154 123800 502210 123856
rect 502154 123700 502156 123720
rect 502156 123700 502208 123720
rect 502208 123700 502210 123720
rect 502154 123664 502210 123700
rect 502062 122712 502118 122768
rect 502062 120944 502118 121000
rect 502062 118224 502118 118280
rect 502430 415520 502486 415576
rect 502338 148844 502394 148880
rect 502338 148824 502340 148844
rect 502340 148824 502392 148844
rect 502392 148824 502394 148844
rect 502338 147484 502394 147520
rect 502338 147464 502340 147484
rect 502340 147464 502392 147484
rect 502392 147464 502394 147484
rect 502338 147228 502340 147248
rect 502340 147228 502392 147248
rect 502392 147228 502394 147248
rect 502338 147192 502394 147228
rect 502338 146920 502394 146976
rect 502338 138352 502394 138408
rect 502338 138252 502340 138272
rect 502340 138252 502392 138272
rect 502392 138252 502394 138272
rect 502338 138216 502394 138252
rect 502338 137436 502340 137456
rect 502340 137436 502392 137456
rect 502392 137436 502394 137456
rect 502338 137400 502394 137436
rect 502338 137264 502394 137320
rect 502706 582800 502762 582856
rect 502706 575456 502762 575512
rect 502890 433200 502946 433256
rect 502890 425040 502946 425096
rect 502614 401376 502670 401432
rect 502614 397840 502670 397896
rect 502522 316784 502578 316840
rect 502522 302912 502578 302968
rect 502706 383696 502762 383752
rect 502614 124616 502670 124672
rect 502614 122168 502670 122224
rect 502798 359216 502854 359272
rect 502890 327392 502946 327448
rect 503902 580352 503958 580408
rect 503718 579672 503774 579728
rect 503718 574096 503774 574152
rect 503810 567024 503866 567080
rect 503810 563488 503866 563544
rect 503810 521056 503866 521112
rect 503534 471824 503590 471880
rect 503258 419056 503314 419112
rect 503442 341536 503498 341592
rect 503166 299376 503222 299432
rect 503074 192480 503130 192536
rect 503074 189760 503130 189816
rect 503074 186632 503130 186688
rect 503074 186496 503130 186552
rect 503074 180104 503130 180160
rect 503074 173032 503130 173088
rect 502982 166388 503038 166424
rect 502982 166368 502984 166388
rect 502984 166368 503036 166388
rect 503036 166368 503038 166388
rect 502982 165416 503038 165472
rect 502982 165008 503038 165064
rect 502982 163804 503038 163840
rect 502982 163784 502984 163804
rect 502984 163784 503036 163804
rect 503036 163784 503038 163804
rect 502982 162852 503038 162888
rect 502982 162832 502984 162852
rect 502984 162832 503036 162852
rect 503036 162832 503038 162852
rect 502982 162444 503038 162480
rect 502982 162424 502984 162444
rect 502984 162424 503036 162444
rect 503036 162424 503038 162444
rect 502982 162288 503038 162344
rect 502982 162016 503038 162072
rect 503258 271088 503314 271144
rect 503442 270544 503498 270600
rect 503350 270272 503406 270328
rect 503534 262384 503590 262440
rect 503442 260072 503498 260128
rect 503626 260208 503682 260264
rect 503350 259392 503406 259448
rect 503534 259528 503590 259584
rect 503534 258712 503590 258768
rect 503442 256672 503498 256728
rect 503534 256128 503590 256184
rect 503350 255312 503406 255368
rect 503626 255040 503682 255096
rect 503534 254904 503590 254960
rect 503350 254496 503406 254552
rect 503350 254088 503406 254144
rect 503442 253172 503444 253192
rect 503444 253172 503496 253192
rect 503496 253172 503498 253192
rect 503442 253136 503498 253172
rect 503442 253020 503498 253056
rect 503442 253000 503444 253020
rect 503444 253000 503496 253020
rect 503496 253000 503498 253020
rect 503442 246608 503498 246664
rect 503534 244160 503590 244216
rect 503534 243072 503590 243128
rect 503442 241440 503498 241496
rect 503442 239536 503498 239592
rect 503442 238040 503498 238096
rect 503350 229064 503406 229120
rect 503350 228928 503406 228984
rect 503534 237632 503590 237688
rect 503534 235728 503590 235784
rect 503534 235456 503590 235512
rect 503534 233144 503590 233200
rect 503442 225392 503498 225448
rect 503442 224848 503498 224904
rect 503442 221992 503498 222048
rect 503442 221876 503498 221912
rect 503442 221856 503444 221876
rect 503444 221856 503496 221876
rect 503496 221856 503498 221876
rect 503442 221448 503498 221504
rect 503626 226480 503682 226536
rect 503626 225120 503682 225176
rect 503626 220360 503682 220416
rect 503626 220244 503682 220280
rect 503626 220224 503628 220244
rect 503628 220224 503680 220244
rect 503680 220224 503682 220244
rect 503534 219816 503590 219872
rect 503626 216008 503682 216064
rect 503534 215872 503590 215928
rect 503534 215736 503590 215792
rect 503442 211792 503498 211848
rect 503442 211248 503498 211304
rect 503626 210740 503628 210760
rect 503628 210740 503680 210760
rect 503680 210740 503682 210760
rect 503626 210704 503682 210740
rect 503626 207712 503682 207768
rect 503534 204876 503590 204912
rect 503534 204856 503536 204876
rect 503536 204856 503588 204876
rect 503588 204856 503590 204876
rect 503534 204040 503590 204096
rect 503626 199316 503628 199336
rect 503628 199316 503680 199336
rect 503680 199316 503682 199336
rect 503626 199280 503682 199316
rect 503534 197376 503590 197432
rect 503626 196832 503682 196888
rect 503534 196188 503536 196208
rect 503536 196188 503588 196208
rect 503588 196188 503590 196208
rect 503534 196152 503590 196188
rect 503534 194404 503590 194440
rect 503534 194384 503536 194404
rect 503536 194384 503588 194404
rect 503588 194384 503590 194404
rect 503534 193568 503590 193624
rect 503626 186768 503682 186824
rect 503626 173168 503682 173224
rect 503626 173032 503682 173088
rect 503626 169088 503682 169144
rect 504178 500112 504234 500168
rect 503902 482432 503958 482488
rect 503810 185816 503866 185872
rect 503810 183504 503866 183560
rect 503810 180240 503866 180296
rect 503810 180140 503812 180160
rect 503812 180140 503864 180160
rect 503864 180140 503866 180160
rect 503810 180104 503866 180140
rect 503810 179424 503866 179480
rect 503718 147872 503774 147928
rect 503718 137264 503774 137320
rect 503718 134952 503774 135008
rect 503718 133900 503720 133920
rect 503720 133900 503772 133920
rect 503772 133900 503774 133920
rect 503718 133864 503774 133900
rect 503718 133728 503774 133784
rect 503718 130620 503774 130656
rect 503718 130600 503720 130620
rect 503720 130600 503772 130620
rect 503772 130600 503774 130620
rect 503626 130192 503682 130248
rect 503626 124888 503682 124944
rect 503718 123936 503774 123992
rect 503994 440272 504050 440328
rect 503902 165824 503958 165880
rect 503902 165572 503958 165608
rect 503902 165552 503904 165572
rect 503904 165552 503956 165572
rect 503956 165552 503958 165572
rect 503902 163648 503958 163704
rect 503902 161744 503958 161800
rect 503626 121352 503682 121408
rect 504086 436736 504142 436792
rect 504178 388320 504234 388376
rect 504270 380160 504326 380216
rect 504178 376896 504234 376952
rect 504178 373360 504234 373416
rect 504178 352144 504234 352200
rect 504178 345072 504234 345128
rect 504178 274660 504180 274680
rect 504180 274660 504232 274680
rect 504232 274660 504234 274680
rect 504178 274624 504234 274660
rect 504086 158752 504142 158808
rect 504086 158480 504142 158536
rect 503994 157392 504050 157448
rect 504086 154944 504142 155000
rect 504086 146140 504088 146160
rect 504088 146140 504140 146160
rect 504140 146140 504142 146160
rect 504086 146104 504142 146140
rect 504086 145988 504142 146024
rect 504086 145968 504088 145988
rect 504088 145968 504140 145988
rect 504140 145968 504142 145988
rect 504086 145832 504142 145888
rect 504086 144336 504142 144392
rect 503994 116048 504050 116104
rect 503994 87624 504050 87680
rect 503994 77288 504050 77344
rect 503994 49000 504050 49056
rect 503994 38800 504050 38856
rect 504914 581984 504970 582040
rect 505006 581576 505062 581632
rect 505190 581576 505246 581632
rect 504914 581168 504970 581224
rect 505006 581032 505062 581088
rect 504914 556144 504970 556200
rect 504822 552084 504878 552120
rect 504822 552064 504824 552084
rect 504824 552064 504876 552084
rect 504876 552064 504878 552084
rect 505006 549364 505062 549400
rect 505006 549344 505008 549364
rect 505008 549344 505060 549364
rect 505060 549344 505062 549364
rect 504454 534112 504510 534168
rect 505006 528128 505062 528184
rect 504454 524592 504510 524648
rect 504454 496576 504510 496632
rect 505006 492668 505008 492688
rect 505008 492668 505060 492688
rect 505060 492668 505062 492688
rect 505006 492632 505062 492668
rect 505006 478916 505062 478952
rect 505006 478896 505008 478916
rect 505008 478896 505060 478916
rect 505060 478896 505062 478916
rect 504546 454144 504602 454200
rect 504638 426128 504694 426184
rect 504546 390768 504602 390824
rect 504546 369860 504548 369880
rect 504548 369860 504600 369880
rect 504600 369860 504602 369880
rect 504546 369824 504602 369860
rect 504546 362788 504548 362808
rect 504548 362788 504600 362808
rect 504600 362788 504602 362808
rect 504546 362752 504602 362788
rect 504546 347520 504602 347576
rect 504546 338816 504602 338872
rect 504546 334464 504602 334520
rect 504454 330928 504510 330984
rect 504454 323856 504510 323912
rect 504454 309984 504510 310040
rect 504454 306448 504510 306504
rect 504454 295840 504510 295896
rect 504454 288768 504510 288824
rect 505006 404912 505062 404968
rect 504822 348608 504878 348664
rect 504730 307128 504786 307184
rect 504730 297336 504786 297392
rect 504730 281696 504786 281752
rect 504730 271768 504786 271824
rect 504730 267008 504786 267064
rect 504730 256944 504786 257000
rect 504638 246472 504694 246528
rect 504638 244704 504694 244760
rect 504638 236020 504694 236056
rect 504638 236000 504640 236020
rect 504640 236000 504692 236020
rect 504692 236000 504694 236020
rect 504546 147600 504602 147656
rect 504546 143928 504602 143984
rect 504546 143520 504602 143576
rect 504546 143404 504602 143440
rect 504546 143384 504548 143404
rect 504548 143384 504600 143404
rect 504600 143384 504602 143404
rect 504546 140800 504602 140856
rect 504546 118224 504602 118280
rect 504546 105984 504602 106040
rect 505006 292304 505062 292360
rect 504914 260480 504970 260536
rect 504822 197104 504878 197160
rect 504822 182960 504878 183016
rect 504270 80144 504326 80200
rect 504270 77288 504326 77344
rect 504454 49000 504510 49056
rect 504454 38664 504510 38720
rect 505006 172624 505062 172680
rect 505190 581032 505246 581088
rect 505190 489504 505246 489560
rect 505558 429664 505614 429720
rect 505650 411984 505706 412040
rect 506018 366288 506074 366344
rect 505834 253408 505890 253464
rect 506018 232464 506074 232520
rect 505834 178220 505890 178256
rect 505834 178200 505836 178220
rect 505836 178200 505888 178220
rect 505888 178200 505890 178220
rect 505834 152632 505890 152688
rect 505834 152108 505890 152144
rect 505834 152088 505836 152108
rect 505836 152088 505888 152108
rect 505888 152088 505890 152108
rect 505834 151852 505836 151872
rect 505836 151852 505888 151872
rect 505888 151852 505890 151872
rect 505834 151816 505890 151852
rect 505834 143384 505890 143440
rect 505834 139848 505890 139904
rect 506386 131960 506442 132016
rect 506662 580896 506718 580952
rect 507030 434560 507086 434616
rect 507030 425176 507086 425232
rect 507030 405592 507086 405648
rect 507030 396072 507086 396128
rect 507030 394576 507086 394632
rect 507030 387096 507086 387152
rect 506846 328344 506902 328400
rect 506846 323584 506902 323640
rect 507030 297336 507086 297392
rect 507030 280744 507086 280800
rect 507030 270680 507086 270736
rect 507030 242120 507086 242176
rect 507030 235320 507086 235376
rect 506938 218320 506994 218376
rect 506846 190032 506902 190088
rect 507030 204176 507086 204232
rect 507858 584024 507914 584080
rect 506662 119312 506718 119368
rect 507674 319504 507730 319560
rect 507674 318824 507730 318880
rect 507674 315968 507730 316024
rect 507674 249872 507730 249928
rect 507582 120536 507638 120592
rect 507490 119992 507546 120048
rect 507766 158072 507822 158128
rect 507766 143792 507822 143848
rect 508502 580624 508558 580680
rect 508410 121488 508466 121544
rect 508594 120944 508650 121000
rect 509238 584160 509294 584216
rect 508870 119720 508926 119776
rect 509054 214784 509110 214840
rect 507858 2760 507914 2816
rect 509974 581576 510030 581632
rect 509974 581168 510030 581224
rect 509974 580216 510030 580272
rect 509790 121760 509846 121816
rect 510434 246336 510490 246392
rect 510250 119040 510306 119096
rect 517518 584432 517574 584488
rect 511446 580080 511502 580136
rect 511354 119856 511410 119912
rect 512090 11600 512146 11656
rect 514666 545400 514722 545456
rect 514850 545264 514906 545320
rect 514666 181092 514668 181112
rect 514668 181092 514720 181112
rect 514720 181092 514722 181112
rect 514666 181056 514722 181092
rect 520278 584296 520334 584352
rect 523038 581304 523094 581360
rect 521566 181092 521568 181112
rect 521568 181092 521620 181112
rect 521620 181092 521622 181112
rect 521566 181056 521622 181092
rect 524418 570152 524474 570208
rect 524418 570016 524474 570072
rect 524326 545264 524382 545320
rect 524510 545128 524566 545184
rect 524418 278704 524474 278760
rect 524602 278704 524658 278760
rect 524418 259392 524474 259448
rect 524602 259392 524658 259448
rect 524418 241712 524474 241768
rect 524418 241576 524474 241632
rect 524418 240080 524474 240136
rect 524602 240080 524658 240136
rect 524418 220768 524474 220824
rect 524602 220768 524658 220824
rect 524418 211112 524474 211168
rect 524602 211112 524658 211168
rect 524418 191800 524474 191856
rect 524602 191800 524658 191856
rect 524418 172488 524474 172544
rect 524602 172488 524658 172544
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 542358 584976 542414 585032
rect 532698 578176 532754 578232
rect 532882 578176 532938 578232
rect 532422 568520 532478 568576
rect 532698 568556 532700 568576
rect 532700 568556 532752 568576
rect 532752 568556 532754 568576
rect 532698 568520 532754 568556
rect 531962 545400 532018 545456
rect 529938 545164 529940 545184
rect 529940 545164 529992 545184
rect 529992 545164 529994 545184
rect 529938 545128 529994 545164
rect 532698 531256 532754 531312
rect 532882 531256 532938 531312
rect 532698 511944 532754 512000
rect 532882 511944 532938 512000
rect 532698 482976 532754 483032
rect 532882 482976 532938 483032
rect 529938 238876 529994 238912
rect 529938 238856 529940 238876
rect 529940 238856 529992 238876
rect 529992 238856 529994 238876
rect 529938 116592 529994 116648
rect 532698 183504 532754 183560
rect 532882 183504 532938 183560
rect 533986 180956 533988 180976
rect 533988 180956 534040 180976
rect 534040 180956 534042 180976
rect 533986 180920 534042 180956
rect 532698 172488 532754 172544
rect 532882 172488 532938 172544
rect 535458 180956 535460 180976
rect 535460 180956 535512 180976
rect 535512 180956 535514 180976
rect 535458 180920 535514 180956
rect 535734 6296 535790 6352
rect 538218 12960 538274 13016
rect 539506 238856 539562 238912
rect 540334 119448 540390 119504
rect 546498 584568 546554 584624
rect 553398 14456 553454 14512
rect 580262 583888 580318 583944
rect 558918 581032 558974 581088
rect 558366 3712 558422 3768
rect 579618 582120 579674 582176
rect 560298 15816 560354 15872
rect 561954 6160 562010 6216
rect 563150 116456 563206 116512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 579986 498616 580042 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 579986 439864 580042 439920
rect 580170 416472 580226 416528
rect 579710 392944 579766 393000
rect 580170 369552 580226 369608
rect 580170 346024 580226 346080
rect 580170 322632 580226 322688
rect 580170 299104 580226 299160
rect 580170 275712 580226 275768
rect 580170 252184 580226 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 580170 205264 580226 205320
rect 579710 181872 579766 181928
rect 579710 181056 579766 181112
rect 580170 170040 580226 170096
rect 580170 158344 580226 158400
rect 580170 123120 580226 123176
rect 580170 76200 580226 76256
rect 580170 64504 580226 64560
rect 580170 40976 580226 41032
rect 580446 451696 580502 451752
rect 580446 404776 580502 404832
rect 580630 357856 580686 357912
rect 580538 310800 580594 310856
rect 580354 111424 580410 111480
rect 580262 17584 580318 17640
<< metal3 >>
rect 92238 700708 92244 700772
rect 92308 700770 92314 700772
rect 154113 700770 154179 700773
rect 92308 700768 154179 700770
rect 92308 700712 154118 700768
rect 154174 700712 154179 700768
rect 92308 700710 154179 700712
rect 92308 700708 92314 700710
rect 154113 700707 154179 700710
rect 89478 700572 89484 700636
rect 89548 700634 89554 700636
rect 218973 700634 219039 700637
rect 89548 700632 219039 700634
rect 89548 700576 218978 700632
rect 219034 700576 219039 700632
rect 89548 700574 219039 700576
rect 89548 700572 89554 700574
rect 218973 700571 219039 700574
rect 93342 700436 93348 700500
rect 93412 700498 93418 700500
rect 267641 700498 267707 700501
rect 93412 700496 267707 700498
rect 93412 700440 267646 700496
rect 267702 700440 267707 700496
rect 93412 700438 267707 700440
rect 93412 700436 93418 700438
rect 267641 700435 267707 700438
rect 91870 700300 91876 700364
rect 91940 700362 91946 700364
rect 348785 700362 348851 700365
rect 91940 700360 348851 700362
rect 91940 700304 348790 700360
rect 348846 700304 348851 700360
rect 91940 700302 348851 700304
rect 91940 700300 91946 700302
rect 348785 700299 348851 700302
rect 89161 699818 89227 699821
rect 90214 699818 90220 699820
rect 89161 699816 90220 699818
rect 89161 699760 89166 699816
rect 89222 699760 90220 699816
rect 89161 699758 90220 699760
rect 89161 699755 89227 699758
rect 90214 699756 90220 699758
rect 90284 699756 90290 699820
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 518942 697174 528570 697234
rect 505686 696900 505692 696964
rect 505756 696962 505762 696964
rect 518942 696962 519002 697174
rect 528510 697098 528570 697174
rect 538262 697174 547890 697234
rect 528510 697038 538138 697098
rect 505756 696902 519002 696962
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 547830 697098 547890 697174
rect 557582 697174 567210 697234
rect 547830 697038 557458 697098
rect 538078 696902 538322 696962
rect 557398 696962 557458 697038
rect 557582 696962 557642 697174
rect 567150 697098 567210 697174
rect 567150 697038 576778 697098
rect 557398 696902 557642 696962
rect 576718 696962 576778 697038
rect 583342 696962 583402 697990
rect 583520 697900 584960 697990
rect 576718 696902 583402 696962
rect 505756 696900 505762 696902
rect -960 696540 480 696780
rect 89529 695468 89595 695469
rect 89478 695404 89484 695468
rect 89548 695466 89595 695468
rect 89548 695464 89640 695466
rect 89590 695408 89640 695464
rect 89548 695406 89640 695408
rect 89548 695404 89595 695406
rect 89529 695403 89595 695404
rect 89529 689346 89595 689349
rect 89846 689346 89852 689348
rect 89529 689344 89852 689346
rect 89529 689288 89534 689344
rect 89590 689288 89852 689344
rect 89529 689286 89852 689288
rect 89529 689283 89595 689286
rect 89846 689284 89852 689286
rect 89916 689284 89922 689348
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 89529 674796 89595 674797
rect 89478 674732 89484 674796
rect 89548 674794 89595 674796
rect 89548 674792 89640 674794
rect 89590 674736 89640 674792
rect 89548 674734 89640 674736
rect 89548 674732 89595 674734
rect 89529 674731 89595 674732
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 89529 665276 89595 665277
rect 89478 665274 89484 665276
rect 89438 665214 89484 665274
rect 89548 665272 89595 665276
rect 89590 665216 89595 665272
rect 89478 665212 89484 665214
rect 89548 665212 89595 665216
rect 89529 665211 89595 665212
rect 583520 662676 584960 662916
rect 89529 655484 89595 655485
rect 89478 655420 89484 655484
rect 89548 655482 89595 655484
rect 89548 655480 89640 655482
rect 89590 655424 89640 655480
rect 89548 655422 89640 655424
rect 89548 655420 89595 655422
rect 89529 655419 89595 655420
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 89529 645964 89595 645965
rect 89478 645962 89484 645964
rect 89438 645902 89484 645962
rect 89548 645960 89595 645964
rect 89590 645904 89595 645960
rect 89478 645900 89484 645902
rect 89548 645900 89595 645904
rect 89529 645899 89595 645900
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 89529 636172 89595 636173
rect 89478 636108 89484 636172
rect 89548 636170 89595 636172
rect 89548 636168 89640 636170
rect 89590 636112 89640 636168
rect 89548 636110 89640 636112
rect 89548 636108 89595 636110
rect 89529 636107 89595 636108
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect 89529 626652 89595 626653
rect 89478 626650 89484 626652
rect 89438 626590 89484 626650
rect 89548 626648 89595 626652
rect 89590 626592 89595 626648
rect 89478 626588 89484 626590
rect 89548 626588 89595 626592
rect 89529 626587 89595 626588
rect 89294 626452 89300 626516
rect 89364 626514 89370 626516
rect 89478 626514 89484 626516
rect 89364 626454 89484 626514
rect 89364 626452 89370 626454
rect 89478 626452 89484 626454
rect 89548 626452 89554 626516
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 83549 597546 83615 597549
rect 83733 597546 83799 597549
rect 83549 597544 83799 597546
rect 83549 597488 83554 597544
rect 83610 597488 83738 597544
rect 83794 597488 83799 597544
rect 83549 597486 83799 597488
rect 83549 597483 83615 597486
rect 83733 597483 83799 597486
rect 89437 596188 89503 596189
rect 89437 596186 89484 596188
rect 89392 596184 89484 596186
rect -960 596050 480 596140
rect 89392 596128 89442 596184
rect 89392 596126 89484 596128
rect 89437 596124 89484 596126
rect 89548 596124 89554 596188
rect 89437 596123 89503 596124
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 87638 585652 87644 585716
rect 87708 585714 87714 585716
rect 412909 585714 412975 585717
rect 87708 585712 412975 585714
rect 87708 585656 412914 585712
rect 412970 585656 412975 585712
rect 87708 585654 412975 585656
rect 87708 585652 87714 585654
rect 412909 585651 412975 585654
rect 99238 585246 99482 585306
rect 89662 584972 89668 585036
rect 89732 585034 89738 585036
rect 99238 585034 99298 585246
rect 99422 585170 99482 585246
rect 99422 585110 148978 585170
rect 89732 584974 99298 585034
rect 89732 584972 89738 584974
rect 88190 584836 88196 584900
rect 88260 584898 88266 584900
rect 148777 584898 148843 584901
rect 88260 584896 148843 584898
rect 88260 584840 148782 584896
rect 148838 584840 148843 584896
rect 88260 584838 148843 584840
rect 148918 584898 148978 585110
rect 205633 585034 205699 585037
rect 225137 585034 225203 585037
rect 542353 585034 542419 585037
rect 195654 584974 198106 585034
rect 157241 584898 157307 584901
rect 148918 584896 157307 584898
rect 148918 584840 157246 584896
rect 157302 584840 157307 584896
rect 148918 584838 157307 584840
rect 88260 584836 88266 584838
rect 148777 584835 148843 584838
rect 157241 584835 157307 584838
rect 157425 584898 157491 584901
rect 172462 584898 172468 584900
rect 157425 584896 172468 584898
rect 157425 584840 157430 584896
rect 157486 584840 172468 584896
rect 157425 584838 172468 584840
rect 157425 584835 157491 584838
rect 172462 584836 172468 584838
rect 172532 584836 172538 584900
rect 191741 584898 191807 584901
rect 195654 584898 195714 584974
rect 191741 584896 195714 584898
rect 191741 584840 191746 584896
rect 191802 584840 195714 584896
rect 191741 584838 195714 584840
rect 198046 584898 198106 584974
rect 205633 585032 206938 585034
rect 205633 584976 205638 585032
rect 205694 584976 206938 585032
rect 205633 584974 206938 584976
rect 205633 584971 205699 584974
rect 205541 584898 205607 584901
rect 198046 584896 205607 584898
rect 198046 584840 205546 584896
rect 205602 584840 205607 584896
rect 198046 584838 205607 584840
rect 206878 584898 206938 584974
rect 207062 584974 215402 585034
rect 207062 584898 207122 584974
rect 206878 584838 207122 584898
rect 191741 584835 191807 584838
rect 205541 584835 205607 584838
rect 91686 584700 91692 584764
rect 91756 584762 91762 584764
rect 158345 584762 158411 584765
rect 91756 584760 158411 584762
rect 91756 584704 158350 584760
rect 158406 584704 158411 584760
rect 91756 584702 158411 584704
rect 91756 584700 91762 584702
rect 158345 584699 158411 584702
rect 172646 584700 172652 584764
rect 172716 584762 172722 584764
rect 182173 584762 182239 584765
rect 172716 584760 182239 584762
rect 172716 584704 182178 584760
rect 182234 584704 182239 584760
rect 172716 584702 182239 584704
rect 215342 584762 215402 584974
rect 225137 585032 542419 585034
rect 225137 584976 225142 585032
rect 225198 584976 542358 585032
rect 542414 584976 542419 585032
rect 225137 584974 542419 584976
rect 225137 584971 225203 584974
rect 542353 584971 542419 584974
rect 218145 584898 218211 584901
rect 227713 584898 227779 584901
rect 218145 584896 227779 584898
rect 218145 584840 218150 584896
rect 218206 584840 227718 584896
rect 227774 584840 227779 584896
rect 218145 584838 227779 584840
rect 218145 584835 218211 584838
rect 227713 584835 227779 584838
rect 427537 584898 427603 584901
rect 501638 584898 501644 584900
rect 427537 584896 501644 584898
rect 427537 584840 427542 584896
rect 427598 584840 501644 584896
rect 427537 584838 501644 584840
rect 427537 584835 427603 584838
rect 501638 584836 501644 584838
rect 501708 584836 501714 584900
rect 218053 584762 218119 584765
rect 215342 584760 218119 584762
rect 215342 584704 218058 584760
rect 218114 584704 218119 584760
rect 215342 584702 218119 584704
rect 172716 584700 172722 584702
rect 182173 584699 182239 584702
rect 218053 584699 218119 584702
rect 234521 584762 234587 584765
rect 238753 584762 238819 584765
rect 234521 584760 238819 584762
rect 234521 584704 234526 584760
rect 234582 584704 238758 584760
rect 238814 584704 238819 584760
rect 234521 584702 238819 584704
rect 234521 584699 234587 584702
rect 238753 584699 238819 584702
rect 372613 584762 372679 584765
rect 465625 584762 465691 584765
rect 372613 584760 465691 584762
rect 372613 584704 372618 584760
rect 372674 584704 465630 584760
rect 465686 584704 465691 584760
rect 372613 584702 465691 584704
rect 372613 584699 372679 584702
rect 465625 584699 465691 584702
rect 472801 584762 472867 584765
rect 506238 584762 506244 584764
rect 472801 584760 506244 584762
rect 472801 584704 472806 584760
rect 472862 584704 506244 584760
rect 472801 584702 506244 584704
rect 472801 584699 472867 584702
rect 506238 584700 506244 584702
rect 506308 584700 506314 584764
rect 88374 584564 88380 584628
rect 88444 584626 88450 584628
rect 291745 584626 291811 584629
rect 88444 584624 291811 584626
rect 88444 584568 291750 584624
rect 291806 584568 291811 584624
rect 88444 584566 291811 584568
rect 88444 584564 88450 584566
rect 291745 584563 291811 584566
rect 315665 584626 315731 584629
rect 546493 584626 546559 584629
rect 315665 584624 546559 584626
rect 315665 584568 315670 584624
rect 315726 584568 546498 584624
rect 546554 584568 546559 584624
rect 315665 584566 546559 584568
rect 315665 584563 315731 584566
rect 546493 584563 546559 584566
rect 97758 584428 97764 584492
rect 97828 584490 97834 584492
rect 182265 584490 182331 584493
rect 97828 584488 182331 584490
rect 97828 584432 182270 584488
rect 182326 584432 182331 584488
rect 97828 584430 182331 584432
rect 97828 584428 97834 584430
rect 182265 584427 182331 584430
rect 233233 584490 233299 584493
rect 233918 584490 233924 584492
rect 233233 584488 233924 584490
rect 233233 584432 233238 584488
rect 233294 584432 233924 584488
rect 233233 584430 233924 584432
rect 233233 584427 233299 584430
rect 233918 584428 233924 584430
rect 233988 584428 233994 584492
rect 275001 584490 275067 584493
rect 517513 584490 517579 584493
rect 275001 584488 517579 584490
rect 275001 584432 275006 584488
rect 275062 584432 517518 584488
rect 517574 584432 517579 584488
rect 275001 584430 517579 584432
rect 275001 584427 275067 584430
rect 517513 584427 517579 584430
rect 87270 584292 87276 584356
rect 87340 584354 87346 584356
rect 175089 584354 175155 584357
rect 87340 584352 175155 584354
rect 87340 584296 175094 584352
rect 175150 584296 175155 584352
rect 87340 584294 175155 584296
rect 87340 584292 87346 584294
rect 175089 584291 175155 584294
rect 277393 584354 277459 584357
rect 520273 584354 520339 584357
rect 277393 584352 520339 584354
rect 277393 584296 277398 584352
rect 277454 584296 520278 584352
rect 520334 584296 520339 584352
rect 277393 584294 520339 584296
rect 277393 584291 277459 584294
rect 520273 584291 520339 584294
rect 88558 584156 88564 584220
rect 88628 584218 88634 584220
rect 241697 584218 241763 584221
rect 88628 584216 241763 584218
rect 88628 584160 241702 584216
rect 241758 584160 241763 584216
rect 88628 584158 241763 584160
rect 88628 584156 88634 584158
rect 241697 584155 241763 584158
rect 258441 584218 258507 584221
rect 509233 584218 509299 584221
rect 258441 584216 509299 584218
rect 258441 584160 258446 584216
rect 258502 584160 509238 584216
rect 509294 584160 509299 584216
rect 258441 584158 509299 584160
rect 258441 584155 258507 584158
rect 509233 584155 509299 584158
rect 92606 584020 92612 584084
rect 92676 584082 92682 584084
rect 201217 584082 201283 584085
rect 92676 584080 201283 584082
rect 92676 584024 201222 584080
rect 201278 584024 201283 584080
rect 92676 584022 201283 584024
rect 92676 584020 92682 584022
rect 201217 584019 201283 584022
rect 222745 584082 222811 584085
rect 507853 584082 507919 584085
rect 222745 584080 507919 584082
rect 222745 584024 222750 584080
rect 222806 584024 507858 584080
rect 507914 584024 507919 584080
rect 222745 584022 507919 584024
rect 222745 584019 222811 584022
rect 507853 584019 507919 584022
rect 84510 583884 84516 583948
rect 84580 583946 84586 583948
rect 179873 583946 179939 583949
rect 84580 583944 179939 583946
rect 84580 583888 179878 583944
rect 179934 583888 179939 583944
rect 84580 583886 179939 583888
rect 84580 583884 84586 583886
rect 179873 583883 179939 583886
rect 186865 583946 186931 583949
rect 494605 583946 494671 583949
rect 186865 583944 494671 583946
rect 186865 583888 186870 583944
rect 186926 583888 494610 583944
rect 494666 583888 494671 583944
rect 186865 583886 494671 583888
rect 186865 583883 186931 583886
rect 494605 583883 494671 583886
rect 496721 583946 496787 583949
rect 496721 583944 499314 583946
rect 496721 583888 496726 583944
rect 496782 583888 499314 583944
rect 496721 583886 499314 583888
rect 496721 583883 496787 583886
rect 92105 583812 92171 583813
rect 92054 583810 92060 583812
rect 92014 583750 92060 583810
rect 92124 583808 92171 583812
rect 92166 583752 92171 583808
rect 92054 583748 92060 583750
rect 92124 583748 92171 583752
rect 93526 583748 93532 583812
rect 93596 583810 93602 583812
rect 139209 583810 139275 583813
rect 93596 583808 139275 583810
rect 93596 583752 139214 583808
rect 139270 583752 139275 583808
rect 93596 583750 139275 583752
rect 93596 583748 93602 583750
rect 92105 583747 92171 583748
rect 139209 583747 139275 583750
rect 233182 583748 233188 583812
rect 233252 583810 233258 583812
rect 234521 583810 234587 583813
rect 233252 583808 234587 583810
rect 233252 583752 234526 583808
rect 234582 583752 234587 583808
rect 233252 583750 234587 583752
rect 233252 583748 233258 583750
rect 234521 583747 234587 583750
rect 298134 583748 298140 583812
rect 298204 583810 298210 583812
rect 298921 583810 298987 583813
rect 298204 583808 298987 583810
rect 298204 583752 298926 583808
rect 298982 583752 298987 583808
rect 298204 583750 298987 583752
rect 298204 583748 298210 583750
rect 298921 583747 298987 583750
rect 451457 583810 451523 583813
rect 499062 583810 499068 583812
rect 451457 583808 499068 583810
rect 451457 583752 451462 583808
rect 451518 583752 499068 583808
rect 451457 583750 499068 583752
rect 451457 583747 451523 583750
rect 499062 583748 499068 583750
rect 499132 583748 499138 583812
rect 499254 583810 499314 583886
rect 499430 583884 499436 583948
rect 499500 583946 499506 583948
rect 580257 583946 580323 583949
rect 499500 583944 580323 583946
rect 499500 583888 580262 583944
rect 580318 583888 580323 583944
rect 499500 583886 580323 583888
rect 499500 583884 499506 583886
rect 580257 583883 580323 583886
rect 509366 583810 509372 583812
rect 499254 583750 509372 583810
rect 509366 583748 509372 583750
rect 509436 583748 509442 583812
rect 84694 582932 84700 582996
rect 84764 582994 84770 582996
rect 303705 582994 303771 582997
rect 84764 582992 303771 582994
rect 84764 582936 303710 582992
rect 303766 582936 303771 582992
rect 84764 582934 303771 582936
rect 84764 582932 84770 582934
rect 303705 582931 303771 582934
rect 314653 582994 314719 582997
rect 500350 582994 500356 582996
rect 314653 582992 500356 582994
rect 314653 582936 314658 582992
rect 314714 582936 500356 582992
rect 314653 582934 500356 582936
rect 314653 582931 314719 582934
rect 500350 582932 500356 582934
rect 500420 582932 500426 582996
rect 89345 582858 89411 582861
rect 89478 582858 89484 582860
rect 89345 582856 89484 582858
rect 89345 582800 89350 582856
rect 89406 582800 89484 582856
rect 89345 582798 89484 582800
rect 89345 582795 89411 582798
rect 89478 582796 89484 582798
rect 89548 582796 89554 582860
rect 106038 582796 106044 582860
rect 106108 582858 106114 582860
rect 213177 582858 213243 582861
rect 106108 582856 213243 582858
rect 106108 582800 213182 582856
rect 213238 582800 213243 582856
rect 106108 582798 213243 582800
rect 106108 582796 106114 582798
rect 213177 582795 213243 582798
rect 318057 582858 318123 582861
rect 502701 582858 502767 582861
rect 318057 582856 502767 582858
rect 318057 582800 318062 582856
rect 318118 582800 502706 582856
rect 502762 582800 502767 582856
rect 318057 582798 502767 582800
rect 318057 582795 318123 582798
rect 502701 582795 502767 582798
rect 301313 582722 301379 582725
rect 501270 582722 501276 582724
rect 301313 582720 501276 582722
rect 301313 582664 301318 582720
rect 301374 582664 501276 582720
rect 301313 582662 501276 582664
rect 301313 582659 301379 582662
rect 501270 582660 501276 582662
rect 501340 582660 501346 582724
rect 206001 582586 206067 582589
rect 506054 582586 506060 582588
rect 206001 582584 506060 582586
rect 206001 582528 206006 582584
rect 206062 582528 506060 582584
rect 206001 582526 506060 582528
rect 206001 582523 206067 582526
rect 506054 582524 506060 582526
rect 506124 582524 506130 582588
rect 86718 582388 86724 582452
rect 86788 582450 86794 582452
rect 94221 582450 94287 582453
rect 101305 582450 101371 582453
rect 107653 582450 107719 582453
rect 86788 582390 93962 582450
rect 86788 582388 86794 582390
rect 89069 582314 89135 582317
rect 93669 582314 93735 582317
rect 89069 582312 93735 582314
rect 89069 582256 89074 582312
rect 89130 582256 93674 582312
rect 93730 582256 93735 582312
rect 89069 582254 93735 582256
rect 89069 582251 89135 582254
rect 93669 582251 93735 582254
rect 89110 582116 89116 582180
rect 89180 582178 89186 582180
rect 93761 582178 93827 582181
rect 89180 582176 93827 582178
rect 89180 582120 93766 582176
rect 93822 582120 93827 582176
rect 89180 582118 93827 582120
rect 93902 582178 93962 582390
rect 94221 582448 101371 582450
rect 94221 582392 94226 582448
rect 94282 582392 101310 582448
rect 101366 582392 101371 582448
rect 94221 582390 101371 582392
rect 94221 582387 94287 582390
rect 101305 582387 101371 582390
rect 101446 582448 107719 582450
rect 101446 582392 107658 582448
rect 107714 582392 107719 582448
rect 101446 582390 107719 582392
rect 94129 582314 94195 582317
rect 101446 582314 101506 582390
rect 107653 582387 107719 582390
rect 113265 582450 113331 582453
rect 132493 582450 132559 582453
rect 156321 582450 156387 582453
rect 113265 582448 115674 582450
rect 113265 582392 113270 582448
rect 113326 582392 115674 582448
rect 113265 582390 115674 582392
rect 113265 582387 113331 582390
rect 94129 582312 101506 582314
rect 94129 582256 94134 582312
rect 94190 582256 101506 582312
rect 94129 582254 101506 582256
rect 101581 582314 101647 582317
rect 113766 582314 113772 582316
rect 101581 582312 113772 582314
rect 101581 582256 101586 582312
rect 101642 582256 113772 582312
rect 101581 582254 113772 582256
rect 94129 582251 94195 582254
rect 101581 582251 101647 582254
rect 113766 582252 113772 582254
rect 113836 582252 113842 582316
rect 115614 582314 115674 582390
rect 132493 582448 133154 582450
rect 132493 582392 132498 582448
rect 132554 582392 133154 582448
rect 132493 582390 133154 582392
rect 132493 582387 132559 582390
rect 123477 582314 123543 582317
rect 115614 582312 123543 582314
rect 115614 582256 123482 582312
rect 123538 582256 123543 582312
rect 115614 582254 123543 582256
rect 123477 582251 123543 582254
rect 123753 582314 123819 582317
rect 132953 582314 133019 582317
rect 123753 582312 133019 582314
rect 123753 582256 123758 582312
rect 123814 582256 132958 582312
rect 133014 582256 133019 582312
rect 123753 582254 133019 582256
rect 133094 582314 133154 582390
rect 153334 582448 156387 582450
rect 153334 582392 156326 582448
rect 156382 582392 156387 582448
rect 153334 582390 156387 582392
rect 142797 582314 142863 582317
rect 133094 582312 142863 582314
rect 133094 582256 142802 582312
rect 142858 582256 142863 582312
rect 133094 582254 142863 582256
rect 123753 582251 123819 582254
rect 132953 582251 133019 582254
rect 142797 582251 142863 582254
rect 147673 582314 147739 582317
rect 150985 582314 151051 582317
rect 147673 582312 151051 582314
rect 147673 582256 147678 582312
rect 147734 582256 150990 582312
rect 151046 582256 151051 582312
rect 147673 582254 151051 582256
rect 147673 582251 147739 582254
rect 150985 582251 151051 582254
rect 151169 582314 151235 582317
rect 153334 582314 153394 582390
rect 156321 582387 156387 582390
rect 196433 582450 196499 582453
rect 505870 582450 505876 582452
rect 196433 582448 505876 582450
rect 196433 582392 196438 582448
rect 196494 582392 505876 582448
rect 196433 582390 505876 582392
rect 196433 582387 196499 582390
rect 505870 582388 505876 582390
rect 505940 582388 505946 582452
rect 151169 582312 153394 582314
rect 151169 582256 151174 582312
rect 151230 582256 153394 582312
rect 151169 582254 153394 582256
rect 156597 582314 156663 582317
rect 162342 582314 162348 582316
rect 156597 582312 162348 582314
rect 156597 582256 156602 582312
rect 156658 582256 162348 582312
rect 156597 582254 162348 582256
rect 151169 582251 151235 582254
rect 156597 582251 156663 582254
rect 162342 582252 162348 582254
rect 162412 582252 162418 582316
rect 162485 582314 162551 582317
rect 166809 582314 166875 582317
rect 162485 582312 166875 582314
rect 162485 582256 162490 582312
rect 162546 582256 166814 582312
rect 166870 582256 166875 582312
rect 162485 582254 166875 582256
rect 162485 582251 162551 582254
rect 166809 582251 166875 582254
rect 166993 582314 167059 582317
rect 171593 582314 171659 582317
rect 166993 582312 171659 582314
rect 166993 582256 166998 582312
rect 167054 582256 171598 582312
rect 171654 582256 171659 582312
rect 166993 582254 171659 582256
rect 166993 582251 167059 582254
rect 171593 582251 171659 582254
rect 171777 582314 171843 582317
rect 181437 582314 181503 582317
rect 171777 582312 181503 582314
rect 171777 582256 171782 582312
rect 171838 582256 181442 582312
rect 181498 582256 181503 582312
rect 171777 582254 181503 582256
rect 171777 582251 171843 582254
rect 181437 582251 181503 582254
rect 181662 582252 181668 582316
rect 181732 582314 181738 582316
rect 190678 582314 190684 582316
rect 181732 582254 190684 582314
rect 181732 582252 181738 582254
rect 190678 582252 190684 582254
rect 190748 582252 190754 582316
rect 190821 582314 190887 582317
rect 200757 582314 200823 582317
rect 190821 582312 200823 582314
rect 190821 582256 190826 582312
rect 190882 582256 200762 582312
rect 200818 582256 200823 582312
rect 190821 582254 200823 582256
rect 190821 582251 190887 582254
rect 200757 582251 200823 582254
rect 200982 582252 200988 582316
rect 201052 582314 201058 582316
rect 211153 582314 211219 582317
rect 201052 582312 211219 582314
rect 201052 582256 211158 582312
rect 211214 582256 211219 582312
rect 201052 582254 211219 582256
rect 201052 582252 201058 582254
rect 211153 582251 211219 582254
rect 282913 582314 282979 582317
rect 292481 582314 292547 582317
rect 282913 582312 292547 582314
rect 282913 582256 282918 582312
rect 282974 582256 292486 582312
rect 292542 582256 292547 582312
rect 282913 582254 292547 582256
rect 282913 582251 282979 582254
rect 292481 582251 292547 582254
rect 302233 582314 302299 582317
rect 311801 582314 311867 582317
rect 302233 582312 311867 582314
rect 302233 582256 302238 582312
rect 302294 582256 311806 582312
rect 311862 582256 311867 582312
rect 302233 582254 311867 582256
rect 302233 582251 302299 582254
rect 311801 582251 311867 582254
rect 316534 582252 316540 582316
rect 316604 582314 316610 582316
rect 326470 582314 326476 582316
rect 316604 582254 326476 582314
rect 316604 582252 316610 582254
rect 326470 582252 326476 582254
rect 326540 582252 326546 582316
rect 412766 582252 412772 582316
rect 412836 582314 412842 582316
rect 423070 582314 423076 582316
rect 412836 582254 423076 582314
rect 412836 582252 412842 582254
rect 423070 582252 423076 582254
rect 423140 582252 423146 582316
rect 431902 582252 431908 582316
rect 431972 582314 431978 582316
rect 442206 582314 442212 582316
rect 431972 582254 442212 582314
rect 431972 582252 431978 582254
rect 442206 582252 442212 582254
rect 442276 582252 442282 582316
rect 451958 582252 451964 582316
rect 452028 582314 452034 582316
rect 461342 582314 461348 582316
rect 452028 582254 461348 582314
rect 452028 582252 452034 582254
rect 461342 582252 461348 582254
rect 461412 582252 461418 582316
rect 470542 582252 470548 582316
rect 470612 582314 470618 582316
rect 480846 582314 480852 582316
rect 470612 582254 480852 582314
rect 470612 582252 470618 582254
rect 480846 582252 480852 582254
rect 480916 582252 480922 582316
rect 489862 582252 489868 582316
rect 489932 582314 489938 582316
rect 490189 582314 490255 582317
rect 489932 582312 490255 582314
rect 489932 582256 490194 582312
rect 490250 582256 490255 582312
rect 489932 582254 490255 582256
rect 489932 582252 489938 582254
rect 490189 582251 490255 582254
rect 490373 582314 490439 582317
rect 510654 582314 510660 582316
rect 490373 582312 510660 582314
rect 490373 582256 490378 582312
rect 490434 582256 510660 582312
rect 490373 582254 510660 582256
rect 490373 582251 490439 582254
rect 510654 582252 510660 582254
rect 510724 582252 510730 582316
rect 191649 582178 191715 582181
rect 93902 582176 191715 582178
rect 93902 582120 191654 582176
rect 191710 582120 191715 582176
rect 93902 582118 191715 582120
rect 89180 582116 89186 582118
rect 93761 582115 93827 582118
rect 191649 582115 191715 582118
rect 192017 582178 192083 582181
rect 200665 582178 200731 582181
rect 192017 582176 200731 582178
rect 192017 582120 192022 582176
rect 192078 582120 200670 582176
rect 200726 582120 200731 582176
rect 192017 582118 200731 582120
rect 192017 582115 192083 582118
rect 200665 582115 200731 582118
rect 200849 582178 200915 582181
rect 210366 582178 210372 582180
rect 200849 582176 210372 582178
rect 200849 582120 200854 582176
rect 200910 582120 210372 582176
rect 200849 582118 210372 582120
rect 200849 582115 200915 582118
rect 210366 582116 210372 582118
rect 210436 582116 210442 582180
rect 229369 582178 229435 582181
rect 258349 582178 258415 582181
rect 229369 582176 258415 582178
rect 229369 582120 229374 582176
rect 229430 582120 258354 582176
rect 258410 582120 258415 582176
rect 229369 582118 258415 582120
rect 229369 582115 229435 582118
rect 258349 582115 258415 582118
rect 260782 582116 260788 582180
rect 260852 582178 260858 582180
rect 273161 582178 273227 582181
rect 260852 582176 273227 582178
rect 260852 582120 273166 582176
rect 273222 582120 273227 582176
rect 260852 582118 273227 582120
rect 260852 582116 260858 582118
rect 273161 582115 273227 582118
rect 277526 582116 277532 582180
rect 277596 582178 277602 582180
rect 287830 582178 287836 582180
rect 277596 582118 287836 582178
rect 277596 582116 277602 582118
rect 287830 582116 287836 582118
rect 287900 582116 287906 582180
rect 297214 582116 297220 582180
rect 297284 582178 297290 582180
rect 306598 582178 306604 582180
rect 297284 582118 306604 582178
rect 297284 582116 297290 582118
rect 306598 582116 306604 582118
rect 306668 582116 306674 582180
rect 316718 582116 316724 582180
rect 316788 582178 316794 582180
rect 326286 582178 326292 582180
rect 316788 582118 326292 582178
rect 316788 582116 316794 582118
rect 326286 582116 326292 582118
rect 326356 582116 326362 582180
rect 326429 582178 326495 582181
rect 329833 582178 329899 582181
rect 326429 582176 329899 582178
rect 326429 582120 326434 582176
rect 326490 582120 329838 582176
rect 329894 582120 329899 582176
rect 326429 582118 329899 582120
rect 326429 582115 326495 582118
rect 329833 582115 329899 582118
rect 393446 582116 393452 582180
rect 393516 582178 393522 582180
rect 403750 582178 403756 582180
rect 393516 582118 403756 582178
rect 393516 582116 393522 582118
rect 403750 582116 403756 582118
rect 403820 582116 403826 582180
rect 412582 582116 412588 582180
rect 412652 582178 412658 582180
rect 422886 582178 422892 582180
rect 412652 582118 422892 582178
rect 412652 582116 412658 582118
rect 422886 582116 422892 582118
rect 422956 582116 422962 582180
rect 424961 582178 425027 582181
rect 491702 582178 491708 582180
rect 424961 582176 491708 582178
rect 424961 582120 424966 582176
rect 425022 582120 491708 582176
rect 424961 582118 491708 582120
rect 424961 582115 425027 582118
rect 491702 582116 491708 582118
rect 491772 582116 491778 582180
rect 491845 582178 491911 582181
rect 579613 582178 579679 582181
rect 491845 582176 579679 582178
rect 491845 582120 491850 582176
rect 491906 582120 579618 582176
rect 579674 582120 579679 582176
rect 491845 582118 579679 582120
rect 491845 582115 491911 582118
rect 579613 582115 579679 582118
rect 85246 581980 85252 582044
rect 85316 582042 85322 582044
rect 89713 582042 89779 582045
rect 85316 582040 89779 582042
rect 85316 581984 89718 582040
rect 89774 581984 89779 582040
rect 85316 581982 89779 581984
rect 85316 581980 85322 581982
rect 89713 581979 89779 581982
rect 89846 581980 89852 582044
rect 89916 582042 89922 582044
rect 93393 582042 93459 582045
rect 89916 582040 93459 582042
rect 89916 581984 93398 582040
rect 93454 581984 93459 582040
rect 89916 581982 93459 581984
rect 89916 581980 89922 581982
rect 93393 581979 93459 581982
rect 118601 582042 118667 582045
rect 128353 582042 128419 582045
rect 118601 582040 128419 582042
rect 118601 581984 118606 582040
rect 118662 581984 128358 582040
rect 128414 581984 128419 582040
rect 118601 581982 128419 581984
rect 118601 581979 118667 581982
rect 128353 581979 128419 581982
rect 137921 582042 137987 582045
rect 147673 582042 147739 582045
rect 137921 582040 147739 582042
rect 137921 581984 137926 582040
rect 137982 581984 147678 582040
rect 147734 581984 147739 582040
rect 137921 581982 147739 581984
rect 137921 581979 137987 581982
rect 147673 581979 147739 581982
rect 151670 581980 151676 582044
rect 151740 582042 151746 582044
rect 155861 582042 155927 582045
rect 151740 582040 155927 582042
rect 151740 581984 155866 582040
rect 155922 581984 155927 582040
rect 151740 581982 155927 581984
rect 151740 581980 151746 581982
rect 155861 581979 155927 581982
rect 156321 582042 156387 582045
rect 156454 582042 156460 582044
rect 156321 582040 156460 582042
rect 156321 581984 156326 582040
rect 156382 581984 156460 582040
rect 156321 581982 156460 581984
rect 156321 581979 156387 581982
rect 156454 581980 156460 581982
rect 156524 581980 156530 582044
rect 157149 582042 157215 582045
rect 167085 582042 167151 582045
rect 157149 582040 167151 582042
rect 157149 581984 157154 582040
rect 157210 581984 167090 582040
rect 167146 581984 167151 582040
rect 157149 581982 167151 581984
rect 157149 581979 157215 581982
rect 167085 581979 167151 581982
rect 176561 582042 176627 582045
rect 186313 582042 186379 582045
rect 176561 582040 186379 582042
rect 176561 581984 176566 582040
rect 176622 581984 186318 582040
rect 186374 581984 186379 582040
rect 176561 581982 186379 581984
rect 176561 581979 176627 581982
rect 186313 581979 186379 581982
rect 195881 582042 195947 582045
rect 203333 582042 203399 582045
rect 195881 582040 203399 582042
rect 195881 581984 195886 582040
rect 195942 581984 203338 582040
rect 203394 581984 203399 582040
rect 195881 581982 203399 581984
rect 195881 581979 195947 581982
rect 203333 581979 203399 581982
rect 210325 582042 210391 582045
rect 220905 582042 220971 582045
rect 210325 582040 220971 582042
rect 210325 581984 210330 582040
rect 210386 581984 220910 582040
rect 220966 581984 220971 582040
rect 210325 581982 220971 581984
rect 210325 581979 210391 581982
rect 220905 581979 220971 581982
rect 221222 581980 221228 582044
rect 221292 582042 221298 582044
rect 229318 582042 229324 582044
rect 221292 581982 229324 582042
rect 221292 581980 221298 581982
rect 229318 581980 229324 581982
rect 229388 581980 229394 582044
rect 229461 582042 229527 582045
rect 236453 582042 236519 582045
rect 229461 582040 236519 582042
rect 229461 581984 229466 582040
rect 229522 581984 236458 582040
rect 236514 581984 236519 582040
rect 229461 581982 236519 581984
rect 229461 581979 229527 581982
rect 236453 581979 236519 581982
rect 238753 582042 238819 582045
rect 249742 582042 249748 582044
rect 238753 582040 249748 582042
rect 238753 581984 238758 582040
rect 238814 581984 249748 582040
rect 238753 581982 249748 581984
rect 238753 581979 238819 581982
rect 249742 581980 249748 581982
rect 249812 581980 249818 582044
rect 258165 582042 258231 582045
rect 268510 582042 268516 582044
rect 258165 582040 268516 582042
rect 258165 581984 258170 582040
rect 258226 581984 268516 582040
rect 258165 581982 268516 581984
rect 258165 581979 258231 581982
rect 268510 581980 268516 581982
rect 268580 581980 268586 582044
rect 277710 581980 277716 582044
rect 277780 582042 277786 582044
rect 287646 582042 287652 582044
rect 277780 581982 287652 582042
rect 277780 581980 277786 581982
rect 287646 581980 287652 581982
rect 287716 581980 287722 582044
rect 297398 581980 297404 582044
rect 297468 582042 297474 582044
rect 306046 582042 306052 582044
rect 297468 581982 306052 582042
rect 297468 581980 297474 581982
rect 306046 581980 306052 581982
rect 306116 581980 306122 582044
rect 306281 582042 306347 582045
rect 497406 582042 497412 582044
rect 306281 582040 497412 582042
rect 306281 581984 306286 582040
rect 306342 581984 497412 582040
rect 306281 581982 497412 581984
rect 306281 581979 306347 581982
rect 497406 581980 497412 581982
rect 497476 581980 497482 582044
rect 497549 582042 497615 582045
rect 504909 582042 504975 582045
rect 497549 582040 504975 582042
rect 497549 581984 497554 582040
rect 497610 581984 504914 582040
rect 504970 581984 504975 582040
rect 497549 581982 504975 581984
rect 497549 581979 497615 581982
rect 504909 581979 504975 581982
rect -960 581620 480 581860
rect 84878 581844 84884 581908
rect 84948 581906 84954 581908
rect 89805 581906 89871 581909
rect 84948 581904 89871 581906
rect 84948 581848 89810 581904
rect 89866 581848 89871 581904
rect 84948 581846 89871 581848
rect 84948 581844 84954 581846
rect 89805 581843 89871 581846
rect 91318 581844 91324 581908
rect 91388 581906 91394 581908
rect 91686 581906 91692 581908
rect 91388 581846 91692 581906
rect 91388 581844 91394 581846
rect 91686 581844 91692 581846
rect 91756 581844 91762 581908
rect 91921 581906 91987 581909
rect 208301 581906 208367 581909
rect 91921 581904 208367 581906
rect 91921 581848 91926 581904
rect 91982 581848 208306 581904
rect 208362 581848 208367 581904
rect 91921 581846 208367 581848
rect 91921 581843 91987 581846
rect 208301 581843 208367 581846
rect 210417 581906 210483 581909
rect 220077 581906 220143 581909
rect 210417 581904 220143 581906
rect 210417 581848 210422 581904
rect 210478 581848 220082 581904
rect 220138 581848 220143 581904
rect 210417 581846 220143 581848
rect 210417 581843 210483 581846
rect 220077 581843 220143 581846
rect 220721 581906 220787 581909
rect 230105 581906 230171 581909
rect 220721 581904 230171 581906
rect 220721 581848 220726 581904
rect 220782 581848 230110 581904
rect 230166 581848 230171 581904
rect 220721 581846 230171 581848
rect 220721 581843 220787 581846
rect 230105 581843 230171 581846
rect 239029 581906 239095 581909
rect 249006 581906 249012 581908
rect 239029 581904 249012 581906
rect 239029 581848 239034 581904
rect 239090 581848 249012 581904
rect 239029 581846 249012 581848
rect 239029 581843 239095 581846
rect 249006 581844 249012 581846
rect 249076 581844 249082 581908
rect 249241 581906 249307 581909
rect 256233 581906 256299 581909
rect 249241 581904 256299 581906
rect 249241 581848 249246 581904
rect 249302 581848 256238 581904
rect 256294 581848 256299 581904
rect 249241 581846 256299 581848
rect 249241 581843 249307 581846
rect 256233 581843 256299 581846
rect 258942 581844 258948 581908
rect 259012 581906 259018 581908
rect 268326 581906 268332 581908
rect 259012 581846 268332 581906
rect 259012 581844 259018 581846
rect 268326 581844 268332 581846
rect 268396 581844 268402 581908
rect 282545 581906 282611 581909
rect 498142 581906 498148 581908
rect 282545 581904 498148 581906
rect 282545 581848 282550 581904
rect 282606 581848 498148 581904
rect 282545 581846 498148 581848
rect 282545 581843 282611 581846
rect 498142 581844 498148 581846
rect 498212 581844 498218 581908
rect 85614 581708 85620 581772
rect 85684 581770 85690 581772
rect 86309 581770 86375 581773
rect 85684 581768 86375 581770
rect 85684 581712 86314 581768
rect 86370 581712 86375 581768
rect 85684 581710 86375 581712
rect 85684 581708 85690 581710
rect 86309 581707 86375 581710
rect 88006 581708 88012 581772
rect 88076 581770 88082 581772
rect 94221 581770 94287 581773
rect 88076 581768 94287 581770
rect 88076 581712 94226 581768
rect 94282 581712 94287 581768
rect 88076 581710 94287 581712
rect 88076 581708 88082 581710
rect 94221 581707 94287 581710
rect 96889 581770 96955 581773
rect 331949 581770 332015 581773
rect 96889 581768 332015 581770
rect 96889 581712 96894 581768
rect 96950 581712 331954 581768
rect 332010 581712 332015 581768
rect 96889 581710 332015 581712
rect 96889 581707 96955 581710
rect 331949 581707 332015 581710
rect 335854 581708 335860 581772
rect 335924 581770 335930 581772
rect 350390 581770 350396 581772
rect 335924 581710 350396 581770
rect 335924 581708 335930 581710
rect 350390 581708 350396 581710
rect 350460 581708 350466 581772
rect 355358 581708 355364 581772
rect 355428 581770 355434 581772
rect 364742 581770 364748 581772
rect 355428 581710 364748 581770
rect 355428 581708 355434 581710
rect 364742 581708 364748 581710
rect 364812 581708 364818 581772
rect 374126 581708 374132 581772
rect 374196 581770 374202 581772
rect 384430 581770 384436 581772
rect 374196 581710 384436 581770
rect 374196 581708 374202 581710
rect 384430 581708 384436 581710
rect 384500 581708 384506 581772
rect 393262 581708 393268 581772
rect 393332 581770 393338 581772
rect 403566 581770 403572 581772
rect 393332 581710 403572 581770
rect 393332 581708 393338 581710
rect 403566 581708 403572 581710
rect 403636 581708 403642 581772
rect 418153 581770 418219 581773
rect 498326 581770 498332 581772
rect 418153 581768 498332 581770
rect 418153 581712 418158 581768
rect 418214 581712 498332 581768
rect 418153 581710 498332 581712
rect 418153 581707 418219 581710
rect 498326 581708 498332 581710
rect 498396 581708 498402 581772
rect 86350 581572 86356 581636
rect 86420 581634 86426 581636
rect 89069 581634 89135 581637
rect 86420 581632 89135 581634
rect 86420 581576 89074 581632
rect 89130 581576 89135 581632
rect 86420 581574 89135 581576
rect 86420 581572 86426 581574
rect 89069 581571 89135 581574
rect 89805 581634 89871 581637
rect 108982 581634 108988 581636
rect 89805 581632 108988 581634
rect 89805 581576 89810 581632
rect 89866 581576 108988 581632
rect 89805 581574 108988 581576
rect 89805 581571 89871 581574
rect 108982 581572 108988 581574
rect 109052 581572 109058 581636
rect 111057 581634 111123 581637
rect 118509 581634 118575 581637
rect 111057 581632 118575 581634
rect 111057 581576 111062 581632
rect 111118 581576 118514 581632
rect 118570 581576 118575 581632
rect 111057 581574 118575 581576
rect 111057 581571 111123 581574
rect 118509 581571 118575 581574
rect 128118 581572 128124 581636
rect 128188 581634 128194 581636
rect 128302 581634 128308 581636
rect 128188 581574 128308 581634
rect 128188 581572 128194 581574
rect 128302 581572 128308 581574
rect 128372 581572 128378 581636
rect 137870 581572 137876 581636
rect 137940 581634 137946 581636
rect 147857 581634 147923 581637
rect 137940 581632 147923 581634
rect 137940 581576 147862 581632
rect 147918 581576 147923 581632
rect 137940 581574 147923 581576
rect 137940 581572 137946 581574
rect 147857 581571 147923 581574
rect 153929 581634 153995 581637
rect 156597 581634 156663 581637
rect 153929 581632 156663 581634
rect 153929 581576 153934 581632
rect 153990 581576 156602 581632
rect 156658 581576 156663 581632
rect 153929 581574 156663 581576
rect 153929 581571 153995 581574
rect 156597 581571 156663 581574
rect 157190 581572 157196 581636
rect 157260 581634 157266 581636
rect 166993 581634 167059 581637
rect 186262 581634 186268 581636
rect 157260 581632 167059 581634
rect 157260 581576 166998 581632
rect 167054 581576 167059 581632
rect 157260 581574 167059 581576
rect 157260 581572 157266 581574
rect 166993 581571 167059 581574
rect 181302 581574 186268 581634
rect 84326 581436 84332 581500
rect 84396 581498 84402 581500
rect 85205 581498 85271 581501
rect 85481 581500 85547 581501
rect 85430 581498 85436 581500
rect 84396 581496 85271 581498
rect 84396 581440 85210 581496
rect 85266 581440 85271 581496
rect 84396 581438 85271 581440
rect 85390 581438 85436 581498
rect 85500 581496 85547 581500
rect 85542 581440 85547 581496
rect 84396 581436 84402 581438
rect 85205 581435 85271 581438
rect 85430 581436 85436 581438
rect 85500 581436 85547 581440
rect 85481 581435 85547 581436
rect 93761 581498 93827 581501
rect 99465 581498 99531 581501
rect 93761 581496 99531 581498
rect 93761 581440 93766 581496
rect 93822 581440 99470 581496
rect 99526 581440 99531 581496
rect 93761 581438 99531 581440
rect 93761 581435 93827 581438
rect 99465 581435 99531 581438
rect 99833 581498 99899 581501
rect 113265 581498 113331 581501
rect 99833 581496 113331 581498
rect 99833 581440 99838 581496
rect 99894 581440 113270 581496
rect 113326 581440 113331 581496
rect 99833 581438 113331 581440
rect 99833 581435 99899 581438
rect 113265 581435 113331 581438
rect 113582 581436 113588 581500
rect 113652 581498 113658 581500
rect 123334 581498 123340 581500
rect 113652 581438 123340 581498
rect 113652 581436 113658 581438
rect 123334 581436 123340 581438
rect 123404 581436 123410 581500
rect 123477 581498 123543 581501
rect 132585 581498 132651 581501
rect 123477 581496 132651 581498
rect 123477 581440 123482 581496
rect 123538 581440 132590 581496
rect 132646 581440 132651 581496
rect 123477 581438 132651 581440
rect 123477 581435 123543 581438
rect 132585 581435 132651 581438
rect 132953 581498 133019 581501
rect 142797 581498 142863 581501
rect 157057 581498 157123 581501
rect 132953 581496 137938 581498
rect 132953 581440 132958 581496
rect 133014 581440 137938 581496
rect 132953 581438 137938 581440
rect 132953 581435 133019 581438
rect 84929 581362 84995 581365
rect 89253 581364 89319 581365
rect 87454 581362 87460 581364
rect 84929 581360 87460 581362
rect 84929 581304 84934 581360
rect 84990 581304 87460 581360
rect 84929 581302 87460 581304
rect 84929 581299 84995 581302
rect 87454 581300 87460 581302
rect 87524 581300 87530 581364
rect 89253 581360 89300 581364
rect 89364 581362 89370 581364
rect 89253 581304 89258 581360
rect 89253 581300 89300 581304
rect 89364 581302 89410 581362
rect 89364 581300 89370 581302
rect 90030 581300 90036 581364
rect 90100 581362 90106 581364
rect 90449 581362 90515 581365
rect 90100 581360 90515 581362
rect 90100 581304 90454 581360
rect 90510 581304 90515 581360
rect 90100 581302 90515 581304
rect 90100 581300 90106 581302
rect 89253 581299 89319 581300
rect 90449 581299 90515 581302
rect 90582 581300 90588 581364
rect 90652 581362 90658 581364
rect 90909 581362 90975 581365
rect 91737 581364 91803 581365
rect 91686 581362 91692 581364
rect 90652 581360 90975 581362
rect 90652 581304 90914 581360
rect 90970 581304 90975 581360
rect 90652 581302 90975 581304
rect 91646 581302 91692 581362
rect 91756 581360 91803 581364
rect 91798 581304 91803 581360
rect 90652 581300 90658 581302
rect 90909 581299 90975 581302
rect 91686 581300 91692 581302
rect 91756 581300 91803 581304
rect 92422 581300 92428 581364
rect 92492 581362 92498 581364
rect 92657 581362 92723 581365
rect 93209 581364 93275 581365
rect 93158 581362 93164 581364
rect 92492 581360 92723 581362
rect 92492 581304 92662 581360
rect 92718 581304 92723 581360
rect 92492 581302 92723 581304
rect 93118 581302 93164 581362
rect 93228 581360 93275 581364
rect 93270 581304 93275 581360
rect 92492 581300 92498 581302
rect 91737 581299 91803 581300
rect 92657 581299 92723 581302
rect 93158 581300 93164 581302
rect 93228 581300 93275 581304
rect 93209 581299 93275 581300
rect 93393 581362 93459 581365
rect 96889 581362 96955 581365
rect 100017 581362 100083 581365
rect 93393 581360 96955 581362
rect 93393 581304 93398 581360
rect 93454 581304 96894 581360
rect 96950 581304 96955 581360
rect 93393 581302 96955 581304
rect 93393 581299 93459 581302
rect 96889 581299 96955 581302
rect 99974 581360 100083 581362
rect 99974 581304 100022 581360
rect 100078 581304 100083 581360
rect 99974 581299 100083 581304
rect 103421 581362 103487 581365
rect 108941 581362 109007 581365
rect 103421 581360 109007 581362
rect 103421 581304 103426 581360
rect 103482 581304 108946 581360
rect 109002 581304 109007 581360
rect 103421 581302 109007 581304
rect 103421 581299 103487 581302
rect 108941 581299 109007 581302
rect 109125 581360 109191 581365
rect 109125 581304 109130 581360
rect 109186 581304 109191 581360
rect 109125 581299 109191 581304
rect 109350 581300 109356 581364
rect 109420 581362 109426 581364
rect 115197 581362 115263 581365
rect 109420 581360 115263 581362
rect 109420 581304 115202 581360
rect 115258 581304 115263 581360
rect 109420 581302 115263 581304
rect 109420 581300 109426 581302
rect 115197 581299 115263 581302
rect 115841 581362 115907 581365
rect 118693 581362 118759 581365
rect 137878 581362 137938 581438
rect 142797 581496 157123 581498
rect 142797 581440 142802 581496
rect 142858 581440 157062 581496
rect 157118 581440 157123 581496
rect 142797 581438 157123 581440
rect 142797 581435 142863 581438
rect 157057 581435 157123 581438
rect 157517 581498 157583 581501
rect 171777 581498 171843 581501
rect 157517 581496 171843 581498
rect 157517 581440 157522 581496
rect 157578 581440 171782 581496
rect 171838 581440 171843 581496
rect 157517 581438 171843 581440
rect 157517 581435 157583 581438
rect 171777 581435 171843 581438
rect 171961 581498 172027 581501
rect 181302 581498 181362 581574
rect 186262 581572 186268 581574
rect 186332 581572 186338 581636
rect 195830 581572 195836 581636
rect 195900 581634 195906 581636
rect 197997 581634 198063 581637
rect 205582 581634 205588 581636
rect 195900 581632 198063 581634
rect 195900 581576 198002 581632
rect 198058 581576 198063 581632
rect 195900 581574 198063 581576
rect 195900 581572 195906 581574
rect 197997 581571 198063 581574
rect 200622 581574 205588 581634
rect 171961 581496 181362 581498
rect 171961 581440 171966 581496
rect 172022 581440 181362 581496
rect 171961 581438 181362 581440
rect 181437 581498 181503 581501
rect 190821 581498 190887 581501
rect 181437 581496 190887 581498
rect 181437 581440 181442 581496
rect 181498 581440 190826 581496
rect 190882 581440 190887 581496
rect 181437 581438 190887 581440
rect 171961 581435 172027 581438
rect 181437 581435 181503 581438
rect 190821 581435 190887 581438
rect 191046 581436 191052 581500
rect 191116 581498 191122 581500
rect 200622 581498 200682 581574
rect 205582 581572 205588 581574
rect 205652 581572 205658 581636
rect 224902 581634 224908 581636
rect 219942 581574 224908 581634
rect 191116 581438 200682 581498
rect 200757 581498 200823 581501
rect 210417 581498 210483 581501
rect 219942 581498 220002 581574
rect 224902 581572 224908 581574
rect 224972 581572 224978 581636
rect 244222 581634 244228 581636
rect 236318 581574 244228 581634
rect 200757 581496 210483 581498
rect 200757 581440 200762 581496
rect 200818 581440 210422 581496
rect 210478 581440 210483 581496
rect 200757 581438 210483 581440
rect 191116 581436 191122 581438
rect 200757 581435 200823 581438
rect 210417 581435 210483 581438
rect 210742 581438 220002 581498
rect 220077 581498 220143 581501
rect 229461 581498 229527 581501
rect 236318 581498 236378 581574
rect 244222 581572 244228 581574
rect 244292 581572 244298 581636
rect 256325 581634 256391 581637
rect 260598 581634 260604 581636
rect 256325 581632 260604 581634
rect 256325 581576 256330 581632
rect 256386 581576 260604 581632
rect 256325 581574 260604 581576
rect 256325 581571 256391 581574
rect 260598 581572 260604 581574
rect 260668 581572 260674 581636
rect 273161 581634 273227 581637
rect 282913 581634 282979 581637
rect 273161 581632 282979 581634
rect 273161 581576 273166 581632
rect 273222 581576 282918 581632
rect 282974 581576 282979 581632
rect 273161 581574 282979 581576
rect 273161 581571 273227 581574
rect 282913 581571 282979 581574
rect 292481 581634 292547 581637
rect 302233 581634 302299 581637
rect 292481 581632 302299 581634
rect 292481 581576 292486 581632
rect 292542 581576 302238 581632
rect 302294 581576 302299 581632
rect 292481 581574 302299 581576
rect 292481 581571 292547 581574
rect 302233 581571 302299 581574
rect 311801 581634 311867 581637
rect 321553 581634 321619 581637
rect 311801 581632 321619 581634
rect 311801 581576 311806 581632
rect 311862 581576 321558 581632
rect 321614 581576 321619 581632
rect 311801 581574 321619 581576
rect 311801 581571 311867 581574
rect 321553 581571 321619 581574
rect 321870 581572 321876 581636
rect 321940 581634 321946 581636
rect 324773 581634 324839 581637
rect 346853 581636 346919 581637
rect 351637 581636 351703 581637
rect 321940 581632 324839 581634
rect 321940 581576 324778 581632
rect 324834 581576 324839 581632
rect 321940 581574 324839 581576
rect 321940 581572 321946 581574
rect 324773 581571 324839 581574
rect 336038 581572 336044 581636
rect 336108 581634 336114 581636
rect 345606 581634 345612 581636
rect 336108 581574 345612 581634
rect 336108 581572 336114 581574
rect 345606 581572 345612 581574
rect 345676 581572 345682 581636
rect 346853 581632 346900 581636
rect 346964 581634 346970 581636
rect 346853 581576 346858 581632
rect 346853 581572 346900 581576
rect 346964 581574 347010 581634
rect 351637 581632 351684 581636
rect 351748 581634 351754 581636
rect 351637 581576 351642 581632
rect 346964 581572 346970 581574
rect 351637 581572 351684 581576
rect 351748 581574 351794 581634
rect 351748 581572 351754 581574
rect 355174 581572 355180 581636
rect 355244 581634 355250 581636
rect 360142 581634 360148 581636
rect 355244 581574 360148 581634
rect 355244 581572 355250 581574
rect 360142 581572 360148 581574
rect 360212 581572 360218 581636
rect 365110 581572 365116 581636
rect 365180 581634 365186 581636
rect 365253 581634 365319 581637
rect 384849 581636 384915 581637
rect 365180 581632 365319 581634
rect 365180 581576 365258 581632
rect 365314 581576 365319 581632
rect 365180 581574 365319 581576
rect 365180 581572 365186 581574
rect 346853 581571 346919 581572
rect 351637 581571 351703 581572
rect 365253 581571 365319 581574
rect 373942 581572 373948 581636
rect 374012 581634 374018 581636
rect 384246 581634 384252 581636
rect 374012 581574 384252 581634
rect 374012 581572 374018 581574
rect 384246 581572 384252 581574
rect 384316 581572 384322 581636
rect 384798 581634 384804 581636
rect 384758 581574 384804 581634
rect 384868 581632 384915 581636
rect 384910 581576 384915 581632
rect 384798 581572 384804 581574
rect 384868 581572 384915 581576
rect 384849 581571 384915 581572
rect 389725 581636 389791 581637
rect 391749 581636 391815 581637
rect 389725 581632 389772 581636
rect 389836 581634 389842 581636
rect 389725 581576 389730 581632
rect 389725 581572 389772 581576
rect 389836 581574 389882 581634
rect 391749 581632 391796 581636
rect 391860 581634 391866 581636
rect 396993 581634 397059 581637
rect 498694 581634 498700 581636
rect 391749 581576 391754 581632
rect 389836 581572 389842 581574
rect 391749 581572 391796 581576
rect 391860 581574 391906 581634
rect 396993 581632 498700 581634
rect 396993 581576 396998 581632
rect 397054 581576 498700 581632
rect 396993 581574 498700 581576
rect 391860 581572 391866 581574
rect 389725 581571 389791 581572
rect 391749 581571 391815 581572
rect 396993 581571 397059 581574
rect 498694 581572 498700 581574
rect 498764 581572 498770 581636
rect 499982 581572 499988 581636
rect 500052 581634 500058 581636
rect 505001 581634 505067 581637
rect 500052 581632 505067 581634
rect 500052 581576 505006 581632
rect 505062 581576 505067 581632
rect 500052 581574 505067 581576
rect 500052 581572 500058 581574
rect 505001 581571 505067 581574
rect 505185 581634 505251 581637
rect 509969 581634 510035 581637
rect 505185 581632 510035 581634
rect 505185 581576 505190 581632
rect 505246 581576 509974 581632
rect 510030 581576 510035 581632
rect 505185 581574 510035 581576
rect 505185 581571 505251 581574
rect 509969 581571 510035 581574
rect 220077 581496 229527 581498
rect 220077 581440 220082 581496
rect 220138 581440 229466 581496
rect 229522 581440 229527 581496
rect 220077 581438 229527 581440
rect 146937 581362 147003 581365
rect 115841 581360 118759 581362
rect 115841 581304 115846 581360
rect 115902 581304 118698 581360
rect 118754 581304 118759 581360
rect 115841 581302 118759 581304
rect 115841 581299 115907 581302
rect 118693 581299 118759 581302
rect 118926 581302 137754 581362
rect 137878 581360 147003 581362
rect 137878 581304 146942 581360
rect 146998 581304 147003 581360
rect 137878 581302 147003 581304
rect 83774 581164 83780 581228
rect 83844 581226 83850 581228
rect 94262 581226 94268 581228
rect 83844 581166 94268 581226
rect 83844 581164 83850 581166
rect 94262 581164 94268 581166
rect 94332 581164 94338 581228
rect 99974 581226 100034 581299
rect 94454 581166 100034 581226
rect 85798 581028 85804 581092
rect 85868 581090 85874 581092
rect 94454 581090 94514 581166
rect 104382 581164 104388 581228
rect 104452 581226 104458 581228
rect 108798 581226 108804 581228
rect 104452 581166 108804 581226
rect 104452 581164 104458 581166
rect 108798 581164 108804 581166
rect 108868 581164 108874 581228
rect 109128 581226 109188 581299
rect 118550 581226 118556 581228
rect 109128 581166 118556 581226
rect 118550 581164 118556 581166
rect 118620 581164 118626 581228
rect 118926 581226 118986 581302
rect 137318 581226 137324 581228
rect 118742 581166 118986 581226
rect 119110 581166 137324 581226
rect 85868 581030 94514 581090
rect 85868 581028 85874 581030
rect 109350 581028 109356 581092
rect 109420 581090 109426 581092
rect 113582 581090 113588 581092
rect 109420 581030 113588 581090
rect 109420 581028 109426 581030
rect 113582 581028 113588 581030
rect 113652 581028 113658 581092
rect 113766 581028 113772 581092
rect 113836 581090 113842 581092
rect 118742 581090 118802 581166
rect 119110 581090 119170 581166
rect 137318 581164 137324 581166
rect 137388 581164 137394 581228
rect 137694 581226 137754 581302
rect 146937 581299 147003 581302
rect 147857 581362 147923 581365
rect 147857 581360 151922 581362
rect 147857 581304 147862 581360
rect 147918 581304 151922 581360
rect 147857 581302 151922 581304
rect 147857 581299 147923 581302
rect 151670 581226 151676 581228
rect 137694 581166 137938 581226
rect 113836 581030 118802 581090
rect 118926 581030 119170 581090
rect 113836 581028 113842 581030
rect 82302 580892 82308 580956
rect 82372 580954 82378 580956
rect 86350 580954 86356 580956
rect 82372 580894 86356 580954
rect 82372 580892 82378 580894
rect 86350 580892 86356 580894
rect 86420 580892 86426 580956
rect 94262 580892 94268 580956
rect 94332 580954 94338 580956
rect 104382 580954 104388 580956
rect 94332 580894 104388 580954
rect 94332 580892 94338 580894
rect 104382 580892 104388 580894
rect 104452 580892 104458 580956
rect 118550 580756 118556 580820
rect 118620 580818 118626 580820
rect 118926 580818 118986 581030
rect 123334 581028 123340 581092
rect 123404 581090 123410 581092
rect 128118 581090 128124 581092
rect 123404 581030 128124 581090
rect 123404 581028 123410 581030
rect 128118 581028 128124 581030
rect 128188 581028 128194 581092
rect 128302 581028 128308 581092
rect 128372 581090 128378 581092
rect 137502 581090 137508 581092
rect 128372 581030 137508 581090
rect 128372 581028 128378 581030
rect 137502 581028 137508 581030
rect 137572 581028 137578 581092
rect 137878 581090 137938 581166
rect 138246 581166 151676 581226
rect 138054 581090 138060 581092
rect 137878 581030 138060 581090
rect 138054 581028 138060 581030
rect 138124 581028 138130 581092
rect 137318 580892 137324 580956
rect 137388 580954 137394 580956
rect 138246 580954 138306 581166
rect 151670 581164 151676 581166
rect 151740 581164 151746 581228
rect 151862 581226 151922 581302
rect 156086 581300 156092 581364
rect 156156 581362 156162 581364
rect 157241 581362 157307 581365
rect 156156 581360 157307 581362
rect 156156 581304 157246 581360
rect 157302 581304 157307 581360
rect 156156 581302 157307 581304
rect 156156 581300 156162 581302
rect 157241 581299 157307 581302
rect 166901 581362 166967 581365
rect 176561 581362 176627 581365
rect 166901 581360 176627 581362
rect 166901 581304 166906 581360
rect 166962 581304 176566 581360
rect 176622 581304 176627 581360
rect 166901 581302 176627 581304
rect 166901 581299 166967 581302
rect 176561 581299 176627 581302
rect 176745 581362 176811 581365
rect 192017 581362 192083 581365
rect 176745 581360 192083 581362
rect 176745 581304 176750 581360
rect 176806 581304 192022 581360
rect 192078 581304 192083 581360
rect 176745 581302 192083 581304
rect 176745 581299 176811 581302
rect 192017 581299 192083 581302
rect 192201 581362 192267 581365
rect 195881 581362 195947 581365
rect 192201 581360 195947 581362
rect 192201 581304 192206 581360
rect 192262 581304 195886 581360
rect 195942 581304 195947 581360
rect 192201 581302 195947 581304
rect 192201 581299 192267 581302
rect 195881 581299 195947 581302
rect 200665 581362 200731 581365
rect 210325 581362 210391 581365
rect 200665 581360 210391 581362
rect 200665 581304 200670 581360
rect 200726 581304 210330 581360
rect 210386 581304 210391 581360
rect 200665 581302 210391 581304
rect 200665 581299 200731 581302
rect 210325 581299 210391 581302
rect 151862 581166 156338 581226
rect 138422 581028 138428 581092
rect 138492 581090 138498 581092
rect 156086 581090 156092 581092
rect 138492 581030 156092 581090
rect 138492 581028 138498 581030
rect 156086 581028 156092 581030
rect 156156 581028 156162 581092
rect 156278 581090 156338 581166
rect 156454 581164 156460 581228
rect 156524 581226 156530 581228
rect 161422 581226 161428 581228
rect 156524 581166 161428 581226
rect 156524 581164 156530 581166
rect 161422 581164 161428 581166
rect 161492 581164 161498 581228
rect 162342 581164 162348 581228
rect 162412 581226 162418 581228
rect 181662 581226 181668 581228
rect 162412 581166 181668 581226
rect 162412 581164 162418 581166
rect 181662 581164 181668 581166
rect 181732 581164 181738 581228
rect 186262 581164 186268 581228
rect 186332 581226 186338 581228
rect 190494 581226 190500 581228
rect 186332 581166 190500 581226
rect 186332 581164 186338 581166
rect 190494 581164 190500 581166
rect 190564 581164 190570 581228
rect 190678 581164 190684 581228
rect 190748 581226 190754 581228
rect 200982 581226 200988 581228
rect 190748 581166 200988 581226
rect 190748 581164 190754 581166
rect 200982 581164 200988 581166
rect 201052 581164 201058 581228
rect 205582 581164 205588 581228
rect 205652 581226 205658 581228
rect 210742 581226 210802 581438
rect 220077 581435 220143 581438
rect 229461 581435 229527 581438
rect 229694 581438 236378 581498
rect 236453 581498 236519 581501
rect 253381 581498 253447 581501
rect 236453 581496 253447 581498
rect 236453 581440 236458 581496
rect 236514 581440 253386 581496
rect 253442 581440 253447 581496
rect 236453 581438 253447 581440
rect 211153 581362 211219 581365
rect 220721 581362 220787 581365
rect 211153 581360 211354 581362
rect 211153 581304 211158 581360
rect 211214 581304 211354 581360
rect 211153 581302 211354 581304
rect 211153 581299 211219 581302
rect 205652 581166 210802 581226
rect 211294 581226 211354 581302
rect 220126 581360 220787 581362
rect 220126 581304 220726 581360
rect 220782 581304 220787 581360
rect 220126 581302 220787 581304
rect 220126 581226 220186 581302
rect 220721 581299 220787 581302
rect 220905 581362 220971 581365
rect 229369 581362 229435 581365
rect 220905 581360 229435 581362
rect 220905 581304 220910 581360
rect 220966 581304 229374 581360
rect 229430 581304 229435 581360
rect 220905 581302 229435 581304
rect 220905 581299 220971 581302
rect 229369 581299 229435 581302
rect 211294 581166 220186 581226
rect 205652 581164 205658 581166
rect 224902 581164 224908 581228
rect 224972 581226 224978 581228
rect 229694 581226 229754 581438
rect 236453 581435 236519 581438
rect 253381 581435 253447 581438
rect 256233 581498 256299 581501
rect 263501 581498 263567 581501
rect 256233 581496 263567 581498
rect 256233 581440 256238 581496
rect 256294 581440 263506 581496
rect 263562 581440 263567 581496
rect 256233 581438 263567 581440
rect 256233 581435 256299 581438
rect 263501 581435 263567 581438
rect 263685 581498 263751 581501
rect 506422 581498 506428 581500
rect 263685 581496 506428 581498
rect 263685 581440 263690 581496
rect 263746 581440 506428 581496
rect 263685 581438 506428 581440
rect 263685 581435 263751 581438
rect 506422 581436 506428 581438
rect 506492 581436 506498 581500
rect 536054 581438 543842 581498
rect 230105 581362 230171 581365
rect 231945 581364 232011 581365
rect 231894 581362 231900 581364
rect 230105 581360 230306 581362
rect 230105 581304 230110 581360
rect 230166 581304 230306 581360
rect 230105 581302 230306 581304
rect 231854 581302 231900 581362
rect 231964 581360 232011 581364
rect 238753 581362 238819 581365
rect 239029 581362 239095 581365
rect 232006 581304 232011 581360
rect 230105 581299 230171 581302
rect 224972 581166 229754 581226
rect 230246 581226 230306 581302
rect 231894 581300 231900 581302
rect 231964 581300 232011 581304
rect 231945 581299 232011 581300
rect 238710 581360 238819 581362
rect 238710 581304 238758 581360
rect 238814 581304 238819 581360
rect 238710 581299 238819 581304
rect 238894 581360 239095 581362
rect 238894 581304 239034 581360
rect 239090 581304 239095 581360
rect 238894 581302 239095 581304
rect 238710 581226 238770 581299
rect 230246 581166 238770 581226
rect 224972 581164 224978 581166
rect 157190 581090 157196 581092
rect 156278 581030 157196 581090
rect 157190 581028 157196 581030
rect 157260 581028 157266 581092
rect 210366 581028 210372 581092
rect 210436 581090 210442 581092
rect 221222 581090 221228 581092
rect 210436 581030 221228 581090
rect 210436 581028 210442 581030
rect 221222 581028 221228 581030
rect 221292 581028 221298 581092
rect 229318 581028 229324 581092
rect 229388 581090 229394 581092
rect 238894 581090 238954 581302
rect 239029 581299 239095 581302
rect 239673 581362 239739 581365
rect 249241 581362 249307 581365
rect 256325 581362 256391 581365
rect 258165 581362 258231 581365
rect 239673 581360 249307 581362
rect 239673 581304 239678 581360
rect 239734 581304 249246 581360
rect 249302 581304 249307 581360
rect 239673 581302 249307 581304
rect 239673 581299 239739 581302
rect 249241 581299 249307 581302
rect 249566 581360 256391 581362
rect 249566 581304 256330 581360
rect 256386 581304 256391 581360
rect 249566 581302 256391 581304
rect 244222 581164 244228 581228
rect 244292 581226 244298 581228
rect 249566 581226 249626 581302
rect 256325 581299 256391 581302
rect 258030 581360 258231 581362
rect 258030 581304 258170 581360
rect 258226 581304 258231 581360
rect 258030 581302 258231 581304
rect 244292 581166 249626 581226
rect 244292 581164 244298 581166
rect 249742 581164 249748 581228
rect 249812 581226 249818 581228
rect 258030 581226 258090 581302
rect 258165 581299 258231 581302
rect 258349 581362 258415 581365
rect 263501 581362 263567 581365
rect 258349 581360 263567 581362
rect 258349 581304 258354 581360
rect 258410 581304 263506 581360
rect 263562 581304 263567 581360
rect 258349 581302 263567 581304
rect 258349 581299 258415 581302
rect 263501 581299 263567 581302
rect 263685 581362 263751 581365
rect 358721 581364 358787 581365
rect 358670 581362 358676 581364
rect 263685 581360 355426 581362
rect 263685 581304 263690 581360
rect 263746 581304 355426 581360
rect 263685 581302 355426 581304
rect 358630 581302 358676 581362
rect 358740 581360 358787 581364
rect 523033 581362 523099 581365
rect 536054 581362 536114 581438
rect 358782 581304 358787 581360
rect 263685 581299 263751 581302
rect 249812 581166 258090 581226
rect 249812 581164 249818 581166
rect 260598 581164 260604 581228
rect 260668 581226 260674 581228
rect 260782 581226 260788 581228
rect 260668 581166 260788 581226
rect 260668 581164 260674 581166
rect 260782 581164 260788 581166
rect 260852 581164 260858 581228
rect 268510 581164 268516 581228
rect 268580 581226 268586 581228
rect 277526 581226 277532 581228
rect 268580 581166 277532 581226
rect 268580 581164 268586 581166
rect 277526 581164 277532 581166
rect 277596 581164 277602 581228
rect 287830 581164 287836 581228
rect 287900 581226 287906 581228
rect 297214 581226 297220 581228
rect 287900 581166 297220 581226
rect 287900 581164 287906 581166
rect 297214 581164 297220 581166
rect 297284 581164 297290 581228
rect 306598 581164 306604 581228
rect 306668 581226 306674 581228
rect 316718 581226 316724 581228
rect 306668 581166 316724 581226
rect 306668 581164 306674 581166
rect 316718 581164 316724 581166
rect 316788 581164 316794 581228
rect 326286 581164 326292 581228
rect 326356 581226 326362 581228
rect 335854 581226 335860 581228
rect 326356 581166 335860 581226
rect 326356 581164 326362 581166
rect 335854 581164 335860 581166
rect 335924 581164 335930 581228
rect 350390 581164 350396 581228
rect 350460 581226 350466 581228
rect 355174 581226 355180 581228
rect 350460 581166 355180 581226
rect 350460 581164 350466 581166
rect 355174 581164 355180 581166
rect 355244 581164 355250 581228
rect 355366 581226 355426 581302
rect 358670 581300 358676 581302
rect 358740 581300 358787 581304
rect 358721 581299 358787 581300
rect 358862 581360 523099 581362
rect 358862 581304 523038 581360
rect 523094 581304 523099 581360
rect 358862 581302 523099 581304
rect 358862 581226 358922 581302
rect 523033 581299 523099 581302
rect 524462 581302 536114 581362
rect 543782 581362 543842 581438
rect 550582 581362 550588 581364
rect 543782 581302 550588 581362
rect 355366 581166 358922 581226
rect 360142 581164 360148 581228
rect 360212 581226 360218 581228
rect 374126 581226 374132 581228
rect 360212 581166 374132 581226
rect 360212 581164 360218 581166
rect 374126 581164 374132 581166
rect 374196 581164 374202 581228
rect 384430 581164 384436 581228
rect 384500 581226 384506 581228
rect 393446 581226 393452 581228
rect 384500 581166 393452 581226
rect 384500 581164 384506 581166
rect 393446 581164 393452 581166
rect 393516 581164 393522 581228
rect 403750 581164 403756 581228
rect 403820 581226 403826 581228
rect 412766 581226 412772 581228
rect 403820 581166 412772 581226
rect 403820 581164 403826 581166
rect 412766 581164 412772 581166
rect 412836 581164 412842 581228
rect 423070 581164 423076 581228
rect 423140 581226 423146 581228
rect 432086 581226 432092 581228
rect 423140 581166 432092 581226
rect 423140 581164 423146 581166
rect 432086 581164 432092 581166
rect 432156 581164 432162 581228
rect 437422 581164 437428 581228
rect 437492 581226 437498 581228
rect 456558 581226 456564 581228
rect 437492 581166 456564 581226
rect 437492 581164 437498 581166
rect 456558 581164 456564 581166
rect 456628 581164 456634 581228
rect 456742 581164 456748 581228
rect 456812 581226 456818 581228
rect 470726 581226 470732 581228
rect 456812 581166 470732 581226
rect 456812 581164 456818 581166
rect 470726 581164 470732 581166
rect 470796 581164 470802 581228
rect 476062 581164 476068 581228
rect 476132 581226 476138 581228
rect 489862 581226 489868 581228
rect 476132 581166 489868 581226
rect 476132 581164 476138 581166
rect 489862 581164 489868 581166
rect 489932 581164 489938 581228
rect 495382 581164 495388 581228
rect 495452 581226 495458 581228
rect 499982 581226 499988 581228
rect 495452 581166 499988 581226
rect 495452 581164 495458 581166
rect 499982 581164 499988 581166
rect 500052 581164 500058 581228
rect 504909 581226 504975 581229
rect 509182 581226 509188 581228
rect 504909 581224 509188 581226
rect 504909 581168 504914 581224
rect 504970 581168 509188 581224
rect 504909 581166 509188 581168
rect 504909 581163 504975 581166
rect 509182 581164 509188 581166
rect 509252 581164 509258 581228
rect 509969 581226 510035 581229
rect 524462 581226 524522 581302
rect 550582 581300 550588 581302
rect 550652 581300 550658 581364
rect 509969 581224 524522 581226
rect 509969 581168 509974 581224
rect 510030 581168 524522 581224
rect 509969 581166 524522 581168
rect 509969 581163 510035 581166
rect 229388 581030 238954 581090
rect 229388 581028 229394 581030
rect 249006 581028 249012 581092
rect 249076 581090 249082 581092
rect 258942 581090 258948 581092
rect 249076 581030 258948 581090
rect 249076 581028 249082 581030
rect 258942 581028 258948 581030
rect 259012 581028 259018 581092
rect 268326 581028 268332 581092
rect 268396 581090 268402 581092
rect 277710 581090 277716 581092
rect 268396 581030 277716 581090
rect 268396 581028 268402 581030
rect 277710 581028 277716 581030
rect 277780 581028 277786 581092
rect 287646 581028 287652 581092
rect 287716 581090 287722 581092
rect 297398 581090 297404 581092
rect 287716 581030 297404 581090
rect 287716 581028 287722 581030
rect 297398 581028 297404 581030
rect 297468 581028 297474 581092
rect 306046 581028 306052 581092
rect 306116 581090 306122 581092
rect 316534 581090 316540 581092
rect 306116 581030 316540 581090
rect 306116 581028 306122 581030
rect 316534 581028 316540 581030
rect 316604 581028 316610 581092
rect 326470 581028 326476 581092
rect 326540 581090 326546 581092
rect 336038 581090 336044 581092
rect 326540 581030 336044 581090
rect 326540 581028 326546 581030
rect 336038 581028 336044 581030
rect 336108 581028 336114 581092
rect 345606 581028 345612 581092
rect 345676 581090 345682 581092
rect 355358 581090 355364 581092
rect 345676 581030 355364 581090
rect 345676 581028 345682 581030
rect 355358 581028 355364 581030
rect 355428 581028 355434 581092
rect 364742 581028 364748 581092
rect 364812 581090 364818 581092
rect 373942 581090 373948 581092
rect 364812 581030 373948 581090
rect 364812 581028 364818 581030
rect 373942 581028 373948 581030
rect 374012 581028 374018 581092
rect 384246 581028 384252 581092
rect 384316 581090 384322 581092
rect 393262 581090 393268 581092
rect 384316 581030 393268 581090
rect 384316 581028 384322 581030
rect 393262 581028 393268 581030
rect 393332 581028 393338 581092
rect 403566 581028 403572 581092
rect 403636 581090 403642 581092
rect 412582 581090 412588 581092
rect 403636 581030 412588 581090
rect 403636 581028 403642 581030
rect 412582 581028 412588 581030
rect 412652 581028 412658 581092
rect 422886 581028 422892 581092
rect 422956 581090 422962 581092
rect 431902 581090 431908 581092
rect 422956 581030 431908 581090
rect 422956 581028 422962 581030
rect 431902 581028 431908 581030
rect 431972 581028 431978 581092
rect 442206 581028 442212 581092
rect 442276 581090 442282 581092
rect 451958 581090 451964 581092
rect 442276 581030 451964 581090
rect 442276 581028 442282 581030
rect 451958 581028 451964 581030
rect 452028 581028 452034 581092
rect 461342 581028 461348 581092
rect 461412 581090 461418 581092
rect 470542 581090 470548 581092
rect 461412 581030 470548 581090
rect 461412 581028 461418 581030
rect 470542 581028 470548 581030
rect 470612 581028 470618 581092
rect 480846 581028 480852 581092
rect 480916 581090 480922 581092
rect 489862 581090 489868 581092
rect 480916 581030 489868 581090
rect 480916 581028 480922 581030
rect 489862 581028 489868 581030
rect 489932 581028 489938 581092
rect 505001 581090 505067 581093
rect 505185 581090 505251 581093
rect 505001 581088 505251 581090
rect 505001 581032 505006 581088
rect 505062 581032 505190 581088
rect 505246 581032 505251 581088
rect 505001 581030 505251 581032
rect 505001 581027 505067 581030
rect 505185 581027 505251 581030
rect 550582 581028 550588 581092
rect 550652 581090 550658 581092
rect 558913 581090 558979 581093
rect 550652 581088 558979 581090
rect 550652 581032 558918 581088
rect 558974 581032 558979 581088
rect 550652 581030 558979 581032
rect 550652 581028 550658 581030
rect 558913 581027 558979 581030
rect 137388 580894 138306 580954
rect 137388 580892 137394 580894
rect 179270 580892 179276 580956
rect 179340 580954 179346 580956
rect 195830 580954 195836 580956
rect 179340 580894 195836 580954
rect 179340 580892 179346 580894
rect 195830 580892 195836 580894
rect 195900 580892 195906 580956
rect 389766 580892 389772 580956
rect 389836 580954 389842 580956
rect 506657 580954 506723 580957
rect 389836 580952 506723 580954
rect 389836 580896 506662 580952
rect 506718 580896 506723 580952
rect 389836 580894 506723 580896
rect 389836 580892 389842 580894
rect 506657 580891 506723 580894
rect 118620 580758 118986 580818
rect 118620 580756 118626 580758
rect 384798 580756 384804 580820
rect 384868 580818 384874 580820
rect 501086 580818 501092 580820
rect 384868 580758 501092 580818
rect 384868 580756 384874 580758
rect 501086 580756 501092 580758
rect 501156 580756 501162 580820
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 82494 579866 82554 580652
rect 161422 580620 161428 580684
rect 161492 580682 161498 580684
rect 169702 580682 169708 580684
rect 161492 580622 169708 580682
rect 161492 580620 161498 580622
rect 169702 580620 169708 580622
rect 169772 580620 169778 580684
rect 391790 580620 391796 580684
rect 391860 580682 391866 580684
rect 508497 580682 508563 580685
rect 391860 580680 508563 580682
rect 391860 580624 508502 580680
rect 508558 580624 508563 580680
rect 583520 580668 584960 580758
rect 391860 580622 508563 580624
rect 391860 580620 391866 580622
rect 508497 580619 508563 580622
rect 99966 580484 99972 580548
rect 100036 580546 100042 580548
rect 113766 580546 113772 580548
rect 100036 580486 113772 580546
rect 100036 580484 100042 580486
rect 113766 580484 113772 580486
rect 113836 580484 113842 580548
rect 114502 580484 114508 580548
rect 114572 580546 114578 580548
rect 123702 580546 123708 580548
rect 114572 580486 123708 580546
rect 114572 580484 114578 580486
rect 123702 580484 123708 580486
rect 123772 580484 123778 580548
rect 124254 580484 124260 580548
rect 124324 580546 124330 580548
rect 137134 580546 137140 580548
rect 124324 580486 137140 580546
rect 124324 580484 124330 580486
rect 137134 580484 137140 580486
rect 137204 580484 137210 580548
rect 142102 580484 142108 580548
rect 142172 580546 142178 580548
rect 151486 580546 151492 580548
rect 142172 580486 151492 580546
rect 142172 580484 142178 580486
rect 151486 580484 151492 580486
rect 151556 580484 151562 580548
rect 151854 580484 151860 580548
rect 151924 580546 151930 580548
rect 161238 580546 161244 580548
rect 151924 580486 161244 580546
rect 151924 580484 151930 580486
rect 161238 580484 161244 580486
rect 161308 580484 161314 580548
rect 166206 580484 166212 580548
rect 166276 580546 166282 580548
rect 167678 580546 167684 580548
rect 166276 580486 167684 580546
rect 166276 580484 166282 580486
rect 167678 580484 167684 580486
rect 167748 580484 167754 580548
rect 197302 580484 197308 580548
rect 197372 580546 197378 580548
rect 206870 580546 206876 580548
rect 197372 580486 206876 580546
rect 197372 580484 197378 580486
rect 206870 580484 206876 580486
rect 206940 580484 206946 580548
rect 216622 580484 216628 580548
rect 216692 580546 216698 580548
rect 226190 580546 226196 580548
rect 216692 580486 226196 580546
rect 216692 580484 216698 580486
rect 226190 580484 226196 580486
rect 226260 580484 226266 580548
rect 358670 580484 358676 580548
rect 358740 580546 358746 580548
rect 502006 580546 502012 580548
rect 358740 580486 502012 580546
rect 358740 580484 358746 580486
rect 502006 580484 502012 580486
rect 502076 580484 502082 580548
rect 86902 580348 86908 580412
rect 86972 580410 86978 580412
rect 231894 580410 231900 580412
rect 86972 580350 231900 580410
rect 86972 580348 86978 580350
rect 231894 580348 231900 580350
rect 231964 580348 231970 580412
rect 245694 580348 245700 580412
rect 245764 580410 245770 580412
rect 254894 580410 254900 580412
rect 245764 580350 254900 580410
rect 245764 580348 245770 580350
rect 254894 580348 254900 580350
rect 254964 580348 254970 580412
rect 260966 580348 260972 580412
rect 261036 580410 261042 580412
rect 270350 580410 270356 580412
rect 261036 580350 270356 580410
rect 261036 580348 261042 580350
rect 270350 580348 270356 580350
rect 270420 580348 270426 580412
rect 272558 580348 272564 580412
rect 272628 580410 272634 580412
rect 273846 580410 273852 580412
rect 272628 580350 273852 580410
rect 272628 580348 272634 580350
rect 273846 580348 273852 580350
rect 273916 580348 273922 580412
rect 282310 580348 282316 580412
rect 282380 580410 282386 580412
rect 283414 580410 283420 580412
rect 282380 580350 283420 580410
rect 282380 580348 282386 580350
rect 283414 580348 283420 580350
rect 283484 580348 283490 580412
rect 291878 580348 291884 580412
rect 291948 580410 291954 580412
rect 293166 580410 293172 580412
rect 291948 580350 293172 580410
rect 291948 580348 291954 580350
rect 293166 580348 293172 580350
rect 293236 580348 293242 580412
rect 330702 580348 330708 580412
rect 330772 580410 330778 580412
rect 331806 580410 331812 580412
rect 330772 580350 331812 580410
rect 330772 580348 330778 580350
rect 331806 580348 331812 580350
rect 331876 580348 331882 580412
rect 338062 580348 338068 580412
rect 338132 580410 338138 580412
rect 341374 580410 341380 580412
rect 338132 580350 341380 580410
rect 338132 580348 338138 580350
rect 341374 580348 341380 580350
rect 341444 580348 341450 580412
rect 346894 580348 346900 580412
rect 346964 580410 346970 580412
rect 503897 580410 503963 580413
rect 346964 580408 503963 580410
rect 346964 580352 503902 580408
rect 503958 580352 503963 580408
rect 346964 580350 503963 580352
rect 346964 580348 346970 580350
rect 503897 580347 503963 580350
rect 91134 580212 91140 580276
rect 91204 580274 91210 580276
rect 321870 580274 321876 580276
rect 91204 580214 321876 580274
rect 91204 580212 91210 580214
rect 321870 580212 321876 580214
rect 321940 580212 321946 580276
rect 351678 580212 351684 580276
rect 351748 580274 351754 580276
rect 509969 580274 510035 580277
rect 351748 580272 510035 580274
rect 351748 580216 509974 580272
rect 510030 580216 510035 580272
rect 351748 580214 510035 580216
rect 351748 580212 351754 580214
rect 509969 580211 510035 580214
rect 91502 580076 91508 580140
rect 91572 580138 91578 580140
rect 93710 580138 93716 580140
rect 91572 580078 93716 580138
rect 91572 580076 91578 580078
rect 93710 580076 93716 580078
rect 93780 580076 93786 580140
rect 169702 580076 169708 580140
rect 169772 580138 169778 580140
rect 179270 580138 179276 580140
rect 169772 580078 179276 580138
rect 169772 580076 169778 580078
rect 179270 580076 179276 580078
rect 179340 580076 179346 580140
rect 318742 580076 318748 580140
rect 318812 580138 318818 580140
rect 328310 580138 328316 580140
rect 318812 580078 328316 580138
rect 318812 580076 318818 580078
rect 328310 580076 328316 580078
rect 328380 580076 328386 580140
rect 432086 580076 432092 580140
rect 432156 580138 432162 580140
rect 437422 580138 437428 580140
rect 432156 580078 437428 580138
rect 432156 580076 432162 580078
rect 437422 580076 437428 580078
rect 437492 580076 437498 580140
rect 456558 580076 456564 580140
rect 456628 580138 456634 580140
rect 456742 580138 456748 580140
rect 456628 580078 456748 580138
rect 456628 580076 456634 580078
rect 456742 580076 456748 580078
rect 456812 580076 456818 580140
rect 470726 580076 470732 580140
rect 470796 580138 470802 580140
rect 476062 580138 476068 580140
rect 470796 580078 476068 580138
rect 470796 580076 470802 580078
rect 476062 580076 476068 580078
rect 476132 580076 476138 580140
rect 491702 580076 491708 580140
rect 491772 580138 491778 580140
rect 511441 580138 511507 580141
rect 491772 580136 511507 580138
rect 491772 580080 511446 580136
rect 511502 580080 511507 580136
rect 491772 580078 511507 580080
rect 491772 580076 491778 580078
rect 511441 580075 511507 580078
rect 86718 579940 86724 580004
rect 86788 580002 86794 580004
rect 87638 580002 87644 580004
rect 86788 579942 87644 580002
rect 86788 579940 86794 579942
rect 87638 579940 87644 579942
rect 87708 579940 87714 580004
rect 88926 579940 88932 580004
rect 88996 580002 89002 580004
rect 94078 580002 94084 580004
rect 88996 579942 94084 580002
rect 88996 579940 89002 579942
rect 94078 579940 94084 579942
rect 94148 579940 94154 580004
rect 489862 579940 489868 580004
rect 489932 580002 489938 580004
rect 495382 580002 495388 580004
rect 489932 579942 495388 580002
rect 489932 579940 489938 579942
rect 495382 579940 495388 579942
rect 495452 579940 495458 580004
rect 90398 579866 90404 579868
rect 82494 579806 90404 579866
rect 90398 579804 90404 579806
rect 90468 579804 90474 579868
rect 92606 579804 92612 579868
rect 92676 579866 92682 579868
rect 97758 579866 97764 579868
rect 92676 579806 97764 579866
rect 92676 579804 92682 579806
rect 97758 579804 97764 579806
rect 97828 579804 97834 579868
rect 8753 579730 8819 579733
rect 503713 579730 503779 579733
rect 8753 579728 503779 579730
rect 8753 579672 8758 579728
rect 8814 579672 503718 579728
rect 503774 579672 503779 579728
rect 8753 579670 503779 579672
rect 8753 579667 8819 579670
rect 503713 579667 503779 579670
rect 532693 578234 532759 578237
rect 532877 578234 532943 578237
rect 532693 578232 532943 578234
rect 532693 578176 532698 578232
rect 532754 578176 532882 578232
rect 532938 578176 532943 578232
rect 532693 578174 532943 578176
rect 532693 578171 532759 578174
rect 532877 578171 532943 578174
rect 82629 577690 82695 577693
rect 508078 577690 508084 577692
rect 82629 577688 82738 577690
rect 82629 577632 82634 577688
rect 82690 577632 82738 577688
rect 82629 577627 82738 577632
rect 501860 577630 508084 577690
rect 508078 577628 508084 577630
rect 508148 577628 508154 577692
rect 82678 577116 82738 577627
rect 502701 575514 502767 575517
rect 506974 575514 506980 575516
rect 502701 575512 506980 575514
rect 502701 575456 502706 575512
rect 502762 575456 506980 575512
rect 502701 575454 506980 575456
rect 502701 575451 502767 575454
rect 506974 575452 506980 575454
rect 507044 575452 507050 575516
rect 503713 574154 503779 574157
rect 501860 574152 503779 574154
rect 501860 574096 503718 574152
rect 503774 574096 503779 574152
rect 501860 574094 503779 574096
rect 503713 574091 503779 574094
rect 501270 573684 501276 573748
rect 501340 573746 501346 573748
rect 502057 573746 502123 573749
rect 501340 573744 502123 573746
rect 501340 573688 502062 573744
rect 502118 573688 502123 573744
rect 501340 573686 502123 573688
rect 501340 573684 501346 573686
rect 502057 573683 502123 573686
rect 78673 573610 78739 573613
rect 78673 573608 82156 573610
rect 78673 573552 78678 573608
rect 78734 573552 82156 573608
rect 78673 573550 82156 573552
rect 78673 573547 78739 573550
rect 501270 573548 501276 573612
rect 501340 573610 501346 573612
rect 501822 573610 501828 573612
rect 501340 573550 501828 573610
rect 501340 573548 501346 573550
rect 501822 573548 501828 573550
rect 501892 573548 501898 573612
rect 501454 572188 501460 572252
rect 501524 572250 501530 572252
rect 502057 572250 502123 572253
rect 501524 572248 502123 572250
rect 501524 572192 502062 572248
rect 502118 572192 502123 572248
rect 501524 572190 502123 572192
rect 501524 572188 501530 572190
rect 502057 572187 502123 572190
rect 501454 571916 501460 571980
rect 501524 571978 501530 571980
rect 501822 571978 501828 571980
rect 501524 571918 501828 571978
rect 501524 571916 501530 571918
rect 501822 571916 501828 571918
rect 501892 571916 501898 571980
rect 79726 570012 79732 570076
rect 79796 570074 79802 570076
rect 501830 570074 501890 570588
rect 524413 570210 524479 570213
rect 524278 570208 524479 570210
rect 524278 570152 524418 570208
rect 524474 570152 524479 570208
rect 524278 570150 524479 570152
rect 505502 570074 505508 570076
rect 79796 570014 82156 570074
rect 501830 570014 505508 570074
rect 79796 570012 79802 570014
rect 505502 570012 505508 570014
rect 505572 570012 505578 570076
rect 524278 570074 524338 570150
rect 524413 570147 524479 570150
rect 524413 570074 524479 570077
rect 524278 570072 524479 570074
rect 524278 570016 524418 570072
rect 524474 570016 524479 570072
rect 524278 570014 524479 570016
rect 524413 570011 524479 570014
rect 583520 568836 584960 569076
rect 532417 568578 532483 568581
rect 532693 568578 532759 568581
rect 532417 568576 532759 568578
rect 532417 568520 532422 568576
rect 532478 568520 532698 568576
rect 532754 568520 532759 568576
rect 532417 568518 532759 568520
rect 532417 568515 532483 568518
rect 532693 568515 532759 568518
rect -960 567354 480 567444
rect 3509 567354 3575 567357
rect -960 567352 3575 567354
rect -960 567296 3514 567352
rect 3570 567296 3575 567352
rect -960 567294 3575 567296
rect -960 567204 480 567294
rect 3509 567291 3575 567294
rect 503805 567082 503871 567085
rect 501860 567080 503871 567082
rect 501860 567024 503810 567080
rect 503866 567024 503871 567080
rect 501860 567022 503871 567024
rect 503805 567019 503871 567022
rect 81617 566538 81683 566541
rect 81617 566536 82156 566538
rect 81617 566480 81622 566536
rect 81678 566480 82156 566536
rect 81617 566478 82156 566480
rect 81617 566475 81683 566478
rect 503805 563546 503871 563549
rect 501860 563544 503871 563546
rect 501860 563488 503810 563544
rect 503866 563488 503871 563544
rect 501860 563486 503871 563488
rect 503805 563483 503871 563486
rect 81341 563002 81407 563005
rect 81341 563000 82156 563002
rect 81341 562944 81346 563000
rect 81402 562944 82156 563000
rect 81341 562942 82156 562944
rect 81341 562939 81407 562942
rect 510102 560010 510108 560012
rect 501860 559950 510108 560010
rect 510102 559948 510108 559950
rect 510172 559948 510178 560012
rect 78673 559466 78739 559469
rect 78673 559464 82156 559466
rect 78673 559408 78678 559464
rect 78734 559408 82156 559464
rect 78673 559406 82156 559408
rect 78673 559403 78739 559406
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 501454 557092 501460 557156
rect 501524 557154 501530 557156
rect 502057 557154 502123 557157
rect 501524 557152 502123 557154
rect 501524 557096 502062 557152
rect 502118 557096 502123 557152
rect 583520 557140 584960 557230
rect 501524 557094 502123 557096
rect 501524 557092 501530 557094
rect 502057 557091 502123 557094
rect 501830 556202 501890 556444
rect 504909 556202 504975 556205
rect 501830 556200 504975 556202
rect 501830 556144 504914 556200
rect 504970 556144 504975 556200
rect 501830 556142 504975 556144
rect 504909 556139 504975 556142
rect 79542 555868 79548 555932
rect 79612 555930 79618 555932
rect 79612 555870 82156 555930
rect 79612 555868 79618 555870
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 82494 551852 82554 552364
rect 501830 552122 501890 552908
rect 504817 552122 504883 552125
rect 501830 552120 504883 552122
rect 501830 552064 504822 552120
rect 504878 552064 504883 552120
rect 501830 552062 504883 552064
rect 504817 552059 504883 552062
rect 82486 551788 82492 551852
rect 82556 551788 82562 551852
rect 505001 549402 505067 549405
rect 501860 549400 505067 549402
rect 501860 549344 505006 549400
rect 505062 549344 505067 549400
rect 501860 549342 505067 549344
rect 505001 549339 505067 549342
rect 79358 548796 79364 548860
rect 79428 548858 79434 548860
rect 79428 548798 82156 548858
rect 79428 548796 79434 548798
rect 501454 547844 501460 547908
rect 501524 547906 501530 547908
rect 502057 547906 502123 547909
rect 501524 547904 502123 547906
rect 501524 547848 502062 547904
rect 502118 547848 502123 547904
rect 501524 547846 502123 547848
rect 501524 547844 501530 547846
rect 502057 547843 502123 547846
rect 507894 545866 507900 545868
rect 501860 545806 507900 545866
rect 507894 545804 507900 545806
rect 507964 545804 507970 545868
rect 583520 545594 584960 545684
rect 583342 545534 584960 545594
rect 507158 545396 507164 545460
rect 507228 545458 507234 545460
rect 514661 545458 514727 545461
rect 507228 545456 514727 545458
rect 507228 545400 514666 545456
rect 514722 545400 514727 545456
rect 507228 545398 514727 545400
rect 507228 545396 507234 545398
rect 514661 545395 514727 545398
rect 531957 545458 532023 545461
rect 531957 545456 547890 545458
rect 531957 545400 531962 545456
rect 532018 545400 547890 545456
rect 531957 545398 547890 545400
rect 531957 545395 532023 545398
rect 81382 545260 81388 545324
rect 81452 545322 81458 545324
rect 514845 545322 514911 545325
rect 524321 545322 524387 545325
rect 81452 545262 82156 545322
rect 514845 545320 524387 545322
rect 514845 545264 514850 545320
rect 514906 545264 524326 545320
rect 524382 545264 524387 545320
rect 514845 545262 524387 545264
rect 547830 545322 547890 545398
rect 557582 545398 567210 545458
rect 547830 545262 557458 545322
rect 81452 545260 81458 545262
rect 514845 545259 514911 545262
rect 524321 545259 524387 545262
rect 524505 545186 524571 545189
rect 529933 545186 529999 545189
rect 524505 545184 529999 545186
rect 524505 545128 524510 545184
rect 524566 545128 529938 545184
rect 529994 545128 529999 545184
rect 524505 545126 529999 545128
rect 557398 545186 557458 545262
rect 557582 545186 557642 545398
rect 567150 545322 567210 545398
rect 583342 545322 583402 545534
rect 583520 545444 584960 545534
rect 567150 545262 576778 545322
rect 557398 545126 557642 545186
rect 576718 545186 576778 545262
rect 576902 545262 583402 545322
rect 576902 545186 576962 545262
rect 576718 545126 576962 545186
rect 524505 545123 524571 545126
rect 529933 545123 529999 545126
rect 506790 543900 506796 543964
rect 506860 543900 506866 543964
rect 506798 543692 506858 543900
rect 506790 543628 506796 543692
rect 506860 543628 506866 543692
rect 502558 542330 502564 542332
rect 501860 542270 502564 542330
rect 502558 542268 502564 542270
rect 502628 542268 502634 542332
rect 82678 541517 82738 541756
rect 82629 541512 82738 541517
rect 82629 541456 82634 541512
rect 82690 541456 82738 541512
rect 82629 541454 82738 541456
rect 82629 541451 82695 541454
rect 82118 539548 82124 539612
rect 82188 539610 82194 539612
rect 82624 539610 82630 539612
rect 82188 539550 82630 539610
rect 82188 539548 82194 539550
rect 82624 539548 82630 539550
rect 82694 539548 82700 539612
rect 506606 538794 506612 538796
rect -960 538658 480 538748
rect 501860 538734 506612 538794
rect 506606 538732 506612 538734
rect 506676 538732 506682 538796
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 81566 538188 81572 538252
rect 81636 538250 81642 538252
rect 81636 538190 82156 538250
rect 81636 538188 81642 538190
rect 79961 534714 80027 534717
rect 79961 534712 82156 534714
rect 79961 534656 79966 534712
rect 80022 534656 82156 534712
rect 79961 534654 82156 534656
rect 79961 534651 80027 534654
rect 501830 534578 501890 535228
rect 501830 534518 502074 534578
rect 502014 534170 502074 534518
rect 504449 534170 504515 534173
rect 502014 534168 504515 534170
rect 502014 534112 504454 534168
rect 504510 534112 504515 534168
rect 502014 534110 504515 534112
rect 504449 534107 504515 534110
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 501830 531450 501890 531692
rect 502926 531450 502932 531452
rect 501830 531390 502932 531450
rect 502926 531388 502932 531390
rect 502996 531388 503002 531452
rect 532693 531314 532759 531317
rect 532877 531314 532943 531317
rect 532693 531312 532943 531314
rect 532693 531256 532698 531312
rect 532754 531256 532882 531312
rect 532938 531256 532943 531312
rect 532693 531254 532943 531256
rect 532693 531251 532759 531254
rect 532877 531251 532943 531254
rect 81198 531116 81204 531180
rect 81268 531178 81274 531180
rect 81268 531118 82156 531178
rect 81268 531116 81274 531118
rect 505001 528186 505067 528189
rect 501860 528184 505067 528186
rect 501860 528128 505006 528184
rect 505062 528128 505067 528184
rect 501860 528126 505067 528128
rect 505001 528123 505067 528126
rect 81750 527580 81756 527644
rect 81820 527642 81826 527644
rect 81820 527582 82156 527642
rect 81820 527580 81826 527582
rect 504449 524650 504515 524653
rect 501860 524648 504515 524650
rect 501860 524592 504454 524648
rect 504510 524592 504515 524648
rect 501860 524590 504515 524592
rect 504449 524587 504515 524590
rect -960 524092 480 524332
rect 82494 523836 82554 524348
rect 82486 523772 82492 523836
rect 82556 523772 82562 523836
rect 583520 521916 584960 522156
rect 503805 521114 503871 521117
rect 501860 521112 503871 521114
rect 501860 521056 503810 521112
rect 503866 521056 503871 521112
rect 501860 521054 503871 521056
rect 503805 521051 503871 521054
rect 78673 520842 78739 520845
rect 78673 520840 82156 520842
rect 78673 520784 78678 520840
rect 78734 520784 82156 520840
rect 78673 520782 82156 520784
rect 78673 520779 78739 520782
rect 501638 520162 501644 520164
rect 501462 520102 501644 520162
rect 501462 519618 501522 520102
rect 501638 520100 501644 520102
rect 501708 520100 501714 520164
rect 501638 519618 501644 519620
rect 501462 519558 501644 519618
rect 501638 519556 501644 519558
rect 501708 519556 501714 519620
rect 82486 519284 82492 519348
rect 82556 519284 82562 519348
rect 82494 519076 82554 519284
rect 82486 519012 82492 519076
rect 82556 519012 82562 519076
rect 82353 518802 82419 518805
rect 82486 518802 82492 518804
rect 82353 518800 82492 518802
rect 82353 518744 82358 518800
rect 82414 518744 82492 518800
rect 82353 518742 82492 518744
rect 82353 518739 82419 518742
rect 82486 518740 82492 518742
rect 82556 518740 82562 518804
rect 501781 518122 501847 518125
rect 501781 518120 501890 518122
rect 501781 518064 501786 518120
rect 501842 518064 501890 518120
rect 501781 518059 501890 518064
rect 501830 517548 501890 518059
rect 81801 517306 81867 517309
rect 81801 517304 82156 517306
rect 81801 517248 81806 517304
rect 81862 517248 82156 517304
rect 81801 517246 82156 517248
rect 81801 517243 81867 517246
rect 501270 517244 501276 517308
rect 501340 517306 501346 517308
rect 501781 517306 501847 517309
rect 501340 517304 501847 517306
rect 501340 517248 501786 517304
rect 501842 517248 501847 517304
rect 501340 517246 501847 517248
rect 501340 517244 501346 517246
rect 501781 517243 501847 517246
rect 502006 517244 502012 517308
rect 502076 517306 502082 517308
rect 502190 517306 502196 517308
rect 502076 517246 502196 517306
rect 502076 517244 502082 517246
rect 502190 517244 502196 517246
rect 502260 517244 502266 517308
rect 74441 513770 74507 513773
rect 501278 513772 501338 514012
rect 74441 513768 82156 513770
rect 74441 513712 74446 513768
rect 74502 513712 82156 513768
rect 74441 513710 82156 513712
rect 74441 513707 74507 513710
rect 501270 513708 501276 513772
rect 501340 513708 501346 513772
rect 501270 511940 501276 512004
rect 501340 512002 501346 512004
rect 502006 512002 502012 512004
rect 501340 511942 502012 512002
rect 501340 511940 501346 511942
rect 502006 511940 502012 511942
rect 502076 511940 502082 512004
rect 532693 512002 532759 512005
rect 532877 512002 532943 512005
rect 532693 512000 532943 512002
rect 532693 511944 532698 512000
rect 532754 511944 532882 512000
rect 532938 511944 532943 512000
rect 532693 511942 532943 511944
rect 532693 511939 532759 511942
rect 532877 511939 532943 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 77150 510172 77156 510236
rect 77220 510234 77226 510236
rect 77220 510174 82156 510234
rect 583520 510220 584960 510310
rect 77220 510172 77226 510174
rect -960 509962 480 510052
rect 2865 509962 2931 509965
rect -960 509960 2931 509962
rect -960 509904 2870 509960
rect 2926 509904 2931 509960
rect -960 509902 2931 509904
rect -960 509812 480 509902
rect 2865 509899 2931 509902
rect 82353 509556 82419 509557
rect 82302 509554 82308 509556
rect 82262 509494 82308 509554
rect 82372 509552 82419 509556
rect 82414 509496 82419 509552
rect 82302 509492 82308 509494
rect 82372 509492 82419 509496
rect 82353 509491 82419 509492
rect 504214 507242 504220 507244
rect 501860 507182 504220 507242
rect 504214 507180 504220 507182
rect 504284 507180 504290 507244
rect 501270 506908 501276 506972
rect 501340 506970 501346 506972
rect 501781 506970 501847 506973
rect 501340 506968 501847 506970
rect 501340 506912 501786 506968
rect 501842 506912 501847 506968
rect 501340 506910 501847 506912
rect 501340 506908 501346 506910
rect 501781 506907 501847 506910
rect 501822 506772 501828 506836
rect 501892 506834 501898 506836
rect 502190 506834 502196 506836
rect 501892 506774 502196 506834
rect 501892 506772 501898 506774
rect 502190 506772 502196 506774
rect 502260 506772 502266 506836
rect 78121 506698 78187 506701
rect 78121 506696 82156 506698
rect 78121 506640 78126 506696
rect 78182 506640 82156 506696
rect 78121 506638 82156 506640
rect 78121 506635 78187 506638
rect 82537 505748 82603 505749
rect 82486 505746 82492 505748
rect 82446 505686 82492 505746
rect 82556 505744 82603 505748
rect 82598 505688 82603 505744
rect 82486 505684 82492 505686
rect 82556 505684 82603 505688
rect 82537 505683 82603 505684
rect 502374 503706 502380 503708
rect 501860 503646 502380 503706
rect 502374 503644 502380 503646
rect 502444 503644 502450 503708
rect 74349 503162 74415 503165
rect 74349 503160 82156 503162
rect 74349 503104 74354 503160
rect 74410 503104 82156 503160
rect 74349 503102 82156 503104
rect 74349 503099 74415 503102
rect 82353 500852 82419 500853
rect 82302 500788 82308 500852
rect 82372 500850 82419 500852
rect 82372 500848 82464 500850
rect 82414 500792 82464 500848
rect 82372 500790 82464 500792
rect 82372 500788 82419 500790
rect 501822 500788 501828 500852
rect 501892 500788 501898 500852
rect 82353 500787 82419 500788
rect 501830 500578 501890 500788
rect 502057 500578 502123 500581
rect 501830 500576 502123 500578
rect 501830 500520 502062 500576
rect 502118 500520 502123 500576
rect 501830 500518 502123 500520
rect 502057 500515 502123 500518
rect 504173 500170 504239 500173
rect 501860 500168 504239 500170
rect 501860 500112 504178 500168
rect 504234 500112 504239 500168
rect 501860 500110 504239 500112
rect 504173 500107 504239 500110
rect 78029 499626 78095 499629
rect 78029 499624 82156 499626
rect 78029 499568 78034 499624
rect 78090 499568 82156 499624
rect 78029 499566 82156 499568
rect 78029 499563 78095 499566
rect 579981 498674 580047 498677
rect 583520 498674 584960 498764
rect 579981 498672 584960 498674
rect 579981 498616 579986 498672
rect 580042 498616 584960 498672
rect 579981 498614 584960 498616
rect 579981 498611 580047 498614
rect 583520 498524 584960 498614
rect 82302 498068 82308 498132
rect 82372 498130 82378 498132
rect 82537 498130 82603 498133
rect 82372 498128 82603 498130
rect 82372 498072 82542 498128
rect 82598 498072 82603 498128
rect 82372 498070 82603 498072
rect 82372 498068 82378 498070
rect 82537 498067 82603 498070
rect 82353 497180 82419 497181
rect 82302 497178 82308 497180
rect 82262 497118 82308 497178
rect 82372 497176 82419 497180
rect 82414 497120 82419 497176
rect 82302 497116 82308 497118
rect 82372 497116 82419 497120
rect 82353 497115 82419 497116
rect 504449 496634 504515 496637
rect 501860 496632 504515 496634
rect 501860 496576 504454 496632
rect 504510 496576 504515 496632
rect 501860 496574 504515 496576
rect 504449 496571 504515 496574
rect 82126 495820 82186 496060
rect 82118 495756 82124 495820
rect 82188 495756 82194 495820
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 501822 493308 501828 493372
rect 501892 493370 501898 493372
rect 502057 493370 502123 493373
rect 501892 493368 502123 493370
rect 501892 493312 502062 493368
rect 502118 493312 502123 493368
rect 501892 493310 502123 493312
rect 501892 493308 501898 493310
rect 502057 493307 502123 493310
rect 501830 492690 501890 493068
rect 505001 492690 505067 492693
rect 501830 492688 505067 492690
rect 501830 492632 505006 492688
rect 505062 492632 505067 492688
rect 501830 492630 505067 492632
rect 505001 492627 505067 492630
rect 506790 492628 506796 492692
rect 506860 492690 506866 492692
rect 506974 492690 506980 492692
rect 506860 492630 506980 492690
rect 506860 492628 506866 492630
rect 506974 492628 506980 492630
rect 507044 492628 507050 492692
rect 81934 491948 81940 492012
rect 82004 492010 82010 492012
rect 82126 492010 82186 492524
rect 82004 491950 82186 492010
rect 82004 491948 82010 491950
rect 505185 489562 505251 489565
rect 501860 489560 505251 489562
rect 501860 489504 505190 489560
rect 505246 489504 505251 489560
rect 501860 489502 505251 489504
rect 505185 489499 505251 489502
rect 81157 489018 81223 489021
rect 81157 489016 82156 489018
rect 81157 488960 81162 489016
rect 81218 488960 82156 489016
rect 81157 488958 82156 488960
rect 81157 488955 81223 488958
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 82537 486164 82603 486165
rect 82486 486100 82492 486164
rect 82556 486162 82603 486164
rect 82556 486160 82648 486162
rect 82598 486104 82648 486160
rect 82556 486102 82648 486104
rect 82556 486100 82603 486102
rect 82537 486099 82603 486100
rect 508262 486026 508268 486028
rect 501860 485966 508268 486026
rect 508262 485964 508268 485966
rect 508332 485964 508338 486028
rect 82494 484940 82554 485452
rect 82486 484876 82492 484940
rect 82556 484876 82562 484940
rect 532693 483034 532759 483037
rect 532877 483034 532943 483037
rect 532693 483032 532943 483034
rect 532693 482976 532698 483032
rect 532754 482976 532882 483032
rect 532938 482976 532943 483032
rect 532693 482974 532943 482976
rect 532693 482971 532759 482974
rect 532877 482971 532943 482974
rect 503897 482490 503963 482493
rect 501860 482488 503963 482490
rect 501860 482432 503902 482488
rect 503958 482432 503963 482488
rect 501860 482430 503963 482432
rect 503897 482427 503963 482430
rect 79869 481946 79935 481949
rect 79869 481944 82156 481946
rect 79869 481888 79874 481944
rect 79930 481888 82156 481944
rect 79869 481886 82156 481888
rect 79869 481883 79935 481886
rect 82353 481266 82419 481269
rect 82486 481266 82492 481268
rect 82353 481264 82492 481266
rect -960 481130 480 481220
rect 82353 481208 82358 481264
rect 82414 481208 82492 481264
rect 82353 481206 82492 481208
rect 82353 481203 82419 481206
rect 82486 481204 82492 481206
rect 82556 481204 82562 481268
rect 3325 481130 3391 481133
rect 82537 481132 82603 481133
rect -960 481128 3391 481130
rect -960 481072 3330 481128
rect 3386 481072 3391 481128
rect -960 481070 3391 481072
rect -960 480980 480 481070
rect 3325 481067 3391 481070
rect 82486 481068 82492 481132
rect 82556 481130 82603 481132
rect 82556 481128 82648 481130
rect 82598 481072 82648 481128
rect 82556 481070 82648 481072
rect 82556 481068 82603 481070
rect 82537 481067 82603 481068
rect 505001 478954 505067 478957
rect 501860 478952 505067 478954
rect 501860 478896 505006 478952
rect 505062 478896 505067 478952
rect 501860 478894 505067 478896
rect 505001 478891 505067 478894
rect 501822 478620 501828 478684
rect 501892 478682 501898 478684
rect 502006 478682 502012 478684
rect 501892 478622 502012 478682
rect 501892 478620 501898 478622
rect 502006 478620 502012 478622
rect 502076 478620 502082 478684
rect 77569 478410 77635 478413
rect 77569 478408 82156 478410
rect 77569 478352 77574 478408
rect 77630 478352 82156 478408
rect 77569 478350 82156 478352
rect 77569 478347 77635 478350
rect 82537 475828 82603 475829
rect 82486 475764 82492 475828
rect 82556 475826 82603 475828
rect 82556 475824 82648 475826
rect 82598 475768 82648 475824
rect 82556 475766 82648 475768
rect 82556 475764 82603 475766
rect 82537 475763 82603 475764
rect 503662 475418 503668 475420
rect 501860 475358 503668 475418
rect 503662 475356 503668 475358
rect 503732 475356 503738 475420
rect 583520 474996 584960 475236
rect 82678 474333 82738 474844
rect 501270 474812 501276 474876
rect 501340 474874 501346 474876
rect 501781 474874 501847 474877
rect 501340 474872 501847 474874
rect 501340 474816 501786 474872
rect 501842 474816 501847 474872
rect 501340 474814 501847 474816
rect 501340 474812 501346 474814
rect 501781 474811 501847 474814
rect 82629 474328 82738 474333
rect 82629 474272 82634 474328
rect 82690 474272 82738 474328
rect 82629 474270 82738 474272
rect 82629 474267 82695 474270
rect 82445 474196 82511 474197
rect 82445 474194 82492 474196
rect 82400 474192 82492 474194
rect 82400 474136 82450 474192
rect 82400 474134 82492 474136
rect 82445 474132 82492 474134
rect 82556 474132 82562 474196
rect 82445 474131 82511 474132
rect 82353 473650 82419 473653
rect 82486 473650 82492 473652
rect 82353 473648 82492 473650
rect 82353 473592 82358 473648
rect 82414 473592 82492 473648
rect 82353 473590 82492 473592
rect 82353 473587 82419 473590
rect 82486 473588 82492 473590
rect 82556 473588 82562 473652
rect 82537 473516 82603 473517
rect 82486 473514 82492 473516
rect 82446 473454 82492 473514
rect 82556 473512 82603 473516
rect 82598 473456 82603 473512
rect 82486 473452 82492 473454
rect 82556 473452 82603 473456
rect 82537 473451 82603 473452
rect 503529 471882 503595 471885
rect 501860 471880 503595 471882
rect 501860 471824 503534 471880
rect 503590 471824 503595 471880
rect 501860 471822 503595 471824
rect 503529 471819 503595 471822
rect 80973 471338 81039 471341
rect 80973 471336 82156 471338
rect 80973 471280 80978 471336
rect 81034 471280 82156 471336
rect 80973 471278 82156 471280
rect 80973 471275 81039 471278
rect 82537 471068 82603 471069
rect 82486 471066 82492 471068
rect 82446 471006 82492 471066
rect 82556 471064 82603 471068
rect 82598 471008 82603 471064
rect 82486 471004 82492 471006
rect 82556 471004 82603 471008
rect 82537 471003 82603 471004
rect 501830 467938 501890 468316
rect 509734 467938 509740 467940
rect 501830 467878 509740 467938
rect 509734 467876 509740 467878
rect 509804 467876 509810 467940
rect 81985 467258 82051 467261
rect 82126 467258 82186 467772
rect 81985 467256 82186 467258
rect 81985 467200 81990 467256
rect 82046 467200 82186 467256
rect 81985 467198 82186 467200
rect 81985 467195 82051 467198
rect -960 466700 480 466940
rect 82445 466172 82511 466173
rect 82445 466170 82492 466172
rect 82400 466168 82492 466170
rect 82400 466112 82450 466168
rect 82400 466110 82492 466112
rect 82445 466108 82492 466110
rect 82556 466108 82562 466172
rect 82445 466107 82511 466108
rect 506790 464810 506796 464812
rect 501860 464750 506796 464810
rect 506790 464748 506796 464750
rect 506860 464748 506866 464812
rect 501454 464476 501460 464540
rect 501524 464538 501530 464540
rect 502190 464538 502196 464540
rect 501524 464478 502196 464538
rect 501524 464476 501530 464478
rect 502190 464476 502196 464478
rect 502260 464476 502266 464540
rect 501638 464340 501644 464404
rect 501708 464402 501714 464404
rect 502149 464402 502215 464405
rect 501708 464400 502215 464402
rect 501708 464344 502154 464400
rect 502210 464344 502215 464400
rect 501708 464342 502215 464344
rect 501708 464340 501714 464342
rect 502149 464339 502215 464342
rect 81065 464266 81131 464269
rect 81065 464264 82156 464266
rect 81065 464208 81070 464264
rect 81126 464208 82156 464264
rect 81065 464206 82156 464208
rect 81065 464203 81131 464206
rect 501454 464204 501460 464268
rect 501524 464266 501530 464268
rect 501781 464266 501847 464269
rect 501524 464264 501847 464266
rect 501524 464208 501786 464264
rect 501842 464208 501847 464264
rect 501524 464206 501847 464208
rect 501524 464204 501530 464206
rect 501781 464203 501847 464206
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 502742 461274 502748 461276
rect 501860 461214 502748 461274
rect 502742 461212 502748 461214
rect 502812 461212 502818 461276
rect 80881 460730 80947 460733
rect 80881 460728 82156 460730
rect 80881 460672 80886 460728
rect 80942 460672 82156 460728
rect 80881 460670 82156 460672
rect 80881 460667 80947 460670
rect 82537 458012 82603 458013
rect 82486 457948 82492 458012
rect 82556 458010 82603 458012
rect 82556 458008 82648 458010
rect 82598 457952 82648 458008
rect 82556 457950 82648 457952
rect 82556 457948 82603 457950
rect 82537 457947 82603 457948
rect 82310 456924 82370 457436
rect 501830 457197 501890 457708
rect 501781 457192 501890 457197
rect 501781 457136 501786 457192
rect 501842 457136 501890 457192
rect 501781 457134 501890 457136
rect 501781 457131 501847 457134
rect 82302 456860 82308 456924
rect 82372 456860 82378 456924
rect 101581 456516 101647 456517
rect 101581 456514 101628 456516
rect 101536 456512 101628 456514
rect 101536 456456 101586 456512
rect 101536 456454 101628 456456
rect 101581 456452 101628 456454
rect 101692 456452 101698 456516
rect 101581 456451 101647 456452
rect 501638 454820 501644 454884
rect 501708 454882 501714 454884
rect 502149 454882 502215 454885
rect 501708 454880 502215 454882
rect 501708 454824 502154 454880
rect 502210 454824 502215 454880
rect 501708 454822 502215 454824
rect 501708 454820 501714 454822
rect 502149 454819 502215 454822
rect 502057 454748 502123 454749
rect 502006 454746 502012 454748
rect 501966 454686 502012 454746
rect 502076 454744 502123 454748
rect 502118 454688 502123 454744
rect 502006 454684 502012 454686
rect 502076 454684 502123 454688
rect 502057 454683 502123 454684
rect 504541 454202 504607 454205
rect 501860 454200 504607 454202
rect 501860 454144 504546 454200
rect 504602 454144 504607 454200
rect 501860 454142 504607 454144
rect 504541 454139 504607 454142
rect 82678 453389 82738 453900
rect 82629 453384 82738 453389
rect 82629 453328 82634 453384
rect 82690 453328 82738 453384
rect 82629 453326 82738 453328
rect 82629 453323 82695 453326
rect -960 452434 480 452524
rect 3918 452434 3924 452436
rect -960 452374 3924 452434
rect -960 452284 480 452374
rect 3918 452372 3924 452374
rect 3988 452372 3994 452436
rect 101489 451892 101555 451893
rect 101438 451828 101444 451892
rect 101508 451890 101555 451892
rect 101508 451888 101600 451890
rect 101550 451832 101600 451888
rect 101508 451830 101600 451832
rect 101508 451828 101555 451830
rect 101489 451827 101555 451828
rect 580441 451754 580507 451757
rect 583520 451754 584960 451844
rect 580441 451752 584960 451754
rect 580441 451696 580446 451752
rect 580502 451696 584960 451752
rect 580441 451694 584960 451696
rect 580441 451691 580507 451694
rect 583520 451604 584960 451694
rect 503662 450666 503668 450668
rect 501860 450606 503668 450666
rect 503662 450604 503668 450606
rect 503732 450604 503738 450668
rect 76833 450394 76899 450397
rect 76833 450392 82156 450394
rect 76833 450336 76838 450392
rect 76894 450336 82156 450392
rect 76833 450334 82156 450336
rect 76833 450331 76899 450334
rect 502057 449034 502123 449037
rect 502190 449034 502196 449036
rect 502057 449032 502196 449034
rect 502057 448976 502062 449032
rect 502118 448976 502196 449032
rect 502057 448974 502196 448976
rect 502057 448971 502123 448974
rect 502190 448972 502196 448974
rect 502260 448972 502266 449036
rect 504582 447130 504588 447132
rect 501860 447070 504588 447130
rect 504582 447068 504588 447070
rect 504652 447068 504658 447132
rect 79685 446858 79751 446861
rect 79685 446856 82156 446858
rect 79685 446800 79690 446856
rect 79746 446800 82156 446856
rect 79685 446798 82156 446800
rect 79685 446795 79751 446798
rect 507158 444484 507164 444548
rect 507228 444484 507234 444548
rect 507166 444412 507226 444484
rect 507158 444348 507164 444412
rect 507228 444348 507234 444412
rect 80789 443322 80855 443325
rect 501462 443324 501522 443836
rect 80789 443320 82156 443322
rect 80789 443264 80794 443320
rect 80850 443264 82156 443320
rect 80789 443262 82156 443264
rect 80789 443259 80855 443262
rect 501454 443260 501460 443324
rect 501524 443260 501530 443324
rect 501270 442444 501276 442508
rect 501340 442444 501346 442508
rect 501454 442444 501460 442508
rect 501524 442506 501530 442508
rect 501965 442506 502031 442509
rect 501524 442504 502031 442506
rect 501524 442448 501970 442504
rect 502026 442448 502031 442504
rect 501524 442446 502031 442448
rect 501524 442444 501530 442446
rect 501278 442234 501338 442444
rect 501965 442443 502031 442446
rect 501454 442234 501460 442236
rect 501278 442174 501460 442234
rect 501454 442172 501460 442174
rect 501524 442172 501530 442236
rect 503989 440330 504055 440333
rect 501860 440328 504055 440330
rect 501860 440272 503994 440328
rect 504050 440272 504055 440328
rect 501860 440270 504055 440272
rect 503989 440267 504055 440270
rect 579981 439922 580047 439925
rect 583520 439922 584960 440012
rect 579981 439920 584960 439922
rect 579981 439864 579986 439920
rect 580042 439864 584960 439920
rect 579981 439862 584960 439864
rect 579981 439859 580047 439862
rect 80697 439786 80763 439789
rect 80697 439784 82156 439786
rect 80697 439728 80702 439784
rect 80758 439728 82156 439784
rect 80697 439726 82156 439728
rect 80697 439723 80763 439726
rect 501270 439724 501276 439788
rect 501340 439786 501346 439788
rect 501965 439786 502031 439789
rect 501340 439784 502031 439786
rect 501340 439728 501970 439784
rect 502026 439728 502031 439784
rect 583520 439772 584960 439862
rect 501340 439726 502031 439728
rect 501340 439724 501346 439726
rect 501965 439723 502031 439726
rect 82537 438972 82603 438973
rect 82486 438908 82492 438972
rect 82556 438970 82603 438972
rect 82556 438968 82648 438970
rect 82598 438912 82648 438968
rect 82556 438910 82648 438912
rect 82556 438908 82603 438910
rect 82537 438907 82603 438908
rect -960 438018 480 438108
rect 501454 438092 501460 438156
rect 501524 438154 501530 438156
rect 502006 438154 502012 438156
rect 501524 438094 502012 438154
rect 501524 438092 501530 438094
rect 502006 438092 502012 438094
rect 502076 438092 502082 438156
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 504081 436794 504147 436797
rect 501860 436792 504147 436794
rect 501860 436736 504086 436792
rect 504142 436736 504147 436792
rect 501860 436734 504147 436736
rect 504081 436731 504147 436734
rect 75085 436250 75151 436253
rect 75085 436248 82156 436250
rect 75085 436192 75090 436248
rect 75146 436192 82156 436248
rect 75085 436190 82156 436192
rect 75085 436187 75151 436190
rect 82537 435436 82603 435437
rect 82486 435434 82492 435436
rect 82446 435374 82492 435434
rect 82556 435432 82603 435436
rect 82598 435376 82603 435432
rect 82486 435372 82492 435374
rect 82556 435372 82603 435376
rect 82537 435371 82603 435372
rect 507025 434620 507091 434621
rect 506974 434556 506980 434620
rect 507044 434618 507091 434620
rect 507044 434616 507136 434618
rect 507086 434560 507136 434616
rect 507044 434558 507136 434560
rect 507044 434556 507091 434558
rect 507025 434555 507091 434556
rect 502885 433258 502951 433261
rect 501860 433256 502951 433258
rect 501860 433200 502890 433256
rect 502946 433200 502951 433256
rect 501860 433198 502951 433200
rect 502885 433195 502951 433198
rect 79174 432652 79180 432716
rect 79244 432714 79250 432716
rect 79244 432654 82156 432714
rect 79244 432652 79250 432654
rect 82537 431220 82603 431221
rect 82486 431218 82492 431220
rect 82446 431158 82492 431218
rect 82556 431216 82603 431220
rect 82598 431160 82603 431216
rect 82486 431156 82492 431158
rect 82556 431156 82603 431160
rect 82537 431155 82603 431156
rect 505553 429722 505619 429725
rect 501860 429720 505619 429722
rect 501860 429664 505558 429720
rect 505614 429664 505619 429720
rect 501860 429662 505619 429664
rect 505553 429659 505619 429662
rect 77569 429178 77635 429181
rect 77569 429176 82156 429178
rect 77569 429120 77574 429176
rect 77630 429120 82156 429176
rect 77569 429118 82156 429120
rect 77569 429115 77635 429118
rect 583520 428076 584960 428316
rect 504214 427892 504220 427956
rect 504284 427892 504290 427956
rect 501270 427756 501276 427820
rect 501340 427818 501346 427820
rect 502149 427818 502215 427821
rect 501340 427816 502215 427818
rect 501340 427760 502154 427816
rect 502210 427760 502215 427816
rect 501340 427758 502215 427760
rect 501340 427756 501346 427758
rect 502149 427755 502215 427758
rect 504222 427684 504282 427892
rect 504214 427620 504220 427684
rect 504284 427620 504290 427684
rect 504633 426186 504699 426189
rect 501860 426184 504699 426186
rect 501860 426128 504638 426184
rect 504694 426128 504699 426184
rect 501860 426126 504699 426128
rect 504633 426123 504699 426126
rect 81249 425642 81315 425645
rect 81249 425640 82156 425642
rect 81249 425584 81254 425640
rect 81310 425584 82156 425640
rect 81249 425582 82156 425584
rect 81249 425579 81315 425582
rect 506790 425444 506796 425508
rect 506860 425444 506866 425508
rect 502885 425098 502951 425101
rect 506798 425100 506858 425444
rect 507025 425236 507091 425237
rect 506974 425234 506980 425236
rect 506934 425174 506980 425234
rect 507044 425232 507091 425236
rect 507086 425176 507091 425232
rect 506974 425172 506980 425174
rect 507044 425172 507091 425176
rect 507158 425172 507164 425236
rect 507228 425172 507234 425236
rect 507025 425171 507091 425172
rect 507166 425100 507226 425172
rect 504398 425098 504404 425100
rect 502885 425096 504404 425098
rect 502885 425040 502890 425096
rect 502946 425040 504404 425096
rect 502885 425038 504404 425040
rect 502885 425035 502951 425038
rect 504398 425036 504404 425038
rect 504468 425036 504474 425100
rect 506790 425036 506796 425100
rect 506860 425036 506866 425100
rect 507158 425036 507164 425100
rect 507228 425036 507234 425100
rect 502006 423874 502012 423876
rect -960 423738 480 423828
rect 501830 423814 502012 423874
rect 2957 423738 3023 423741
rect 501830 423740 501890 423814
rect 502006 423812 502012 423814
rect 502076 423812 502082 423876
rect -960 423736 3023 423738
rect -960 423680 2962 423736
rect 3018 423680 3023 423736
rect -960 423678 3023 423680
rect -960 423588 480 423678
rect 2957 423675 3023 423678
rect 501822 423676 501828 423740
rect 501892 423676 501898 423740
rect 501822 423404 501828 423468
rect 501892 423466 501898 423468
rect 502057 423466 502123 423469
rect 501892 423464 502123 423466
rect 501892 423408 502062 423464
rect 502118 423408 502123 423464
rect 501892 423406 502123 423408
rect 501892 423404 501898 423406
rect 502057 423403 502123 423406
rect 507710 422650 507716 422652
rect 501860 422590 507716 422650
rect 507710 422588 507716 422590
rect 507780 422588 507786 422652
rect 78990 422044 78996 422108
rect 79060 422106 79066 422108
rect 79060 422046 82156 422106
rect 79060 422044 79066 422046
rect 503253 419114 503319 419117
rect 501860 419112 503319 419114
rect 501860 419056 503258 419112
rect 503314 419056 503319 419112
rect 501860 419054 503319 419056
rect 503253 419051 503319 419054
rect 76741 418570 76807 418573
rect 76741 418568 82156 418570
rect 76741 418512 76746 418568
rect 76802 418512 82156 418568
rect 76741 418510 82156 418512
rect 76741 418507 76807 418510
rect 501270 418236 501276 418300
rect 501340 418298 501346 418300
rect 502149 418298 502215 418301
rect 501340 418296 502215 418298
rect 501340 418240 502154 418296
rect 502210 418240 502215 418296
rect 501340 418238 502215 418240
rect 501340 418236 501346 418238
rect 502149 418235 502215 418238
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 502425 415578 502491 415581
rect 501860 415576 502491 415578
rect 501860 415520 502430 415576
rect 502486 415520 502491 415576
rect 501860 415518 502491 415520
rect 502425 415515 502491 415518
rect 81709 415034 81775 415037
rect 81709 415032 82156 415034
rect 81709 414976 81714 415032
rect 81770 414976 82156 415032
rect 81709 414974 82156 414976
rect 81709 414971 81775 414974
rect 502057 414084 502123 414085
rect 502006 414020 502012 414084
rect 502076 414082 502123 414084
rect 502076 414080 502168 414082
rect 502118 414024 502168 414080
rect 502076 414022 502168 414024
rect 502076 414020 502123 414022
rect 502057 414019 502123 414020
rect 502057 413810 502123 413813
rect 502190 413810 502196 413812
rect 502057 413808 502196 413810
rect 502057 413752 502062 413808
rect 502118 413752 502196 413808
rect 502057 413750 502196 413752
rect 502057 413747 502123 413750
rect 502190 413748 502196 413750
rect 502260 413748 502266 413812
rect 505645 412042 505711 412045
rect 501860 412040 505711 412042
rect 501860 411984 505650 412040
rect 505706 411984 505711 412040
rect 501860 411982 505711 411984
rect 505645 411979 505711 411982
rect 79409 411498 79475 411501
rect 79409 411496 82156 411498
rect 79409 411440 79414 411496
rect 79470 411440 82156 411496
rect 79409 411438 82156 411440
rect 79409 411435 79475 411438
rect 501270 411436 501276 411500
rect 501340 411498 501346 411500
rect 501965 411498 502031 411501
rect 501340 411496 502031 411498
rect 501340 411440 501970 411496
rect 502026 411440 502031 411496
rect 501340 411438 502031 411440
rect 501340 411436 501346 411438
rect 501965 411435 502031 411438
rect 501965 410138 502031 410141
rect 501278 410136 502031 410138
rect 501278 410080 501970 410136
rect 502026 410080 502031 410136
rect 501278 410078 502031 410080
rect 501278 410004 501338 410078
rect 501965 410075 502031 410078
rect 501270 409940 501276 410004
rect 501340 409940 501346 410004
rect -960 409172 480 409412
rect 504030 408580 504036 408644
rect 504100 408642 504106 408644
rect 504398 408642 504404 408644
rect 504100 408582 504404 408642
rect 504100 408580 504106 408582
rect 504398 408580 504404 408582
rect 504468 408580 504474 408644
rect 503846 408506 503852 408508
rect 501860 408446 503852 408506
rect 503846 408444 503852 408446
rect 503916 408444 503922 408508
rect 77661 407962 77727 407965
rect 77661 407960 82156 407962
rect 77661 407904 77666 407960
rect 77722 407904 82156 407960
rect 77661 407902 82156 407904
rect 77661 407899 77727 407902
rect 82537 406468 82603 406469
rect 82486 406466 82492 406468
rect 82446 406406 82492 406466
rect 82556 406464 82603 406468
rect 82598 406408 82603 406464
rect 82486 406404 82492 406406
rect 82556 406404 82603 406408
rect 82537 406403 82603 406404
rect 501822 405724 501828 405788
rect 501892 405786 501898 405788
rect 501965 405786 502031 405789
rect 501892 405784 502031 405786
rect 501892 405728 501970 405784
rect 502026 405728 502031 405784
rect 501892 405726 502031 405728
rect 501892 405724 501898 405726
rect 501965 405723 502031 405726
rect 501822 405588 501828 405652
rect 501892 405650 501898 405652
rect 502057 405650 502123 405653
rect 507025 405652 507091 405653
rect 501892 405648 502123 405650
rect 501892 405592 502062 405648
rect 502118 405592 502123 405648
rect 501892 405590 502123 405592
rect 501892 405588 501898 405590
rect 502057 405587 502123 405590
rect 506974 405588 506980 405652
rect 507044 405650 507091 405652
rect 507044 405648 507136 405650
rect 507086 405592 507136 405648
rect 507044 405590 507136 405592
rect 507044 405588 507091 405590
rect 507025 405587 507091 405588
rect 505001 404970 505067 404973
rect 501860 404968 505067 404970
rect 501860 404912 505006 404968
rect 505062 404912 505067 404968
rect 501860 404910 505067 404912
rect 505001 404907 505067 404910
rect 580441 404834 580507 404837
rect 583520 404834 584960 404924
rect 580441 404832 584960 404834
rect 580441 404776 580446 404832
rect 580502 404776 584960 404832
rect 580441 404774 584960 404776
rect 580441 404771 580507 404774
rect 583520 404684 584960 404774
rect 80605 404426 80671 404429
rect 80605 404424 82156 404426
rect 80605 404368 80610 404424
rect 80666 404368 82156 404424
rect 80605 404366 82156 404368
rect 80605 404363 80671 404366
rect 501454 403684 501460 403748
rect 501524 403746 501530 403748
rect 502057 403746 502123 403749
rect 501524 403744 502123 403746
rect 501524 403688 502062 403744
rect 502118 403688 502123 403744
rect 501524 403686 502123 403688
rect 501524 403684 501530 403686
rect 502057 403683 502123 403686
rect 82537 401572 82603 401573
rect 82486 401570 82492 401572
rect 82446 401510 82492 401570
rect 82556 401568 82603 401572
rect 82598 401512 82603 401568
rect 82486 401508 82492 401510
rect 82556 401508 82603 401512
rect 82537 401507 82603 401508
rect 502609 401434 502675 401437
rect 501860 401432 502675 401434
rect 501860 401376 502614 401432
rect 502670 401376 502675 401432
rect 501860 401374 502675 401376
rect 502609 401371 502675 401374
rect 78765 400890 78831 400893
rect 78765 400888 82156 400890
rect 78765 400832 78770 400888
rect 78826 400832 82156 400888
rect 78765 400830 82156 400832
rect 78765 400827 78831 400830
rect 501822 400828 501828 400892
rect 501892 400890 501898 400892
rect 502190 400890 502196 400892
rect 501892 400830 502196 400890
rect 501892 400828 501898 400830
rect 502190 400828 502196 400830
rect 502260 400828 502266 400892
rect 501822 400692 501828 400756
rect 501892 400754 501898 400756
rect 501965 400754 502031 400757
rect 501892 400752 502031 400754
rect 501892 400696 501970 400752
rect 502026 400696 502031 400752
rect 501892 400694 502031 400696
rect 501892 400692 501898 400694
rect 501965 400691 502031 400694
rect 82353 400210 82419 400213
rect 82486 400210 82492 400212
rect 82353 400208 82492 400210
rect 82353 400152 82358 400208
rect 82414 400152 82492 400208
rect 82353 400150 82492 400152
rect 82353 400147 82419 400150
rect 82486 400148 82492 400150
rect 82556 400148 82562 400212
rect 504030 398788 504036 398852
rect 504100 398788 504106 398852
rect 502057 398716 502123 398717
rect 502006 398714 502012 398716
rect 501966 398654 502012 398714
rect 502076 398712 502123 398716
rect 502118 398656 502123 398712
rect 502006 398652 502012 398654
rect 502076 398652 502123 398656
rect 504038 398714 504098 398788
rect 504398 398714 504404 398716
rect 504038 398654 504404 398714
rect 504398 398652 504404 398654
rect 504468 398652 504474 398716
rect 502057 398651 502123 398652
rect 502609 397898 502675 397901
rect 501860 397896 502675 397898
rect 501860 397840 502614 397896
rect 502670 397840 502675 397896
rect 501860 397838 502675 397840
rect 502609 397835 502675 397838
rect 82494 396813 82554 397324
rect 82445 396808 82554 396813
rect 82445 396752 82450 396808
rect 82506 396752 82554 396808
rect 82445 396750 82554 396752
rect 82445 396747 82511 396750
rect 82445 396132 82511 396133
rect 507025 396132 507091 396133
rect 82445 396128 82492 396132
rect 82556 396130 82562 396132
rect 506974 396130 506980 396132
rect 82445 396072 82450 396128
rect 82445 396068 82492 396072
rect 82556 396070 82602 396130
rect 506934 396070 506980 396130
rect 507044 396128 507091 396132
rect 507086 396072 507091 396128
rect 82556 396068 82562 396070
rect 506974 396068 506980 396070
rect 507044 396068 507091 396072
rect 82445 396067 82511 396068
rect 507025 396067 507091 396068
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 502241 394636 502307 394637
rect 507025 394636 507091 394637
rect 502190 394572 502196 394636
rect 502260 394634 502307 394636
rect 502260 394632 502352 394634
rect 502302 394576 502352 394632
rect 502260 394574 502352 394576
rect 502260 394572 502307 394574
rect 506974 394572 506980 394636
rect 507044 394634 507091 394636
rect 507044 394632 507136 394634
rect 507086 394576 507136 394632
rect 507044 394574 507136 394576
rect 507044 394572 507091 394574
rect 502241 394571 502307 394572
rect 507025 394571 507091 394572
rect 503294 394362 503300 394364
rect 501860 394302 503300 394362
rect 503294 394300 503300 394302
rect 503364 394300 503370 394364
rect 80830 394028 80836 394092
rect 80900 394090 80906 394092
rect 82302 394090 82308 394092
rect 80900 394030 82308 394090
rect 80900 394028 80906 394030
rect 82302 394028 82308 394030
rect 82372 394028 82378 394092
rect 78765 393818 78831 393821
rect 78765 393816 82156 393818
rect 78765 393760 78770 393816
rect 78826 393760 82156 393816
rect 78765 393758 82156 393760
rect 78765 393755 78831 393758
rect 80830 393076 80836 393140
rect 80900 393138 80906 393140
rect 82629 393138 82695 393141
rect 80900 393136 82695 393138
rect 80900 393080 82634 393136
rect 82690 393080 82695 393136
rect 80900 393078 82695 393080
rect 80900 393076 80906 393078
rect 82629 393075 82695 393078
rect 579705 393002 579771 393005
rect 583520 393002 584960 393092
rect 579705 393000 584960 393002
rect 579705 392944 579710 393000
rect 579766 392944 584960 393000
rect 579705 392942 584960 392944
rect 579705 392939 579771 392942
rect 583520 392852 584960 392942
rect 501638 391852 501644 391916
rect 501708 391852 501714 391916
rect 501646 391778 501706 391852
rect 501822 391778 501828 391780
rect 501646 391718 501828 391778
rect 501822 391716 501828 391718
rect 501892 391716 501898 391780
rect 82261 391234 82327 391237
rect 82486 391234 82492 391236
rect 82261 391232 82492 391234
rect 82261 391176 82266 391232
rect 82322 391176 82492 391232
rect 82261 391174 82492 391176
rect 82261 391171 82327 391174
rect 82486 391172 82492 391174
rect 82556 391172 82562 391236
rect 82077 391098 82143 391101
rect 82077 391096 82186 391098
rect 82077 391040 82082 391096
rect 82138 391040 82186 391096
rect 82077 391035 82186 391040
rect 82126 390524 82186 391035
rect 504541 390826 504607 390829
rect 501860 390824 504607 390826
rect 501860 390768 504546 390824
rect 504602 390768 504607 390824
rect 501860 390766 504607 390768
rect 504541 390763 504607 390766
rect 503294 388316 503300 388380
rect 503364 388378 503370 388380
rect 504173 388378 504239 388381
rect 503364 388376 504239 388378
rect 503364 388320 504178 388376
rect 504234 388320 504239 388376
rect 503364 388318 504239 388320
rect 503364 388316 503370 388318
rect 504173 388315 504239 388318
rect 504030 387290 504036 387292
rect 501860 387230 504036 387290
rect 504030 387228 504036 387230
rect 504100 387228 504106 387292
rect 502241 387156 502307 387157
rect 507025 387156 507091 387157
rect 502190 387154 502196 387156
rect 502150 387094 502196 387154
rect 502260 387152 502307 387156
rect 506974 387154 506980 387156
rect 502302 387096 502307 387152
rect 502190 387092 502196 387094
rect 502260 387092 502307 387096
rect 506934 387094 506980 387154
rect 507044 387152 507091 387156
rect 507086 387096 507091 387152
rect 506974 387092 506980 387094
rect 507044 387092 507091 387096
rect 502241 387091 502307 387092
rect 507025 387091 507091 387092
rect 80830 386956 80836 387020
rect 80900 387018 80906 387020
rect 80900 386958 82156 387018
rect 80900 386956 80906 386958
rect 82537 385796 82603 385797
rect 82486 385794 82492 385796
rect 82446 385734 82492 385794
rect 82556 385792 82603 385796
rect 82598 385736 82603 385792
rect 82486 385732 82492 385734
rect 82556 385732 82603 385736
rect 82537 385731 82603 385732
rect 80830 385596 80836 385660
rect 80900 385658 80906 385660
rect 82077 385658 82143 385661
rect 82353 385660 82419 385661
rect 82302 385658 82308 385660
rect 80900 385656 82143 385658
rect 80900 385600 82082 385656
rect 82138 385600 82143 385656
rect 80900 385598 82143 385600
rect 82262 385598 82308 385658
rect 82372 385656 82419 385660
rect 82414 385600 82419 385656
rect 80900 385596 80906 385598
rect 82077 385595 82143 385598
rect 82302 385596 82308 385598
rect 82372 385596 82419 385600
rect 82353 385595 82419 385596
rect 501454 385052 501460 385116
rect 501524 385114 501530 385116
rect 502006 385114 502012 385116
rect 501524 385054 502012 385114
rect 501524 385052 501530 385054
rect 502006 385052 502012 385054
rect 502076 385052 502082 385116
rect 502701 383754 502767 383757
rect 501860 383752 502767 383754
rect 501860 383696 502706 383752
rect 502762 383696 502767 383752
rect 501860 383694 502767 383696
rect 502701 383691 502767 383694
rect 78806 383420 78812 383484
rect 78876 383482 78882 383484
rect 78876 383422 82156 383482
rect 78876 383420 78882 383422
rect 503294 382468 503300 382532
rect 503364 382530 503370 382532
rect 507526 382530 507532 382532
rect 503364 382470 507532 382530
rect 503364 382468 503370 382470
rect 507526 382468 507532 382470
rect 507596 382468 507602 382532
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3049 380626 3115 380629
rect -960 380624 3115 380626
rect -960 380568 3054 380624
rect 3110 380568 3115 380624
rect -960 380566 3115 380568
rect -960 380476 480 380566
rect 3049 380563 3115 380566
rect 504265 380218 504331 380221
rect 501860 380216 504331 380218
rect 501860 380160 504270 380216
rect 504326 380160 504331 380216
rect 501860 380158 504331 380160
rect 504265 380155 504331 380158
rect 77569 379946 77635 379949
rect 77569 379944 82156 379946
rect 77569 379888 77574 379944
rect 77630 379888 82156 379944
rect 77569 379886 82156 379888
rect 77569 379883 77635 379886
rect 504173 376954 504239 376957
rect 501860 376952 504239 376954
rect 501860 376896 504178 376952
rect 504234 376896 504239 376952
rect 501860 376894 504239 376896
rect 504173 376891 504239 376894
rect 78622 376348 78628 376412
rect 78692 376410 78698 376412
rect 78692 376350 82156 376410
rect 78692 376348 78698 376350
rect 504173 373418 504239 373421
rect 501860 373416 504239 373418
rect 501860 373360 504178 373416
rect 504234 373360 504239 373416
rect 501860 373358 504239 373360
rect 504173 373355 504239 373358
rect 77569 372874 77635 372877
rect 77569 372872 82156 372874
rect 77569 372816 77574 372872
rect 77630 372816 82156 372872
rect 77569 372814 82156 372816
rect 77569 372811 77635 372814
rect 82445 371924 82511 371925
rect 82445 371922 82492 371924
rect 82400 371920 82492 371922
rect 82400 371864 82450 371920
rect 82400 371862 82492 371864
rect 82445 371860 82492 371862
rect 82556 371860 82562 371924
rect 82445 371859 82511 371860
rect 504541 369882 504607 369885
rect 501860 369880 504607 369882
rect 501860 369824 504546 369880
rect 504602 369824 504607 369880
rect 501860 369822 504607 369824
rect 504541 369819 504607 369822
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect 82494 369069 82554 369308
rect 82353 369068 82419 369069
rect 82302 369066 82308 369068
rect 82262 369006 82308 369066
rect 82372 369064 82419 369068
rect 82414 369008 82419 369064
rect 82302 369004 82308 369006
rect 82372 369004 82419 369008
rect 82494 369064 82603 369069
rect 82494 369008 82542 369064
rect 82598 369008 82603 369064
rect 82494 369006 82603 369008
rect 82353 369003 82419 369004
rect 82537 369003 82603 369006
rect 82302 368868 82308 368932
rect 82372 368930 82378 368932
rect 82629 368930 82695 368933
rect 82372 368928 82695 368930
rect 82372 368872 82634 368928
rect 82690 368872 82695 368928
rect 82372 368870 82695 368872
rect 82372 368868 82378 368870
rect 82629 368867 82695 368870
rect 82486 368732 82492 368796
rect 82556 368794 82562 368796
rect 82629 368794 82695 368797
rect 82556 368792 82695 368794
rect 82556 368736 82634 368792
rect 82690 368736 82695 368792
rect 82556 368734 82695 368736
rect 82556 368732 82562 368734
rect 82629 368731 82695 368734
rect 82445 368116 82511 368117
rect 82445 368112 82492 368116
rect 82556 368114 82562 368116
rect 82445 368056 82450 368112
rect 82445 368052 82492 368056
rect 82556 368054 82602 368114
rect 82556 368052 82562 368054
rect 82445 368051 82511 368052
rect 506013 366346 506079 366349
rect 501860 366344 506079 366346
rect -960 366210 480 366300
rect 501860 366288 506018 366344
rect 506074 366288 506079 366344
rect 501860 366286 506079 366288
rect 506013 366283 506079 366286
rect 3601 366210 3667 366213
rect -960 366208 3667 366210
rect -960 366152 3606 366208
rect 3662 366152 3667 366208
rect -960 366150 3667 366152
rect -960 366060 480 366150
rect 3601 366147 3667 366150
rect 82445 364852 82511 364853
rect 82445 364848 82492 364852
rect 82556 364850 82562 364852
rect 82445 364792 82450 364848
rect 82445 364788 82492 364792
rect 82556 364790 82602 364850
rect 82556 364788 82562 364790
rect 82445 364787 82511 364788
rect 82353 364714 82419 364717
rect 82486 364714 82492 364716
rect 82353 364712 82492 364714
rect 82353 364656 82358 364712
rect 82414 364656 82492 364712
rect 82353 364654 82492 364656
rect 82353 364651 82419 364654
rect 82486 364652 82492 364654
rect 82556 364652 82562 364716
rect 82353 362946 82419 362949
rect 82486 362946 82492 362948
rect 82353 362944 82492 362946
rect 82353 362888 82358 362944
rect 82414 362888 82492 362944
rect 82353 362886 82492 362888
rect 82353 362883 82419 362886
rect 82486 362884 82492 362886
rect 82556 362884 82562 362948
rect 82486 362748 82492 362812
rect 82556 362810 82562 362812
rect 82629 362810 82695 362813
rect 504541 362810 504607 362813
rect 82556 362808 82695 362810
rect 82556 362752 82634 362808
rect 82690 362752 82695 362808
rect 82556 362750 82695 362752
rect 501860 362808 504607 362810
rect 501860 362752 504546 362808
rect 504602 362752 504607 362808
rect 501860 362750 504607 362752
rect 82556 362748 82562 362750
rect 82629 362747 82695 362750
rect 504541 362747 504607 362750
rect 77569 362266 77635 362269
rect 77569 362264 82156 362266
rect 77569 362208 77574 362264
rect 77630 362208 82156 362264
rect 77569 362206 82156 362208
rect 77569 362203 77635 362206
rect 82353 360228 82419 360229
rect 82302 360226 82308 360228
rect 82262 360166 82308 360226
rect 82372 360224 82419 360228
rect 82414 360168 82419 360224
rect 82302 360164 82308 360166
rect 82372 360164 82419 360168
rect 82353 360163 82419 360164
rect 82629 360092 82695 360093
rect 82624 360090 82630 360092
rect 82538 360030 82630 360090
rect 82624 360028 82630 360030
rect 82694 360028 82700 360092
rect 82629 360027 82695 360028
rect 82445 359410 82511 359413
rect 82624 359410 82630 359412
rect 82445 359408 82630 359410
rect 82445 359352 82450 359408
rect 82506 359352 82630 359408
rect 82445 359350 82630 359352
rect 82445 359347 82511 359350
rect 82624 359348 82630 359350
rect 82694 359348 82700 359412
rect 502793 359274 502859 359277
rect 501860 359272 502859 359274
rect 501860 359216 502798 359272
rect 502854 359216 502859 359272
rect 501860 359214 502859 359216
rect 502793 359211 502859 359214
rect 74165 358730 74231 358733
rect 74165 358728 82156 358730
rect 74165 358672 74170 358728
rect 74226 358672 82156 358728
rect 74165 358670 82156 358672
rect 74165 358667 74231 358670
rect 501454 358532 501460 358596
rect 501524 358594 501530 358596
rect 502006 358594 502012 358596
rect 501524 358534 502012 358594
rect 501524 358532 501530 358534
rect 502006 358532 502012 358534
rect 502076 358532 502082 358596
rect 82629 358052 82695 358053
rect 82624 358050 82630 358052
rect 82538 357990 82630 358050
rect 82624 357988 82630 357990
rect 82694 357988 82700 358052
rect 82629 357987 82695 357988
rect 580625 357914 580691 357917
rect 583520 357914 584960 358004
rect 580625 357912 584960 357914
rect 580625 357856 580630 357912
rect 580686 357856 584960 357912
rect 580625 357854 584960 357856
rect 580625 357851 580691 357854
rect 583520 357764 584960 357854
rect 503110 355738 503116 355740
rect 501860 355678 503116 355738
rect 503110 355676 503116 355678
rect 503180 355676 503186 355740
rect 82126 354653 82186 355164
rect 82077 354648 82186 354653
rect 82077 354592 82082 354648
rect 82138 354592 82186 354648
rect 82077 354590 82186 354592
rect 82077 354587 82143 354590
rect 504173 352202 504239 352205
rect 501860 352200 504239 352202
rect 501860 352144 504178 352200
rect 504234 352144 504239 352200
rect 501860 352142 504239 352144
rect 504173 352139 504239 352142
rect -960 351780 480 352020
rect 79777 351658 79843 351661
rect 79777 351656 82156 351658
rect 79777 351600 79782 351656
rect 79838 351600 82156 351656
rect 79777 351598 82156 351600
rect 79777 351595 79843 351598
rect 501270 351596 501276 351660
rect 501340 351658 501346 351660
rect 501965 351658 502031 351661
rect 501340 351656 502031 351658
rect 501340 351600 501970 351656
rect 502026 351600 502031 351656
rect 501340 351598 502031 351600
rect 501340 351596 501346 351598
rect 501965 351595 502031 351598
rect 501454 350508 501460 350572
rect 501524 350570 501530 350572
rect 502057 350570 502123 350573
rect 501524 350568 502123 350570
rect 501524 350512 502062 350568
rect 502118 350512 502123 350568
rect 501524 350510 502123 350512
rect 501524 350508 501530 350510
rect 502057 350507 502123 350510
rect 501454 349828 501460 349892
rect 501524 349890 501530 349892
rect 504582 349890 504588 349892
rect 501524 349830 504588 349890
rect 501524 349828 501530 349830
rect 504582 349828 504588 349830
rect 504652 349828 504658 349892
rect 504030 349556 504036 349620
rect 504100 349618 504106 349620
rect 504582 349618 504588 349620
rect 504100 349558 504588 349618
rect 504100 349556 504106 349558
rect 504582 349556 504588 349558
rect 504652 349556 504658 349620
rect 504817 348666 504883 348669
rect 501860 348664 504883 348666
rect 501860 348608 504822 348664
rect 504878 348608 504883 348664
rect 501860 348606 504883 348608
rect 504817 348603 504883 348606
rect 79133 348122 79199 348125
rect 79133 348120 82156 348122
rect 79133 348064 79138 348120
rect 79194 348064 82156 348120
rect 79133 348062 82156 348064
rect 79133 348059 79199 348062
rect 504398 347652 504404 347716
rect 504468 347652 504474 347716
rect 504406 347578 504466 347652
rect 504541 347578 504607 347581
rect 504406 347576 504607 347578
rect 504406 347520 504546 347576
rect 504602 347520 504607 347576
rect 504406 347518 504607 347520
rect 504541 347515 504607 347518
rect 82537 347036 82603 347037
rect 82486 347034 82492 347036
rect 82446 346974 82492 347034
rect 82556 347032 82603 347036
rect 82598 346976 82603 347032
rect 82486 346972 82492 346974
rect 82556 346972 82603 346976
rect 82537 346971 82603 346972
rect 501454 346428 501460 346492
rect 501524 346490 501530 346492
rect 502057 346490 502123 346493
rect 501524 346488 502123 346490
rect 501524 346432 502062 346488
rect 502118 346432 502123 346488
rect 501524 346430 502123 346432
rect 501524 346428 501530 346430
rect 502057 346427 502123 346430
rect 501454 346292 501460 346356
rect 501524 346354 501530 346356
rect 501965 346354 502031 346357
rect 501524 346352 502031 346354
rect 501524 346296 501970 346352
rect 502026 346296 502031 346352
rect 501524 346294 502031 346296
rect 501524 346292 501530 346294
rect 501965 346291 502031 346294
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 504173 345130 504239 345133
rect 501860 345128 504239 345130
rect 501860 345072 504178 345128
rect 504234 345072 504239 345128
rect 501860 345070 504239 345072
rect 504173 345067 504239 345070
rect 506974 345068 506980 345132
rect 507044 345130 507050 345132
rect 507342 345130 507348 345132
rect 507044 345070 507348 345130
rect 507044 345068 507050 345070
rect 507342 345068 507348 345070
rect 507412 345068 507418 345132
rect 502149 344996 502215 344997
rect 502149 344994 502196 344996
rect 502104 344992 502196 344994
rect 502104 344936 502154 344992
rect 502104 344934 502196 344936
rect 502149 344932 502196 344934
rect 502260 344932 502266 344996
rect 502149 344931 502215 344932
rect 501270 344796 501276 344860
rect 501340 344796 501346 344860
rect 77569 344586 77635 344589
rect 77569 344584 82156 344586
rect 77569 344528 77574 344584
rect 77630 344528 82156 344584
rect 77569 344526 82156 344528
rect 77569 344523 77635 344526
rect 501278 344314 501338 344796
rect 501454 344314 501460 344316
rect 501278 344254 501460 344314
rect 501454 344252 501460 344254
rect 501524 344252 501530 344316
rect 82629 341732 82695 341733
rect 82624 341730 82630 341732
rect 82538 341670 82630 341730
rect 82624 341668 82630 341670
rect 82694 341668 82700 341732
rect 82629 341667 82695 341668
rect 503437 341594 503503 341597
rect 501860 341592 503503 341594
rect 501860 341536 503442 341592
rect 503498 341536 503503 341592
rect 501860 341534 503503 341536
rect 503437 341531 503503 341534
rect 73613 341050 73679 341053
rect 73613 341048 82156 341050
rect 73613 340992 73618 341048
rect 73674 340992 82156 341048
rect 73613 340990 82156 340992
rect 73613 340987 73679 340990
rect 82169 339690 82235 339693
rect 82486 339690 82492 339692
rect 82169 339688 82492 339690
rect 82169 339632 82174 339688
rect 82230 339632 82492 339688
rect 82169 339630 82492 339632
rect 82169 339627 82235 339630
rect 82486 339628 82492 339630
rect 82556 339628 82562 339692
rect 82353 339012 82419 339013
rect 82302 339010 82308 339012
rect 82262 338950 82308 339010
rect 82372 339008 82419 339012
rect 82414 338952 82419 339008
rect 82302 338948 82308 338950
rect 82372 338948 82419 338952
rect 501454 338948 501460 339012
rect 501524 339010 501530 339012
rect 502006 339010 502012 339012
rect 501524 338950 502012 339010
rect 501524 338948 501530 338950
rect 502006 338948 502012 338950
rect 502076 338948 502082 339012
rect 504030 338948 504036 339012
rect 504100 339010 504106 339012
rect 504582 339010 504588 339012
rect 504100 338950 504588 339010
rect 504100 338948 504106 338950
rect 504582 338948 504588 338950
rect 504652 338948 504658 339012
rect 82353 338947 82419 338948
rect 502006 338812 502012 338876
rect 502076 338874 502082 338876
rect 502149 338874 502215 338877
rect 504541 338876 504607 338877
rect 504541 338874 504588 338876
rect 502076 338872 502215 338874
rect 502076 338816 502154 338872
rect 502210 338816 502215 338872
rect 502076 338814 502215 338816
rect 504496 338872 504588 338874
rect 504496 338816 504546 338872
rect 504496 338814 504588 338816
rect 502076 338812 502082 338814
rect 502149 338811 502215 338814
rect 504541 338812 504588 338814
rect 504652 338812 504658 338876
rect 504541 338811 504607 338812
rect 80830 337996 80836 338060
rect 80900 338058 80906 338060
rect 82169 338058 82235 338061
rect 80900 338056 82235 338058
rect 80900 338000 82174 338056
rect 82230 338000 82235 338056
rect 80900 337998 82235 338000
rect 80900 337996 80906 337998
rect 82169 337995 82235 337998
rect -960 337514 480 337604
rect 2957 337514 3023 337517
rect -960 337512 3023 337514
rect -960 337456 2962 337512
rect 3018 337456 3023 337512
rect -960 337454 3023 337456
rect -960 337364 480 337454
rect 2957 337451 3023 337454
rect 79961 337514 80027 337517
rect 501830 337514 501890 338028
rect 502057 337514 502123 337517
rect 79961 337512 82156 337514
rect 79961 337456 79966 337512
rect 80022 337456 82156 337512
rect 79961 337454 82156 337456
rect 501830 337512 502123 337514
rect 501830 337456 502062 337512
rect 502118 337456 502123 337512
rect 501830 337454 502123 337456
rect 79961 337451 80027 337454
rect 502057 337451 502123 337454
rect 82537 336970 82603 336973
rect 82494 336968 82603 336970
rect 82494 336912 82542 336968
rect 82598 336912 82603 336968
rect 82494 336907 82603 336912
rect 82494 336836 82554 336907
rect 82486 336772 82492 336836
rect 82556 336772 82562 336836
rect 82537 335068 82603 335069
rect 82486 335066 82492 335068
rect 82446 335006 82492 335066
rect 82556 335064 82603 335068
rect 82598 335008 82603 335064
rect 82486 335004 82492 335006
rect 82556 335004 82603 335008
rect 82537 335003 82603 335004
rect 504541 334522 504607 334525
rect 501860 334520 504607 334522
rect 501860 334464 504546 334520
rect 504602 334464 504607 334520
rect 501860 334462 504607 334464
rect 504541 334459 504607 334462
rect 583520 334236 584960 334476
rect 76465 333978 76531 333981
rect 76465 333976 82156 333978
rect 76465 333920 76470 333976
rect 76526 333920 82156 333976
rect 76465 333918 82156 333920
rect 76465 333915 76531 333918
rect 82169 332210 82235 332213
rect 82486 332210 82492 332212
rect 82169 332208 82492 332210
rect 82169 332152 82174 332208
rect 82230 332152 82492 332208
rect 82169 332150 82492 332152
rect 82169 332147 82235 332150
rect 82486 332148 82492 332150
rect 82556 332148 82562 332212
rect 82353 331260 82419 331261
rect 82302 331258 82308 331260
rect 82262 331198 82308 331258
rect 82372 331256 82419 331260
rect 82414 331200 82419 331256
rect 82302 331196 82308 331198
rect 82372 331196 82419 331200
rect 82486 331196 82492 331260
rect 82556 331258 82562 331260
rect 82629 331258 82695 331261
rect 82556 331256 82695 331258
rect 82556 331200 82634 331256
rect 82690 331200 82695 331256
rect 82556 331198 82695 331200
rect 82556 331196 82562 331198
rect 82353 331195 82419 331196
rect 82629 331195 82695 331198
rect 82537 331124 82603 331125
rect 82486 331122 82492 331124
rect 82446 331062 82492 331122
rect 82556 331120 82603 331124
rect 82598 331064 82603 331120
rect 82486 331060 82492 331062
rect 82556 331060 82603 331064
rect 82537 331059 82603 331060
rect 504449 330986 504515 330989
rect 501860 330984 504515 330986
rect 501860 330928 504454 330984
rect 504510 330928 504515 330984
rect 501860 330926 504515 330928
rect 504449 330923 504515 330926
rect 77569 330442 77635 330445
rect 77569 330440 82156 330442
rect 77569 330384 77574 330440
rect 77630 330384 82156 330440
rect 77569 330382 82156 330384
rect 77569 330379 77635 330382
rect 506841 328404 506907 328405
rect 506790 328340 506796 328404
rect 506860 328402 506907 328404
rect 506860 328400 506952 328402
rect 506902 328344 506952 328400
rect 506860 328342 506952 328344
rect 506860 328340 506907 328342
rect 506841 328339 506907 328340
rect 80830 328068 80836 328132
rect 80900 328130 80906 328132
rect 82169 328130 82235 328133
rect 80900 328128 82235 328130
rect 80900 328072 82174 328128
rect 82230 328072 82235 328128
rect 80900 328070 82235 328072
rect 80900 328068 80906 328070
rect 82169 328067 82235 328070
rect 78254 327796 78260 327860
rect 78324 327858 78330 327860
rect 80830 327858 80836 327860
rect 78324 327798 80836 327858
rect 78324 327796 78330 327798
rect 80830 327796 80836 327798
rect 80900 327796 80906 327860
rect 81893 327450 81959 327453
rect 502885 327450 502951 327453
rect 81893 327448 82186 327450
rect 81893 327392 81898 327448
rect 81954 327392 82186 327448
rect 81893 327390 82186 327392
rect 501860 327448 502951 327450
rect 501860 327392 502890 327448
rect 502946 327392 502951 327448
rect 501860 327390 502951 327392
rect 81893 327387 81959 327390
rect 82126 326876 82186 327390
rect 502885 327387 502951 327390
rect 504582 326498 504588 326500
rect 503854 326438 504588 326498
rect 503854 326226 503914 326438
rect 504582 326436 504588 326438
rect 504652 326436 504658 326500
rect 504030 326300 504036 326364
rect 504100 326362 504106 326364
rect 504582 326362 504588 326364
rect 504100 326302 504588 326362
rect 504100 326300 504106 326302
rect 504582 326300 504588 326302
rect 504652 326300 504658 326364
rect 504030 326226 504036 326228
rect 503854 326166 504036 326226
rect 504030 326164 504036 326166
rect 504100 326164 504106 326228
rect 501638 325620 501644 325684
rect 501708 325682 501714 325684
rect 501965 325682 502031 325685
rect 501708 325680 502031 325682
rect 501708 325624 501970 325680
rect 502026 325624 502031 325680
rect 501708 325622 502031 325624
rect 501708 325620 501714 325622
rect 501965 325619 502031 325622
rect 504449 323914 504515 323917
rect 501860 323912 504515 323914
rect 501860 323856 504454 323912
rect 504510 323856 504515 323912
rect 501860 323854 504515 323856
rect 504449 323851 504515 323854
rect 77661 323642 77727 323645
rect 506841 323644 506907 323645
rect 506790 323642 506796 323644
rect 77661 323640 82156 323642
rect 77661 323584 77666 323640
rect 77722 323584 82156 323640
rect 77661 323582 82156 323584
rect 506750 323582 506796 323642
rect 506860 323640 506907 323644
rect 506902 323584 506907 323640
rect 77661 323579 77727 323582
rect 506790 323580 506796 323582
rect 506860 323580 506907 323584
rect 506841 323579 506907 323580
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 502149 320378 502215 320381
rect 501860 320376 502215 320378
rect 501860 320320 502154 320376
rect 502210 320320 502215 320376
rect 501860 320318 502215 320320
rect 502149 320315 502215 320318
rect 82678 319565 82738 320076
rect 82629 319560 82738 319565
rect 82629 319504 82634 319560
rect 82690 319504 82738 319560
rect 82629 319502 82738 319504
rect 82629 319499 82695 319502
rect 507526 319500 507532 319564
rect 507596 319562 507602 319564
rect 507669 319562 507735 319565
rect 507596 319560 507735 319562
rect 507596 319504 507674 319560
rect 507730 319504 507735 319560
rect 507596 319502 507735 319504
rect 507596 319500 507602 319502
rect 507669 319499 507735 319502
rect 507526 318820 507532 318884
rect 507596 318882 507602 318884
rect 507669 318882 507735 318885
rect 507596 318880 507735 318882
rect 507596 318824 507674 318880
rect 507730 318824 507735 318880
rect 507596 318822 507735 318824
rect 507596 318820 507602 318822
rect 507669 318819 507735 318822
rect 82445 317388 82511 317389
rect 82445 317386 82492 317388
rect 82400 317384 82492 317386
rect 82400 317328 82450 317384
rect 82400 317326 82492 317328
rect 82445 317324 82492 317326
rect 82556 317324 82562 317388
rect 82445 317323 82511 317324
rect 502517 316842 502583 316845
rect 501860 316840 502583 316842
rect 501860 316784 502522 316840
rect 502578 316784 502583 316840
rect 501860 316782 502583 316784
rect 502517 316779 502583 316782
rect 504582 316780 504588 316844
rect 504652 316842 504658 316844
rect 504652 316782 504834 316842
rect 504652 316780 504658 316782
rect 504030 316644 504036 316708
rect 504100 316706 504106 316708
rect 504582 316706 504588 316708
rect 504100 316646 504588 316706
rect 504100 316644 504106 316646
rect 504582 316644 504588 316646
rect 504652 316644 504658 316708
rect 80513 316570 80579 316573
rect 80513 316568 82156 316570
rect 80513 316512 80518 316568
rect 80574 316512 82156 316568
rect 80513 316510 82156 316512
rect 80513 316507 80579 316510
rect 504030 316508 504036 316572
rect 504100 316570 504106 316572
rect 504774 316570 504834 316782
rect 504100 316510 504834 316570
rect 504100 316508 504106 316510
rect 82445 316300 82511 316301
rect 82445 316296 82492 316300
rect 82556 316298 82562 316300
rect 82445 316240 82450 316296
rect 82445 316236 82492 316240
rect 82556 316238 82602 316298
rect 82556 316236 82562 316238
rect 82445 316235 82511 316236
rect 507342 315964 507348 316028
rect 507412 316026 507418 316028
rect 507669 316026 507735 316029
rect 507412 316024 507735 316026
rect 507412 315968 507674 316024
rect 507730 315968 507735 316024
rect 507412 315966 507735 315968
rect 507412 315964 507418 315966
rect 507669 315963 507735 315966
rect 501822 315828 501828 315892
rect 501892 315890 501898 315892
rect 501965 315890 502031 315893
rect 501892 315888 502031 315890
rect 501892 315832 501970 315888
rect 502026 315832 502031 315888
rect 501892 315830 502031 315832
rect 501892 315828 501898 315830
rect 501965 315827 502031 315830
rect 503294 313306 503300 313308
rect 501860 313246 503300 313306
rect 503294 313244 503300 313246
rect 503364 313244 503370 313308
rect 82678 312493 82738 313004
rect 82629 312488 82738 312493
rect 82629 312432 82634 312488
rect 82690 312432 82738 312488
rect 82629 312430 82738 312432
rect 82629 312427 82695 312430
rect 82445 312356 82511 312357
rect 82445 312354 82492 312356
rect 82400 312352 82492 312354
rect 82400 312296 82450 312352
rect 82400 312294 82492 312296
rect 82445 312292 82492 312294
rect 82556 312292 82562 312356
rect 82445 312291 82511 312292
rect 580533 310858 580599 310861
rect 583520 310858 584960 310948
rect 580533 310856 584960 310858
rect 580533 310800 580538 310856
rect 580594 310800 584960 310856
rect 580533 310798 584960 310800
rect 580533 310795 580599 310798
rect 583520 310708 584960 310798
rect 504449 310042 504515 310045
rect 501860 310040 504515 310042
rect 501860 309984 504454 310040
rect 504510 309984 504515 310040
rect 501860 309982 504515 309984
rect 504449 309979 504515 309982
rect 77569 309498 77635 309501
rect 77569 309496 82156 309498
rect 77569 309440 77574 309496
rect 77630 309440 82156 309496
rect 77569 309438 82156 309440
rect 77569 309435 77635 309438
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 501638 308484 501644 308548
rect 501708 308546 501714 308548
rect 501965 308546 502031 308549
rect 501708 308544 502031 308546
rect 501708 308488 501970 308544
rect 502026 308488 502031 308544
rect 501708 308486 502031 308488
rect 501708 308484 501714 308486
rect 501965 308483 502031 308486
rect 82445 307460 82511 307461
rect 82445 307458 82492 307460
rect 82400 307456 82492 307458
rect 82400 307400 82450 307456
rect 82400 307398 82492 307400
rect 82445 307396 82492 307398
rect 82556 307396 82562 307460
rect 82445 307395 82511 307396
rect 504582 307124 504588 307188
rect 504652 307186 504658 307188
rect 504725 307186 504791 307189
rect 504652 307184 504791 307186
rect 504652 307128 504730 307184
rect 504786 307128 504791 307184
rect 504652 307126 504791 307128
rect 504652 307124 504658 307126
rect 504725 307123 504791 307126
rect 504030 306988 504036 307052
rect 504100 307050 504106 307052
rect 504582 307050 504588 307052
rect 504100 306990 504588 307050
rect 504100 306988 504106 306990
rect 504582 306988 504588 306990
rect 504652 306988 504658 307052
rect 501454 306852 501460 306916
rect 501524 306914 501530 306916
rect 501638 306914 501644 306916
rect 501524 306854 501644 306914
rect 501524 306852 501530 306854
rect 501638 306852 501644 306854
rect 501708 306852 501714 306916
rect 504449 306506 504515 306509
rect 501860 306504 504515 306506
rect 501860 306448 504454 306504
rect 504510 306448 504515 306504
rect 501860 306446 504515 306448
rect 504449 306443 504515 306446
rect 82678 305421 82738 305932
rect 82629 305416 82738 305421
rect 82629 305360 82634 305416
rect 82690 305360 82738 305416
rect 82629 305358 82738 305360
rect 82629 305355 82695 305358
rect 502517 302970 502583 302973
rect 501860 302968 502583 302970
rect 501860 302912 502522 302968
rect 502578 302912 502583 302968
rect 501860 302910 502583 302912
rect 502517 302907 502583 302910
rect 82126 301885 82186 302396
rect 82126 301880 82235 301885
rect 82126 301824 82174 301880
rect 82230 301824 82235 301880
rect 82126 301822 82235 301824
rect 82169 301819 82235 301822
rect 503161 299434 503227 299437
rect 501860 299432 503227 299434
rect 501860 299376 503166 299432
rect 503222 299376 503227 299432
rect 501860 299374 503227 299376
rect 503161 299371 503227 299374
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 81014 298828 81020 298892
rect 81084 298890 81090 298892
rect 81084 298830 82156 298890
rect 81084 298828 81090 298830
rect 82537 297804 82603 297805
rect 82486 297740 82492 297804
rect 82556 297802 82603 297804
rect 82556 297800 82648 297802
rect 82598 297744 82648 297800
rect 82556 297742 82648 297744
rect 82556 297740 82603 297742
rect 82537 297739 82603 297740
rect 82486 297468 82492 297532
rect 82556 297530 82562 297532
rect 82629 297530 82695 297533
rect 82556 297528 82695 297530
rect 82556 297472 82634 297528
rect 82690 297472 82695 297528
rect 82556 297470 82695 297472
rect 82556 297468 82562 297470
rect 82629 297467 82695 297470
rect 504030 297468 504036 297532
rect 504100 297530 504106 297532
rect 504582 297530 504588 297532
rect 504100 297470 504588 297530
rect 504100 297468 504106 297470
rect 504582 297468 504588 297470
rect 504652 297468 504658 297532
rect 504398 297332 504404 297396
rect 504468 297394 504474 297396
rect 504725 297394 504791 297397
rect 507025 297396 507091 297397
rect 506974 297394 506980 297396
rect 504468 297392 504791 297394
rect 504468 297336 504730 297392
rect 504786 297336 504791 297392
rect 504468 297334 504791 297336
rect 506934 297334 506980 297394
rect 507044 297392 507091 297396
rect 507086 297336 507091 297392
rect 504468 297332 504474 297334
rect 504725 297331 504791 297334
rect 506974 297332 506980 297334
rect 507044 297332 507091 297336
rect 507025 297331 507091 297332
rect 82353 296850 82419 296853
rect 82486 296850 82492 296852
rect 82353 296848 82492 296850
rect 82353 296792 82358 296848
rect 82414 296792 82492 296848
rect 82353 296790 82492 296792
rect 82353 296787 82419 296790
rect 82486 296788 82492 296790
rect 82556 296788 82562 296852
rect 504449 295898 504515 295901
rect 501860 295896 504515 295898
rect 501860 295840 504454 295896
rect 504510 295840 504515 295896
rect 501860 295838 504515 295840
rect 504449 295835 504515 295838
rect 77569 295490 77635 295493
rect 78254 295490 78260 295492
rect 77569 295488 78260 295490
rect 77569 295432 77574 295488
rect 77630 295432 78260 295488
rect 77569 295430 78260 295432
rect 77569 295427 77635 295430
rect 78254 295428 78260 295430
rect 78324 295428 78330 295492
rect 82310 294813 82370 295324
rect 82261 294808 82370 294813
rect 82261 294752 82266 294808
rect 82322 294752 82370 294808
rect 82261 294750 82370 294752
rect 82261 294747 82327 294750
rect -960 294402 480 294492
rect 3233 294402 3299 294405
rect -960 294400 3299 294402
rect -960 294344 3238 294400
rect 3294 294344 3299 294400
rect -960 294342 3299 294344
rect -960 294252 480 294342
rect 3233 294339 3299 294342
rect 80830 293388 80836 293452
rect 80900 293450 80906 293452
rect 82486 293450 82492 293452
rect 80900 293390 82492 293450
rect 80900 293388 80906 293390
rect 82486 293388 82492 293390
rect 82556 293388 82562 293452
rect 505001 292362 505067 292365
rect 501860 292360 505067 292362
rect 501860 292304 505006 292360
rect 505062 292304 505067 292360
rect 501860 292302 505067 292304
rect 505001 292299 505067 292302
rect 82486 292028 82492 292092
rect 82556 292090 82562 292092
rect 82629 292090 82695 292093
rect 82556 292088 82695 292090
rect 82556 292032 82634 292088
rect 82690 292032 82695 292088
rect 82556 292030 82695 292032
rect 82556 292028 82562 292030
rect 82629 292027 82695 292030
rect 81893 291274 81959 291277
rect 82126 291274 82186 291788
rect 82353 291274 82419 291277
rect 81893 291272 82186 291274
rect 81893 291216 81898 291272
rect 81954 291216 82186 291272
rect 81893 291214 82186 291216
rect 82310 291272 82419 291274
rect 82310 291216 82358 291272
rect 82414 291216 82419 291272
rect 81893 291211 81959 291214
rect 82310 291211 82419 291216
rect 82310 291140 82370 291211
rect 82302 291076 82308 291140
rect 82372 291076 82378 291140
rect 501965 290460 502031 290461
rect 501965 290458 502012 290460
rect 501920 290456 502012 290458
rect 501920 290400 501970 290456
rect 501920 290398 502012 290400
rect 501965 290396 502012 290398
rect 502076 290396 502082 290460
rect 506974 290396 506980 290460
rect 507044 290458 507050 290460
rect 507342 290458 507348 290460
rect 507044 290398 507348 290458
rect 507044 290396 507050 290398
rect 507342 290396 507348 290398
rect 507412 290396 507418 290460
rect 501965 290395 502031 290396
rect 501454 290260 501460 290324
rect 501524 290322 501530 290324
rect 501965 290322 502031 290325
rect 501524 290320 502031 290322
rect 501524 290264 501970 290320
rect 502026 290264 502031 290320
rect 501524 290262 502031 290264
rect 501524 290260 501530 290262
rect 501965 290259 502031 290262
rect 501965 290186 502031 290189
rect 504214 290186 504220 290188
rect 501965 290184 504220 290186
rect 501965 290128 501970 290184
rect 502026 290128 504220 290184
rect 501965 290126 504220 290128
rect 501965 290123 502031 290126
rect 504214 290124 504220 290126
rect 504284 290124 504290 290188
rect 501454 289988 501460 290052
rect 501524 290050 501530 290052
rect 502241 290050 502307 290053
rect 501524 290048 502307 290050
rect 501524 289992 502246 290048
rect 502302 289992 502307 290048
rect 501524 289990 502307 289992
rect 501524 289988 501530 289990
rect 502241 289987 502307 289990
rect 82537 289100 82603 289101
rect 82486 289098 82492 289100
rect 82446 289038 82492 289098
rect 82556 289096 82603 289100
rect 82598 289040 82603 289096
rect 82486 289036 82492 289038
rect 82556 289036 82603 289040
rect 501270 289036 501276 289100
rect 501340 289098 501346 289100
rect 501638 289098 501644 289100
rect 501340 289038 501644 289098
rect 501340 289036 501346 289038
rect 501638 289036 501644 289038
rect 501708 289036 501714 289100
rect 82537 289035 82603 289036
rect 504449 288826 504515 288829
rect 501860 288824 504515 288826
rect 501860 288768 504454 288824
rect 504510 288768 504515 288824
rect 501860 288766 504515 288768
rect 504449 288763 504515 288766
rect 76649 288282 76715 288285
rect 76649 288280 82156 288282
rect 76649 288224 76654 288280
rect 76710 288224 82156 288280
rect 76649 288222 82156 288224
rect 76649 288219 76715 288222
rect 583520 287316 584960 287556
rect 504030 286996 504036 287060
rect 504100 287058 504106 287060
rect 504214 287058 504220 287060
rect 504100 286998 504220 287058
rect 504100 286996 504106 286998
rect 504214 286996 504220 286998
rect 504284 286996 504290 287060
rect 501454 286316 501460 286380
rect 501524 286378 501530 286380
rect 501822 286378 501828 286380
rect 501524 286318 501828 286378
rect 501524 286316 501530 286318
rect 501822 286316 501828 286318
rect 501892 286316 501898 286380
rect 79501 284746 79567 284749
rect 501278 284748 501338 285260
rect 79501 284744 82156 284746
rect 79501 284688 79506 284744
rect 79562 284688 82156 284744
rect 79501 284686 82156 284688
rect 79501 284683 79567 284686
rect 501270 284684 501276 284748
rect 501340 284684 501346 284748
rect 501454 282372 501460 282436
rect 501524 282434 501530 282436
rect 501965 282434 502031 282437
rect 501524 282432 502031 282434
rect 501524 282376 501970 282432
rect 502026 282376 502031 282432
rect 501524 282374 502031 282376
rect 501524 282372 501530 282374
rect 501965 282371 502031 282374
rect 501965 282300 502031 282301
rect 501965 282298 502012 282300
rect 501920 282296 502012 282298
rect 501920 282240 501970 282296
rect 501920 282238 502012 282240
rect 501965 282236 502012 282238
rect 502076 282236 502082 282300
rect 501965 282235 502031 282236
rect 504725 281754 504791 281757
rect 501860 281752 504791 281754
rect 501860 281696 504730 281752
rect 504786 281696 504791 281752
rect 501860 281694 504791 281696
rect 504725 281691 504791 281694
rect 501270 281420 501276 281484
rect 501340 281482 501346 281484
rect 501965 281482 502031 281485
rect 501340 281480 502031 281482
rect 501340 281424 501970 281480
rect 502026 281424 502031 281480
rect 501340 281422 502031 281424
rect 501340 281420 501346 281422
rect 501965 281419 502031 281422
rect 75637 281210 75703 281213
rect 75637 281208 82156 281210
rect 75637 281152 75642 281208
rect 75698 281152 82156 281208
rect 75637 281150 82156 281152
rect 75637 281147 75703 281150
rect 78254 280876 78260 280940
rect 78324 280938 78330 280940
rect 82302 280938 82308 280940
rect 78324 280878 82308 280938
rect 78324 280876 78330 280878
rect 82302 280876 82308 280878
rect 82372 280876 82378 280940
rect 507025 280802 507091 280805
rect 507342 280802 507348 280804
rect 507025 280800 507348 280802
rect 507025 280744 507030 280800
rect 507086 280744 507348 280800
rect 507025 280742 507348 280744
rect 507025 280739 507091 280742
rect 507342 280740 507348 280742
rect 507412 280740 507418 280804
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 524413 278762 524479 278765
rect 524597 278762 524663 278765
rect 524413 278760 524663 278762
rect 524413 278704 524418 278760
rect 524474 278704 524602 278760
rect 524658 278704 524663 278760
rect 524413 278702 524663 278704
rect 524413 278699 524479 278702
rect 524597 278699 524663 278702
rect 502241 278218 502307 278221
rect 501860 278216 502307 278218
rect 501860 278160 502246 278216
rect 502302 278160 502307 278216
rect 501860 278158 502307 278160
rect 502241 278155 502307 278158
rect 75453 277674 75519 277677
rect 75453 277672 82156 277674
rect 75453 277616 75458 277672
rect 75514 277616 82156 277672
rect 75453 277614 82156 277616
rect 75453 277611 75519 277614
rect 501638 276524 501644 276588
rect 501708 276524 501714 276588
rect 501454 276252 501460 276316
rect 501524 276314 501530 276316
rect 501646 276314 501706 276524
rect 501524 276254 501706 276314
rect 501524 276252 501530 276254
rect 501822 275844 501828 275908
rect 501892 275906 501898 275908
rect 501892 275846 502258 275906
rect 501892 275844 501898 275846
rect 501454 275226 501460 275228
rect 501278 275166 501460 275226
rect 501278 274954 501338 275166
rect 501454 275164 501460 275166
rect 501524 275164 501530 275228
rect 501454 275028 501460 275092
rect 501524 275090 501530 275092
rect 501965 275090 502031 275093
rect 501524 275088 502031 275090
rect 501524 275032 501970 275088
rect 502026 275032 502031 275088
rect 501524 275030 502031 275032
rect 501524 275028 501530 275030
rect 501965 275027 502031 275030
rect 501454 274954 501460 274956
rect 501278 274894 501460 274954
rect 501454 274892 501460 274894
rect 501524 274892 501530 274956
rect 502006 274892 502012 274956
rect 502076 274954 502082 274956
rect 502198 274954 502258 275846
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 502076 274894 502258 274954
rect 502076 274892 502082 274894
rect 504173 274682 504239 274685
rect 501860 274680 504239 274682
rect 501860 274624 504178 274680
rect 504234 274624 504239 274680
rect 501860 274622 504239 274624
rect 504173 274619 504239 274622
rect 79317 274138 79383 274141
rect 79317 274136 82156 274138
rect 79317 274080 79322 274136
rect 79378 274080 82156 274136
rect 79317 274078 82156 274080
rect 79317 274075 79383 274078
rect 501270 274076 501276 274140
rect 501340 274138 501346 274140
rect 502190 274138 502196 274140
rect 501340 274078 502196 274138
rect 501340 274076 501346 274078
rect 502190 274076 502196 274078
rect 502260 274076 502266 274140
rect 78254 274002 78260 274004
rect 78078 273942 78260 274002
rect 78078 273458 78138 273942
rect 78254 273940 78260 273942
rect 78324 273940 78330 274004
rect 78254 273458 78260 273460
rect 78078 273398 78260 273458
rect 78254 273396 78260 273398
rect 78324 273396 78330 273460
rect 501638 273322 501644 273324
rect 501278 273262 501644 273322
rect 501278 272914 501338 273262
rect 501638 273260 501644 273262
rect 501708 273260 501714 273324
rect 501454 273124 501460 273188
rect 501524 273186 501530 273188
rect 501965 273186 502031 273189
rect 501524 273184 502031 273186
rect 501524 273128 501970 273184
rect 502026 273128 502031 273184
rect 501524 273126 502031 273128
rect 501524 273124 501530 273126
rect 501965 273123 502031 273126
rect 501454 272914 501460 272916
rect 501278 272854 501460 272914
rect 501454 272852 501460 272854
rect 501524 272852 501530 272916
rect 501638 272580 501644 272644
rect 501708 272642 501714 272644
rect 501965 272642 502031 272645
rect 501708 272640 502031 272642
rect 501708 272584 501970 272640
rect 502026 272584 502031 272640
rect 501708 272582 502031 272584
rect 501708 272580 501714 272582
rect 501965 272579 502031 272582
rect 501454 272444 501460 272508
rect 501524 272506 501530 272508
rect 501965 272506 502031 272509
rect 501524 272504 502031 272506
rect 501524 272448 501970 272504
rect 502026 272448 502031 272504
rect 501524 272446 502031 272448
rect 501524 272444 501530 272446
rect 501965 272443 502031 272446
rect 501270 272308 501276 272372
rect 501340 272370 501346 272372
rect 501965 272370 502031 272373
rect 501340 272368 502031 272370
rect 501340 272312 501970 272368
rect 502026 272312 502031 272368
rect 501340 272310 502031 272312
rect 501340 272308 501346 272310
rect 501965 272307 502031 272310
rect 504582 271764 504588 271828
rect 504652 271826 504658 271828
rect 504725 271826 504791 271829
rect 504652 271824 504791 271826
rect 504652 271768 504730 271824
rect 504786 271768 504791 271824
rect 504652 271766 504791 271768
rect 504652 271764 504658 271766
rect 504725 271763 504791 271766
rect 503253 271146 503319 271149
rect 501860 271144 503319 271146
rect 501860 271088 503258 271144
rect 503314 271088 503319 271144
rect 501860 271086 503319 271088
rect 503253 271083 503319 271086
rect 501270 270812 501276 270876
rect 501340 270874 501346 270876
rect 501965 270874 502031 270877
rect 501340 270872 502031 270874
rect 501340 270816 501970 270872
rect 502026 270816 502031 270872
rect 501340 270814 502031 270816
rect 501340 270812 501346 270814
rect 501965 270811 502031 270814
rect 507025 270738 507091 270741
rect 506982 270736 507091 270738
rect 506982 270680 507030 270736
rect 507086 270680 507091 270736
rect 506982 270675 507091 270680
rect 80830 270540 80836 270604
rect 80900 270602 80906 270604
rect 80900 270542 82156 270602
rect 80900 270540 80906 270542
rect 502006 270540 502012 270604
rect 502076 270602 502082 270604
rect 503437 270602 503503 270605
rect 506982 270604 507042 270675
rect 502076 270600 503503 270602
rect 502076 270544 503442 270600
rect 503498 270544 503503 270600
rect 502076 270542 503503 270544
rect 502076 270540 502082 270542
rect 503437 270539 503503 270542
rect 506974 270540 506980 270604
rect 507044 270540 507050 270604
rect 501270 270404 501276 270468
rect 501340 270466 501346 270468
rect 501965 270466 502031 270469
rect 501340 270464 502031 270466
rect 501340 270408 501970 270464
rect 502026 270408 502031 270464
rect 501340 270406 502031 270408
rect 501340 270404 501346 270406
rect 501965 270403 502031 270406
rect 503345 270330 503411 270333
rect 504582 270330 504588 270332
rect 503345 270328 504588 270330
rect 503345 270272 503350 270328
rect 503406 270272 504588 270328
rect 503345 270270 504588 270272
rect 503345 270267 503411 270270
rect 504582 270268 504588 270270
rect 504652 270268 504658 270332
rect 78254 269588 78260 269652
rect 78324 269650 78330 269652
rect 82629 269650 82695 269653
rect 78324 269648 82695 269650
rect 78324 269592 82634 269648
rect 82690 269592 82695 269648
rect 78324 269590 82695 269592
rect 78324 269588 78330 269590
rect 82629 269587 82695 269590
rect 501270 268228 501276 268292
rect 501340 268290 501346 268292
rect 501965 268290 502031 268293
rect 501340 268288 502031 268290
rect 501340 268232 501970 268288
rect 502026 268232 502031 268288
rect 501340 268230 502031 268232
rect 501340 268228 501346 268230
rect 501965 268227 502031 268230
rect 501830 267202 501890 267580
rect 502006 267202 502012 267204
rect 501830 267142 502012 267202
rect 502006 267140 502012 267142
rect 502076 267140 502082 267204
rect 77569 267066 77635 267069
rect 77569 267064 82156 267066
rect 77569 267008 77574 267064
rect 77630 267008 82156 267064
rect 77569 267006 82156 267008
rect 77569 267003 77635 267006
rect 501270 267004 501276 267068
rect 501340 267066 501346 267068
rect 501965 267066 502031 267069
rect 501340 267064 502031 267066
rect 501340 267008 501970 267064
rect 502026 267008 502031 267064
rect 501340 267006 502031 267008
rect 501340 267004 501346 267006
rect 501965 267003 502031 267006
rect 504582 267004 504588 267068
rect 504652 267066 504658 267068
rect 504725 267066 504791 267069
rect 504652 267064 504791 267066
rect 504652 267008 504730 267064
rect 504786 267008 504791 267064
rect 504652 267006 504791 267008
rect 504652 267004 504658 267006
rect 504725 267003 504791 267006
rect 82445 266250 82511 266253
rect 82624 266250 82630 266252
rect 82445 266248 82630 266250
rect 82445 266192 82450 266248
rect 82506 266192 82630 266248
rect 82445 266190 82630 266192
rect 82445 266187 82511 266190
rect 82624 266188 82630 266190
rect 82694 266188 82700 266252
rect -960 265706 480 265796
rect 2957 265706 3023 265709
rect -960 265704 3023 265706
rect -960 265648 2962 265704
rect 3018 265648 3023 265704
rect -960 265646 3023 265648
rect -960 265556 480 265646
rect 2957 265643 3023 265646
rect 82629 264074 82695 264077
rect 82629 264072 82738 264074
rect 82629 264016 82634 264072
rect 82690 264016 82738 264072
rect 82629 264011 82738 264016
rect 82678 263500 82738 264011
rect 501270 263468 501276 263532
rect 501340 263468 501346 263532
rect 501830 263530 501890 264044
rect 583520 263938 584960 264028
rect 518942 263878 528570 263938
rect 507526 263604 507532 263668
rect 507596 263666 507602 263668
rect 518942 263666 519002 263878
rect 528510 263802 528570 263878
rect 538262 263878 547890 263938
rect 528510 263742 538138 263802
rect 507596 263606 519002 263666
rect 538078 263666 538138 263742
rect 538262 263666 538322 263878
rect 547830 263802 547890 263878
rect 557582 263878 567210 263938
rect 547830 263742 557458 263802
rect 538078 263606 538322 263666
rect 557398 263666 557458 263742
rect 557582 263666 557642 263878
rect 567150 263802 567210 263878
rect 583342 263878 584960 263938
rect 583342 263802 583402 263878
rect 567150 263742 576778 263802
rect 557398 263606 557642 263666
rect 576718 263666 576778 263742
rect 576902 263742 583402 263802
rect 583520 263788 584960 263878
rect 576902 263666 576962 263742
rect 576718 263606 576962 263666
rect 507596 263604 507602 263606
rect 501965 263530 502031 263533
rect 501830 263528 502031 263530
rect 501830 263472 501970 263528
rect 502026 263472 502031 263528
rect 501830 263470 502031 263472
rect 501278 263394 501338 263468
rect 501965 263467 502031 263470
rect 502006 263394 502012 263396
rect 501278 263334 502012 263394
rect 502006 263332 502012 263334
rect 502076 263332 502082 263396
rect 77886 262788 77892 262852
rect 77956 262850 77962 262852
rect 82624 262850 82630 262852
rect 77956 262790 82630 262850
rect 77956 262788 77962 262790
rect 82624 262788 82630 262790
rect 82694 262788 82700 262852
rect 501638 262380 501644 262444
rect 501708 262442 501714 262444
rect 503529 262442 503595 262445
rect 501708 262440 503595 262442
rect 501708 262384 503534 262440
rect 503590 262384 503595 262440
rect 501708 262382 503595 262384
rect 501708 262380 501714 262382
rect 503529 262379 503595 262382
rect 506974 261428 506980 261492
rect 507044 261490 507050 261492
rect 507342 261490 507348 261492
rect 507044 261430 507348 261490
rect 507044 261428 507050 261430
rect 507342 261428 507348 261430
rect 507412 261428 507418 261492
rect 78254 260748 78260 260812
rect 78324 260810 78330 260812
rect 82624 260810 82630 260812
rect 78324 260750 82630 260810
rect 78324 260748 78330 260750
rect 82624 260748 82630 260750
rect 82694 260748 82700 260812
rect 504909 260538 504975 260541
rect 501860 260536 504975 260538
rect 501860 260480 504914 260536
rect 504970 260480 504975 260536
rect 501860 260478 504975 260480
rect 504909 260475 504975 260478
rect 82445 260266 82511 260269
rect 82624 260266 82630 260268
rect 82445 260264 82630 260266
rect 82445 260208 82450 260264
rect 82506 260208 82630 260264
rect 82445 260206 82630 260208
rect 82445 260203 82511 260206
rect 82624 260204 82630 260206
rect 82694 260204 82700 260268
rect 501270 260204 501276 260268
rect 501340 260266 501346 260268
rect 503621 260266 503687 260269
rect 501340 260264 503687 260266
rect 501340 260208 503626 260264
rect 503682 260208 503687 260264
rect 501340 260206 503687 260208
rect 501340 260204 501346 260206
rect 503621 260203 503687 260206
rect 503437 260130 503503 260133
rect 501830 260128 503503 260130
rect 501830 260072 503442 260128
rect 503498 260072 503503 260128
rect 501830 260070 503503 260072
rect 79225 259994 79291 259997
rect 79225 259992 82156 259994
rect 79225 259936 79230 259992
rect 79286 259936 82156 259992
rect 79225 259934 82156 259936
rect 79225 259931 79291 259934
rect 501830 259860 501890 260070
rect 503437 260067 503503 260070
rect 501822 259796 501828 259860
rect 501892 259796 501898 259860
rect 503529 259586 503595 259589
rect 502198 259584 503595 259586
rect 502198 259528 503534 259584
rect 503590 259528 503595 259584
rect 502198 259526 503595 259528
rect 502198 259450 502258 259526
rect 503529 259523 503595 259526
rect 503345 259450 503411 259453
rect 502198 259448 503411 259450
rect 502198 259392 503350 259448
rect 503406 259392 503411 259448
rect 502198 259390 503411 259392
rect 503345 259387 503411 259390
rect 524413 259450 524479 259453
rect 524597 259450 524663 259453
rect 524413 259448 524663 259450
rect 524413 259392 524418 259448
rect 524474 259392 524602 259448
rect 524658 259392 524663 259448
rect 524413 259390 524663 259392
rect 524413 259387 524479 259390
rect 524597 259387 524663 259390
rect 501270 258708 501276 258772
rect 501340 258770 501346 258772
rect 503529 258770 503595 258773
rect 501340 258768 503595 258770
rect 501340 258712 503534 258768
rect 503590 258712 503595 258768
rect 501340 258710 503595 258712
rect 501340 258708 501346 258710
rect 503529 258707 503595 258710
rect 504725 257002 504791 257005
rect 501860 257000 504791 257002
rect 501860 256944 504730 257000
rect 504786 256944 504791 257000
rect 501860 256942 504791 256944
rect 504725 256939 504791 256942
rect 77477 256730 77543 256733
rect 77477 256728 82156 256730
rect 77477 256672 77482 256728
rect 77538 256672 82156 256728
rect 77477 256670 82156 256672
rect 77477 256667 77543 256670
rect 501270 256668 501276 256732
rect 501340 256730 501346 256732
rect 503437 256730 503503 256733
rect 501340 256728 503503 256730
rect 501340 256672 503442 256728
rect 503498 256672 503503 256728
rect 501340 256670 503503 256672
rect 501340 256668 501346 256670
rect 503437 256667 503503 256670
rect 501454 256260 501460 256324
rect 501524 256322 501530 256324
rect 501822 256322 501828 256324
rect 501524 256262 501828 256322
rect 501524 256260 501530 256262
rect 501822 256260 501828 256262
rect 501892 256260 501898 256324
rect 501454 256124 501460 256188
rect 501524 256186 501530 256188
rect 503529 256186 503595 256189
rect 501524 256184 503595 256186
rect 501524 256128 503534 256184
rect 503590 256128 503595 256184
rect 501524 256126 503595 256128
rect 501524 256124 501530 256126
rect 503529 256123 503595 256126
rect 502190 255642 502196 255644
rect 501462 255582 502196 255642
rect 77702 255444 77708 255508
rect 77772 255506 77778 255508
rect 77886 255506 77892 255508
rect 77772 255446 77892 255506
rect 77772 255444 77778 255446
rect 77886 255444 77892 255446
rect 77956 255444 77962 255508
rect 501462 254962 501522 255582
rect 502190 255580 502196 255582
rect 502260 255580 502266 255644
rect 501638 255444 501644 255508
rect 501708 255506 501714 255508
rect 502190 255506 502196 255508
rect 501708 255446 502196 255506
rect 501708 255444 501714 255446
rect 502190 255444 502196 255446
rect 502260 255444 502266 255508
rect 501638 255308 501644 255372
rect 501708 255370 501714 255372
rect 503345 255370 503411 255373
rect 501708 255368 503411 255370
rect 501708 255312 503350 255368
rect 503406 255312 503411 255368
rect 501708 255310 503411 255312
rect 501708 255308 501714 255310
rect 503345 255307 503411 255310
rect 501822 255036 501828 255100
rect 501892 255098 501898 255100
rect 503621 255098 503687 255101
rect 501892 255096 503687 255098
rect 501892 255040 503626 255096
rect 503682 255040 503687 255096
rect 501892 255038 503687 255040
rect 501892 255036 501898 255038
rect 503621 255035 503687 255038
rect 503529 254962 503595 254965
rect 501462 254960 503595 254962
rect 501462 254904 503534 254960
rect 503590 254904 503595 254960
rect 501462 254902 503595 254904
rect 503529 254899 503595 254902
rect 82537 254828 82603 254829
rect 82486 254764 82492 254828
rect 82556 254826 82603 254828
rect 82556 254824 82648 254826
rect 82598 254768 82648 254824
rect 82556 254766 82648 254768
rect 82556 254764 82603 254766
rect 82537 254763 82603 254764
rect 501822 254492 501828 254556
rect 501892 254554 501898 254556
rect 503345 254554 503411 254557
rect 501892 254552 503411 254554
rect 501892 254496 503350 254552
rect 503406 254496 503411 254552
rect 501892 254494 503411 254496
rect 501892 254492 501898 254494
rect 503345 254491 503411 254494
rect 501638 254084 501644 254148
rect 501708 254146 501714 254148
rect 503345 254146 503411 254149
rect 501708 254144 503411 254146
rect 501708 254088 503350 254144
rect 503406 254088 503411 254144
rect 501708 254086 503411 254088
rect 501708 254084 501714 254086
rect 503345 254083 503411 254086
rect 77886 253948 77892 254012
rect 77956 254010 77962 254012
rect 82486 254010 82492 254012
rect 77956 253950 82492 254010
rect 77956 253948 77962 253950
rect 82486 253948 82492 253950
rect 82556 253948 82562 254012
rect 505829 253466 505895 253469
rect 501860 253464 505895 253466
rect 501860 253408 505834 253464
rect 505890 253408 505895 253464
rect 501860 253406 505895 253408
rect 505829 253403 505895 253406
rect 79041 253194 79107 253197
rect 79041 253192 82156 253194
rect 79041 253136 79046 253192
rect 79102 253136 82156 253192
rect 79041 253134 82156 253136
rect 79041 253131 79107 253134
rect 501270 253132 501276 253196
rect 501340 253132 501346 253196
rect 501454 253132 501460 253196
rect 501524 253194 501530 253196
rect 503437 253194 503503 253197
rect 501524 253192 503503 253194
rect 501524 253136 503442 253192
rect 503498 253136 503503 253192
rect 501524 253134 503503 253136
rect 501524 253132 501530 253134
rect 501278 253058 501338 253132
rect 503437 253131 503503 253134
rect 503437 253058 503503 253061
rect 501278 253056 503503 253058
rect 501278 253000 503442 253056
rect 503498 253000 503503 253056
rect 501278 252998 503503 253000
rect 503437 252995 503503 252998
rect 82537 252788 82603 252789
rect 82486 252786 82492 252788
rect 82446 252726 82492 252786
rect 82556 252784 82603 252788
rect 82598 252728 82603 252784
rect 82486 252724 82492 252726
rect 82556 252724 82603 252728
rect 82537 252723 82603 252724
rect 77702 252316 77708 252380
rect 77772 252378 77778 252380
rect 78254 252378 78260 252380
rect 77772 252318 78260 252378
rect 77772 252316 77778 252318
rect 78254 252316 78260 252318
rect 78324 252316 78330 252380
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect 501638 251908 501644 251972
rect 501708 251970 501714 251972
rect 504030 251970 504036 251972
rect 501708 251910 504036 251970
rect 501708 251908 501714 251910
rect 504030 251908 504036 251910
rect 504100 251908 504106 251972
rect 501638 251772 501644 251836
rect 501708 251834 501714 251836
rect 502190 251834 502196 251836
rect 501708 251774 502196 251834
rect 501708 251772 501714 251774
rect 502190 251772 502196 251774
rect 502260 251772 502266 251836
rect -960 251290 480 251380
rect 3325 251290 3391 251293
rect -960 251288 3391 251290
rect -960 251232 3330 251288
rect 3386 251232 3391 251288
rect -960 251230 3391 251232
rect -960 251140 480 251230
rect 3325 251227 3391 251230
rect 507669 249930 507735 249933
rect 501860 249928 507735 249930
rect 501860 249872 507674 249928
rect 507730 249872 507735 249928
rect 501860 249870 507735 249872
rect 507669 249867 507735 249870
rect 503478 249732 503484 249796
rect 503548 249794 503554 249796
rect 504214 249794 504220 249796
rect 503548 249734 504220 249794
rect 503548 249732 503554 249734
rect 504214 249732 504220 249734
rect 504284 249732 504290 249796
rect 76005 249658 76071 249661
rect 76005 249656 82156 249658
rect 76005 249600 76010 249656
rect 76066 249600 82156 249656
rect 76005 249598 82156 249600
rect 76005 249595 76071 249598
rect 501270 249596 501276 249660
rect 501340 249658 501346 249660
rect 504398 249658 504404 249660
rect 501340 249598 504404 249658
rect 501340 249596 501346 249598
rect 504398 249596 504404 249598
rect 504468 249596 504474 249660
rect 501454 249324 501460 249388
rect 501524 249324 501530 249388
rect 501462 249116 501522 249324
rect 501454 249052 501460 249116
rect 501524 249052 501530 249116
rect 88701 248028 88767 248029
rect 88701 248026 88748 248028
rect 88656 248024 88748 248026
rect 88656 247968 88706 248024
rect 88656 247966 88748 247968
rect 88701 247964 88748 247966
rect 88812 247964 88818 248028
rect 88701 247963 88767 247964
rect 77385 247890 77451 247893
rect 77518 247890 77524 247892
rect 77385 247888 77524 247890
rect 77385 247832 77390 247888
rect 77446 247832 77524 247888
rect 77385 247830 77524 247832
rect 77385 247827 77451 247830
rect 77518 247828 77524 247830
rect 77588 247828 77594 247892
rect 88425 247756 88491 247757
rect 88374 247692 88380 247756
rect 88444 247754 88491 247756
rect 88444 247752 88536 247754
rect 88486 247696 88536 247752
rect 88444 247694 88536 247696
rect 88444 247692 88491 247694
rect 88425 247691 88491 247692
rect 501454 246604 501460 246668
rect 501524 246666 501530 246668
rect 503437 246666 503503 246669
rect 501524 246664 503503 246666
rect 501524 246608 503442 246664
rect 503498 246608 503503 246664
rect 501524 246606 503503 246608
rect 501524 246604 501530 246606
rect 503437 246603 503503 246606
rect 504214 246468 504220 246532
rect 504284 246530 504290 246532
rect 504633 246530 504699 246533
rect 504284 246528 504699 246530
rect 504284 246472 504638 246528
rect 504694 246472 504699 246528
rect 504284 246470 504699 246472
rect 504284 246468 504290 246470
rect 504633 246467 504699 246470
rect 510429 246394 510495 246397
rect 501860 246392 510495 246394
rect 501860 246336 510434 246392
rect 510490 246336 510495 246392
rect 501860 246334 510495 246336
rect 510429 246331 510495 246334
rect 82310 245581 82370 246092
rect 501454 246060 501460 246124
rect 501524 246122 501530 246124
rect 504030 246122 504036 246124
rect 501524 246062 504036 246122
rect 501524 246060 501530 246062
rect 504030 246060 504036 246062
rect 504100 246060 504106 246124
rect 82310 245576 82419 245581
rect 82310 245520 82358 245576
rect 82414 245520 82419 245576
rect 82310 245518 82419 245520
rect 82353 245515 82419 245518
rect 502190 244898 502196 244900
rect 501278 244838 502196 244898
rect 501278 244354 501338 244838
rect 502190 244836 502196 244838
rect 502260 244836 502266 244900
rect 502190 244700 502196 244764
rect 502260 244762 502266 244764
rect 504633 244762 504699 244765
rect 502260 244760 504699 244762
rect 502260 244704 504638 244760
rect 504694 244704 504699 244760
rect 502260 244702 504699 244704
rect 502260 244700 502266 244702
rect 504633 244699 504699 244702
rect 501454 244564 501460 244628
rect 501524 244626 501530 244628
rect 501822 244626 501828 244628
rect 501524 244566 501828 244626
rect 501524 244564 501530 244566
rect 501822 244564 501828 244566
rect 501892 244564 501898 244628
rect 501454 244428 501460 244492
rect 501524 244490 501530 244492
rect 502006 244490 502012 244492
rect 501524 244430 502012 244490
rect 501524 244428 501530 244430
rect 502006 244428 502012 244430
rect 502076 244428 502082 244492
rect 501454 244354 501460 244356
rect 501278 244294 501460 244354
rect 501454 244292 501460 244294
rect 501524 244292 501530 244356
rect 502006 244156 502012 244220
rect 502076 244218 502082 244220
rect 503529 244218 503595 244221
rect 502076 244216 503595 244218
rect 502076 244160 503534 244216
rect 503590 244160 503595 244216
rect 502076 244158 503595 244160
rect 502076 244156 502082 244158
rect 503529 244155 503595 244158
rect 503529 243130 503595 243133
rect 501860 243128 503595 243130
rect 501860 243072 503534 243128
rect 503590 243072 503595 243128
rect 501860 243070 503595 243072
rect 503529 243067 503595 243070
rect 501638 242660 501644 242724
rect 501708 242722 501714 242724
rect 501708 242662 502074 242722
rect 501708 242660 501714 242662
rect 78254 242524 78260 242588
rect 78324 242586 78330 242588
rect 78324 242526 82156 242586
rect 78324 242524 78330 242526
rect 501270 242524 501276 242588
rect 501340 242524 501346 242588
rect 80421 241498 80487 241501
rect 81014 241498 81020 241500
rect 80421 241496 81020 241498
rect 80421 241440 80426 241496
rect 80482 241440 81020 241496
rect 80421 241438 81020 241440
rect 80421 241435 80487 241438
rect 81014 241436 81020 241438
rect 81084 241436 81090 241500
rect 501278 241498 501338 242524
rect 501454 242388 501460 242452
rect 501524 242450 501530 242452
rect 501524 242390 501706 242450
rect 501524 242388 501530 242390
rect 501454 242116 501460 242180
rect 501524 242178 501530 242180
rect 501646 242178 501706 242390
rect 501822 242252 501828 242316
rect 501892 242314 501898 242316
rect 502014 242314 502074 242662
rect 501892 242254 502074 242314
rect 501892 242252 501898 242254
rect 501524 242118 501706 242178
rect 501524 242116 501530 242118
rect 503478 242116 503484 242180
rect 503548 242178 503554 242180
rect 504030 242178 504036 242180
rect 503548 242118 504036 242178
rect 503548 242116 503554 242118
rect 504030 242116 504036 242118
rect 504100 242116 504106 242180
rect 507025 242178 507091 242181
rect 507342 242178 507348 242180
rect 507025 242176 507348 242178
rect 507025 242120 507030 242176
rect 507086 242120 507348 242176
rect 507025 242118 507348 242120
rect 507025 242115 507091 242118
rect 507342 242116 507348 242118
rect 507412 242116 507418 242180
rect 501638 241980 501644 242044
rect 501708 242042 501714 242044
rect 503478 242042 503484 242044
rect 501708 241982 503484 242042
rect 501708 241980 501714 241982
rect 503478 241980 503484 241982
rect 503548 241980 503554 242044
rect 501454 241708 501460 241772
rect 501524 241770 501530 241772
rect 507526 241770 507532 241772
rect 501524 241710 507532 241770
rect 501524 241708 501530 241710
rect 507526 241708 507532 241710
rect 507596 241708 507602 241772
rect 524413 241770 524479 241773
rect 524278 241768 524479 241770
rect 524278 241712 524418 241768
rect 524474 241712 524479 241768
rect 524278 241710 524479 241712
rect 524278 241634 524338 241710
rect 524413 241707 524479 241710
rect 524413 241634 524479 241637
rect 524278 241632 524479 241634
rect 524278 241576 524418 241632
rect 524474 241576 524479 241632
rect 524278 241574 524479 241576
rect 524413 241571 524479 241574
rect 501454 241498 501460 241500
rect 501278 241438 501460 241498
rect 501454 241436 501460 241438
rect 501524 241436 501530 241500
rect 501638 241436 501644 241500
rect 501708 241498 501714 241500
rect 503437 241498 503503 241501
rect 501708 241496 503503 241498
rect 501708 241440 503442 241496
rect 503498 241440 503503 241496
rect 501708 241438 503503 241440
rect 501708 241436 501714 241438
rect 503437 241435 503503 241438
rect 80830 241362 80836 241364
rect 80654 241302 80836 241362
rect 80654 240818 80714 241302
rect 80830 241300 80836 241302
rect 80900 241300 80906 241364
rect 81198 241300 81204 241364
rect 81268 241300 81274 241364
rect 81382 241300 81388 241364
rect 81452 241300 81458 241364
rect 81206 240820 81266 241300
rect 81390 240820 81450 241300
rect 80830 240818 80836 240820
rect 80654 240758 80836 240818
rect 80830 240756 80836 240758
rect 80900 240756 80906 240820
rect 81198 240756 81204 240820
rect 81268 240756 81274 240820
rect 81382 240756 81388 240820
rect 81452 240756 81458 240820
rect 583520 240396 584960 240636
rect 524413 240138 524479 240141
rect 524597 240138 524663 240141
rect 524413 240136 524663 240138
rect 524413 240080 524418 240136
rect 524474 240080 524602 240136
rect 524658 240080 524663 240136
rect 524413 240078 524663 240080
rect 524413 240075 524479 240078
rect 524597 240075 524663 240078
rect 503437 239594 503503 239597
rect 501860 239592 503503 239594
rect 501860 239536 503442 239592
rect 503498 239536 503503 239592
rect 501860 239534 503503 239536
rect 503437 239531 503503 239534
rect 80421 239458 80487 239461
rect 82537 239460 82603 239461
rect 81014 239458 81020 239460
rect 80421 239456 81020 239458
rect 80421 239400 80426 239456
rect 80482 239400 81020 239456
rect 80421 239398 81020 239400
rect 80421 239395 80487 239398
rect 81014 239396 81020 239398
rect 81084 239396 81090 239460
rect 82532 239458 82538 239460
rect 82446 239398 82538 239458
rect 82532 239396 82538 239398
rect 82602 239396 82608 239460
rect 82537 239395 82603 239396
rect 81433 239050 81499 239053
rect 504398 239050 504404 239052
rect 81433 239048 82156 239050
rect 81433 238992 81438 239048
rect 81494 238992 82156 239048
rect 81433 238990 82156 238992
rect 501278 238990 504404 239050
rect 81433 238987 81499 238990
rect 82445 238372 82511 238373
rect 82445 238370 82492 238372
rect 82400 238368 82492 238370
rect 82400 238312 82450 238368
rect 82400 238310 82492 238312
rect 82445 238308 82492 238310
rect 82556 238308 82562 238372
rect 82445 238307 82511 238308
rect 501278 238100 501338 238990
rect 504398 238988 504404 238990
rect 504468 238988 504474 239052
rect 529933 238914 529999 238917
rect 539501 238914 539567 238917
rect 529933 238912 539567 238914
rect 529933 238856 529938 238912
rect 529994 238856 539506 238912
rect 539562 238856 539567 238912
rect 529933 238854 539567 238856
rect 529933 238851 529999 238854
rect 539501 238851 539567 238854
rect 501270 238036 501276 238100
rect 501340 238036 501346 238100
rect 501822 238036 501828 238100
rect 501892 238098 501898 238100
rect 503437 238098 503503 238101
rect 501892 238096 503503 238098
rect 501892 238040 503442 238096
rect 503498 238040 503503 238096
rect 501892 238038 503503 238040
rect 501892 238036 501898 238038
rect 503437 238035 503503 238038
rect 501454 237764 501460 237828
rect 501524 237764 501530 237828
rect 501638 237764 501644 237828
rect 501708 237764 501714 237828
rect 77385 237690 77451 237693
rect 78070 237690 78076 237692
rect 77385 237688 78076 237690
rect 77385 237632 77390 237688
rect 77446 237632 78076 237688
rect 77385 237630 78076 237632
rect 77385 237627 77451 237630
rect 78070 237628 78076 237630
rect 78140 237628 78146 237692
rect 501462 237556 501522 237764
rect 501646 237556 501706 237764
rect 501822 237628 501828 237692
rect 501892 237690 501898 237692
rect 503529 237690 503595 237693
rect 501892 237688 503595 237690
rect 501892 237632 503534 237688
rect 503590 237632 503595 237688
rect 501892 237630 503595 237632
rect 501892 237628 501898 237630
rect 503529 237627 503595 237630
rect 501454 237492 501460 237556
rect 501524 237492 501530 237556
rect 501638 237492 501644 237556
rect 501708 237492 501714 237556
rect 501270 237220 501276 237284
rect 501340 237282 501346 237284
rect 501822 237282 501828 237284
rect 501340 237222 501828 237282
rect 501340 237220 501346 237222
rect 501822 237220 501828 237222
rect 501892 237220 501898 237284
rect -960 237010 480 237100
rect 3233 237010 3299 237013
rect 80329 237012 80395 237013
rect 80278 237010 80284 237012
rect -960 237008 3299 237010
rect -960 236952 3238 237008
rect 3294 236952 3299 237008
rect -960 236950 3299 236952
rect 80238 236950 80284 237010
rect 80348 237008 80395 237012
rect 80390 236952 80395 237008
rect -960 236860 480 236950
rect 3233 236947 3299 236950
rect 80278 236948 80284 236950
rect 80348 236948 80395 236952
rect 82486 236948 82492 237012
rect 82556 237010 82562 237012
rect 82629 237010 82695 237013
rect 82556 237008 82695 237010
rect 82556 236952 82634 237008
rect 82690 236952 82695 237008
rect 82556 236950 82695 236952
rect 82556 236948 82562 236950
rect 80329 236947 80395 236948
rect 82629 236947 82695 236950
rect 80329 236194 80395 236197
rect 82486 236194 82492 236196
rect 80329 236192 82492 236194
rect 80329 236136 80334 236192
rect 80390 236136 82492 236192
rect 80329 236134 82492 236136
rect 80329 236131 80395 236134
rect 82486 236132 82492 236134
rect 82556 236132 82562 236196
rect 504633 236058 504699 236061
rect 501860 236056 504699 236058
rect 501860 236000 504638 236056
rect 504694 236000 504699 236056
rect 501860 235998 504699 236000
rect 504633 235995 504699 235998
rect 501270 235724 501276 235788
rect 501340 235786 501346 235788
rect 503529 235786 503595 235789
rect 501340 235784 503595 235786
rect 501340 235728 503534 235784
rect 503590 235728 503595 235784
rect 501340 235726 503595 235728
rect 501340 235724 501346 235726
rect 503529 235723 503595 235726
rect 501270 235588 501276 235652
rect 501340 235650 501346 235652
rect 503478 235650 503484 235652
rect 501340 235590 503484 235650
rect 501340 235588 501346 235590
rect 503478 235588 503484 235590
rect 503548 235588 503554 235652
rect 503529 235514 503595 235517
rect 504582 235514 504588 235516
rect 503529 235512 504588 235514
rect 82445 235108 82511 235109
rect 82445 235106 82492 235108
rect 82400 235104 82492 235106
rect 82400 235048 82450 235104
rect 82400 235046 82492 235048
rect 82445 235044 82492 235046
rect 82556 235044 82562 235108
rect 82445 235043 82511 235044
rect 82445 234970 82511 234973
rect 82678 234970 82738 235484
rect 503529 235456 503534 235512
rect 503590 235456 504588 235512
rect 503529 235454 504588 235456
rect 503529 235451 503595 235454
rect 504582 235452 504588 235454
rect 504652 235452 504658 235516
rect 507025 235380 507091 235381
rect 504030 235316 504036 235380
rect 504100 235378 504106 235380
rect 504582 235378 504588 235380
rect 504100 235318 504588 235378
rect 504100 235316 504106 235318
rect 504582 235316 504588 235318
rect 504652 235316 504658 235380
rect 506974 235378 506980 235380
rect 506934 235318 506980 235378
rect 507044 235376 507091 235380
rect 507086 235320 507091 235376
rect 506974 235316 506980 235318
rect 507044 235316 507091 235320
rect 507025 235315 507091 235316
rect 82445 234968 82738 234970
rect 82445 234912 82450 234968
rect 82506 234912 82738 234968
rect 82445 234910 82738 234912
rect 82445 234907 82511 234910
rect 82486 234772 82492 234836
rect 82556 234834 82562 234836
rect 82629 234834 82695 234837
rect 82556 234832 82695 234834
rect 82556 234776 82634 234832
rect 82690 234776 82695 234832
rect 82556 234774 82695 234776
rect 82556 234772 82562 234774
rect 82629 234771 82695 234774
rect 81433 233746 81499 233749
rect 82486 233746 82492 233748
rect 81433 233744 82492 233746
rect 81433 233688 81438 233744
rect 81494 233688 82492 233744
rect 81433 233686 82492 233688
rect 81433 233683 81499 233686
rect 82486 233684 82492 233686
rect 82556 233684 82562 233748
rect 82486 233412 82492 233476
rect 82556 233474 82562 233476
rect 82629 233474 82695 233477
rect 82556 233472 82695 233474
rect 82556 233416 82634 233472
rect 82690 233416 82695 233472
rect 82556 233414 82695 233416
rect 82556 233412 82562 233414
rect 82629 233411 82695 233414
rect 502006 233140 502012 233204
rect 502076 233202 502082 233204
rect 503529 233202 503595 233205
rect 502076 233200 503595 233202
rect 502076 233144 503534 233200
rect 503590 233144 503595 233200
rect 502076 233142 503595 233144
rect 502076 233140 502082 233142
rect 503529 233139 503595 233142
rect 88701 233068 88767 233069
rect 88701 233066 88748 233068
rect 88656 233064 88748 233066
rect 88656 233008 88706 233064
rect 88656 233006 88748 233008
rect 88701 233004 88748 233006
rect 88812 233004 88818 233068
rect 88701 233003 88767 233004
rect 87873 232796 87939 232797
rect 87822 232732 87828 232796
rect 87892 232794 87939 232796
rect 87892 232792 87984 232794
rect 87934 232736 87984 232792
rect 87892 232734 87984 232736
rect 87892 232732 87939 232734
rect 87873 232731 87939 232732
rect 82302 232596 82308 232660
rect 82372 232596 82378 232660
rect 82486 232596 82492 232660
rect 82556 232658 82562 232660
rect 82629 232658 82695 232661
rect 82556 232656 82695 232658
rect 82556 232600 82634 232656
rect 82690 232600 82695 232656
rect 82556 232598 82695 232600
rect 82556 232596 82562 232598
rect 82310 232386 82370 232596
rect 82629 232595 82695 232598
rect 506013 232522 506079 232525
rect 501860 232520 506079 232522
rect 501860 232464 506018 232520
rect 506074 232464 506079 232520
rect 501860 232462 506079 232464
rect 506013 232459 506079 232462
rect 82537 232386 82603 232389
rect 82310 232384 82603 232386
rect 82310 232328 82542 232384
rect 82598 232328 82603 232384
rect 82310 232326 82603 232328
rect 82537 232323 82603 232326
rect 78949 231978 79015 231981
rect 78949 231976 82156 231978
rect 78949 231920 78954 231976
rect 79010 231920 82156 231976
rect 78949 231918 82156 231920
rect 78949 231915 79015 231918
rect 502374 231780 502380 231844
rect 502444 231780 502450 231844
rect 502382 231300 502442 231780
rect 502374 231236 502380 231300
rect 502444 231236 502450 231300
rect 82486 230964 82492 231028
rect 82556 231026 82562 231028
rect 82556 230966 82738 231026
rect 82556 230964 82562 230966
rect 78254 230828 78260 230892
rect 78324 230890 78330 230892
rect 82486 230890 82492 230892
rect 78324 230830 82492 230890
rect 78324 230828 78330 230830
rect 82486 230828 82492 230830
rect 82556 230828 82562 230892
rect 82302 230556 82308 230620
rect 82372 230618 82378 230620
rect 82678 230618 82738 230966
rect 82372 230558 82738 230618
rect 82372 230556 82378 230558
rect 81433 229530 81499 229533
rect 82486 229530 82492 229532
rect 81433 229528 82492 229530
rect 81433 229472 81438 229528
rect 81494 229472 82492 229528
rect 81433 229470 82492 229472
rect 81433 229467 81499 229470
rect 82486 229468 82492 229470
rect 82556 229468 82562 229532
rect 81433 229258 81499 229261
rect 82486 229258 82492 229260
rect 81433 229256 82492 229258
rect 81433 229200 81438 229256
rect 81494 229200 82492 229256
rect 81433 229198 82492 229200
rect 81433 229195 81499 229198
rect 82486 229196 82492 229198
rect 82556 229196 82562 229260
rect 503345 229122 503411 229125
rect 503478 229122 503484 229124
rect 503345 229120 503484 229122
rect 503345 229064 503350 229120
rect 503406 229064 503484 229120
rect 503345 229062 503484 229064
rect 503345 229059 503411 229062
rect 503478 229060 503484 229062
rect 503548 229060 503554 229124
rect 503345 228986 503411 228989
rect 501860 228984 503411 228986
rect 501860 228928 503350 228984
rect 503406 228928 503411 228984
rect 501860 228926 503411 228928
rect 503345 228923 503411 228926
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 76557 228442 76623 228445
rect 76557 228440 82156 228442
rect 76557 228384 76562 228440
rect 76618 228384 82156 228440
rect 76557 228382 82156 228384
rect 76557 228379 76623 228382
rect 81433 227898 81499 227901
rect 82486 227898 82492 227900
rect 81433 227896 82492 227898
rect 81433 227840 81438 227896
rect 81494 227840 82492 227896
rect 81433 227838 82492 227840
rect 81433 227835 81499 227838
rect 82486 227836 82492 227838
rect 82556 227836 82562 227900
rect 84561 226812 84627 226813
rect 84510 226748 84516 226812
rect 84580 226810 84627 226812
rect 86125 226812 86191 226813
rect 84580 226808 84672 226810
rect 84622 226752 84672 226808
rect 84580 226750 84672 226752
rect 86125 226808 86172 226812
rect 86236 226810 86242 226812
rect 86125 226752 86130 226808
rect 84580 226748 84627 226750
rect 84561 226747 84627 226748
rect 86125 226748 86172 226752
rect 86236 226750 86282 226810
rect 86236 226748 86242 226750
rect 86125 226747 86191 226748
rect 501822 226612 501828 226676
rect 501892 226674 501898 226676
rect 502190 226674 502196 226676
rect 501892 226614 502196 226674
rect 501892 226612 501898 226614
rect 502190 226612 502196 226614
rect 502260 226612 502266 226676
rect 502190 226476 502196 226540
rect 502260 226538 502266 226540
rect 503621 226538 503687 226541
rect 502260 226536 503687 226538
rect 502260 226480 503626 226536
rect 503682 226480 503687 226536
rect 502260 226478 503687 226480
rect 502260 226476 502266 226478
rect 503621 226475 503687 226478
rect 82302 225660 82308 225724
rect 82372 225722 82378 225724
rect 82629 225722 82695 225725
rect 82372 225720 82695 225722
rect 82372 225664 82634 225720
rect 82690 225664 82695 225720
rect 82372 225662 82695 225664
rect 82372 225660 82378 225662
rect 82629 225659 82695 225662
rect 503437 225450 503503 225453
rect 501860 225448 503503 225450
rect 501860 225392 503442 225448
rect 503498 225392 503503 225448
rect 501860 225390 503503 225392
rect 503437 225387 503503 225390
rect 501270 225116 501276 225180
rect 501340 225178 501346 225180
rect 503621 225178 503687 225181
rect 501340 225176 503687 225178
rect 501340 225120 503626 225176
rect 503682 225120 503687 225176
rect 501340 225118 503687 225120
rect 501340 225116 501346 225118
rect 503621 225115 503687 225118
rect 82678 224365 82738 224876
rect 501270 224844 501276 224908
rect 501340 224906 501346 224908
rect 503437 224906 503503 224909
rect 501340 224904 503503 224906
rect 501340 224848 503442 224904
rect 503498 224848 503503 224904
rect 501340 224846 503503 224848
rect 501340 224844 501346 224846
rect 503437 224843 503503 224846
rect 82629 224360 82738 224365
rect 82629 224304 82634 224360
rect 82690 224304 82738 224360
rect 82629 224302 82738 224304
rect 82629 224299 82695 224302
rect 501454 223682 501460 223684
rect 501278 223622 501460 223682
rect 81433 223410 81499 223413
rect 82486 223410 82492 223412
rect 81433 223408 82492 223410
rect 81433 223352 81438 223408
rect 81494 223352 82492 223408
rect 81433 223350 82492 223352
rect 81433 223347 81499 223350
rect 82486 223348 82492 223350
rect 82556 223348 82562 223412
rect -960 222594 480 222684
rect 3325 222594 3391 222597
rect -960 222592 3391 222594
rect -960 222536 3330 222592
rect 3386 222536 3391 222592
rect -960 222534 3391 222536
rect 501278 222594 501338 223622
rect 501454 223620 501460 223622
rect 501524 223620 501530 223684
rect 501454 222594 501460 222596
rect 501278 222534 501460 222594
rect -960 222444 480 222534
rect 3325 222531 3391 222534
rect 501454 222532 501460 222534
rect 501524 222532 501530 222596
rect 501270 222124 501276 222188
rect 501340 222186 501346 222188
rect 501340 222126 504650 222186
rect 501340 222124 501346 222126
rect 503437 222050 503503 222053
rect 503437 222048 503684 222050
rect 503437 221992 503442 222048
rect 503498 221992 503684 222048
rect 503437 221990 503684 221992
rect 503437 221987 503503 221990
rect 503437 221914 503503 221917
rect 501860 221912 503503 221914
rect 501860 221856 503442 221912
rect 503498 221856 503503 221912
rect 501860 221854 503503 221856
rect 503437 221851 503503 221854
rect 501270 221580 501276 221644
rect 501340 221642 501346 221644
rect 503624 221642 503684 221990
rect 504030 221988 504036 222052
rect 504100 222050 504106 222052
rect 504398 222050 504404 222052
rect 504100 221990 504404 222050
rect 504100 221988 504106 221990
rect 504398 221988 504404 221990
rect 504468 221988 504474 222052
rect 504590 221916 504650 222126
rect 504582 221852 504588 221916
rect 504652 221852 504658 221916
rect 501340 221582 503684 221642
rect 501340 221580 501346 221582
rect 501270 221444 501276 221508
rect 501340 221506 501346 221508
rect 501822 221506 501828 221508
rect 501340 221446 501828 221506
rect 501340 221444 501346 221446
rect 501822 221444 501828 221446
rect 501892 221444 501898 221508
rect 502006 221444 502012 221508
rect 502076 221506 502082 221508
rect 503437 221506 503503 221509
rect 502076 221504 503503 221506
rect 502076 221448 503442 221504
rect 503498 221448 503503 221504
rect 502076 221446 503503 221448
rect 502076 221444 502082 221446
rect 503437 221443 503503 221446
rect 81525 221370 81591 221373
rect 81525 221368 82156 221370
rect 81525 221312 81530 221368
rect 81586 221312 82156 221368
rect 81525 221310 82156 221312
rect 81525 221307 81591 221310
rect 524413 220826 524479 220829
rect 524597 220826 524663 220829
rect 524413 220824 524663 220826
rect 524413 220768 524418 220824
rect 524474 220768 524602 220824
rect 524658 220768 524663 220824
rect 524413 220766 524663 220768
rect 524413 220763 524479 220766
rect 524597 220763 524663 220766
rect 503621 220418 503687 220421
rect 501278 220416 503687 220418
rect 501278 220360 503626 220416
rect 503682 220360 503687 220416
rect 501278 220358 503687 220360
rect 82486 220084 82492 220148
rect 82556 220146 82562 220148
rect 82556 220086 82738 220146
rect 82556 220084 82562 220086
rect 78254 219948 78260 220012
rect 78324 220010 78330 220012
rect 82486 220010 82492 220012
rect 78324 219950 82492 220010
rect 78324 219948 78330 219950
rect 82486 219948 82492 219950
rect 82556 219948 82562 220012
rect 82486 219812 82492 219876
rect 82556 219874 82562 219876
rect 82678 219874 82738 220086
rect 82556 219814 82738 219874
rect 82556 219812 82562 219814
rect 501278 219738 501338 220358
rect 503621 220355 503687 220358
rect 501454 220220 501460 220284
rect 501524 220282 501530 220284
rect 503621 220282 503687 220285
rect 501524 220280 503687 220282
rect 501524 220224 503626 220280
rect 503682 220224 503687 220280
rect 501524 220222 503687 220224
rect 501524 220220 501530 220222
rect 503621 220219 503687 220222
rect 501822 219948 501828 220012
rect 501892 220010 501898 220012
rect 502190 220010 502196 220012
rect 501892 219950 502196 220010
rect 501892 219948 501898 219950
rect 502190 219948 502196 219950
rect 502260 219948 502266 220012
rect 502190 219812 502196 219876
rect 502260 219874 502266 219876
rect 503529 219874 503595 219877
rect 502260 219872 503595 219874
rect 502260 219816 503534 219872
rect 503590 219816 503595 219872
rect 502260 219814 503595 219816
rect 502260 219812 502266 219814
rect 503529 219811 503595 219814
rect 501454 219738 501460 219740
rect 501278 219678 501460 219738
rect 501454 219676 501460 219678
rect 501524 219676 501530 219740
rect 506933 218378 506999 218381
rect 501860 218376 506999 218378
rect 501860 218320 506938 218376
rect 506994 218320 506999 218376
rect 501860 218318 506999 218320
rect 506933 218315 506999 218318
rect 80329 217834 80395 217837
rect 80329 217832 82156 217834
rect 80329 217776 80334 217832
rect 80390 217776 82156 217832
rect 80329 217774 82156 217776
rect 80329 217771 80395 217774
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 502006 216276 502012 216340
rect 502076 216276 502082 216340
rect 502014 216202 502074 216276
rect 502014 216142 502258 216202
rect 502198 216066 502258 216142
rect 503621 216066 503687 216069
rect 502198 216064 503687 216066
rect 502198 216008 503626 216064
rect 503682 216008 503687 216064
rect 502198 216006 503687 216008
rect 503621 216003 503687 216006
rect 501454 215868 501460 215932
rect 501524 215930 501530 215932
rect 503529 215930 503595 215933
rect 501524 215928 503595 215930
rect 501524 215872 503534 215928
rect 503590 215872 503595 215928
rect 501524 215870 503595 215872
rect 501524 215868 501530 215870
rect 503529 215867 503595 215870
rect 502190 215732 502196 215796
rect 502260 215794 502266 215796
rect 503529 215794 503595 215797
rect 502260 215792 503595 215794
rect 502260 215736 503534 215792
rect 503590 215736 503595 215792
rect 502260 215734 503595 215736
rect 502260 215732 502266 215734
rect 503529 215731 503595 215734
rect 509049 214842 509115 214845
rect 501860 214840 509115 214842
rect 501860 214784 509054 214840
rect 509110 214784 509115 214840
rect 501860 214782 509115 214784
rect 509049 214779 509115 214782
rect 504030 214508 504036 214572
rect 504100 214570 504106 214572
rect 504398 214570 504404 214572
rect 504100 214510 504404 214570
rect 504100 214508 504106 214510
rect 504398 214508 504404 214510
rect 504468 214508 504474 214572
rect 81525 214298 81591 214301
rect 81525 214296 82156 214298
rect 81525 214240 81530 214296
rect 81586 214240 82156 214296
rect 81525 214238 82156 214240
rect 81525 214235 81591 214238
rect 502190 211788 502196 211852
rect 502260 211850 502266 211852
rect 503437 211850 503503 211853
rect 502260 211848 503503 211850
rect 502260 211792 503442 211848
rect 503498 211792 503503 211848
rect 502260 211790 503503 211792
rect 502260 211788 502266 211790
rect 503437 211787 503503 211790
rect 501270 211516 501276 211580
rect 501340 211578 501346 211580
rect 504582 211578 504588 211580
rect 501340 211518 504588 211578
rect 501340 211516 501346 211518
rect 504582 211516 504588 211518
rect 504652 211516 504658 211580
rect 503437 211306 503503 211309
rect 501860 211304 503503 211306
rect 501860 211248 503442 211304
rect 503498 211248 503503 211304
rect 501860 211246 503503 211248
rect 503437 211243 503503 211246
rect 524413 211170 524479 211173
rect 524597 211170 524663 211173
rect 524413 211168 524663 211170
rect 524413 211112 524418 211168
rect 524474 211112 524602 211168
rect 524658 211112 524663 211168
rect 524413 211110 524663 211112
rect 524413 211107 524479 211110
rect 524597 211107 524663 211110
rect 79409 210762 79475 210765
rect 503621 210762 503687 210765
rect 504030 210762 504036 210764
rect 79409 210760 82156 210762
rect 79409 210704 79414 210760
rect 79470 210704 82156 210760
rect 79409 210702 82156 210704
rect 503621 210760 504036 210762
rect 503621 210704 503626 210760
rect 503682 210704 504036 210760
rect 503621 210702 504036 210704
rect 79409 210699 79475 210702
rect 503621 210699 503687 210702
rect 504030 210700 504036 210702
rect 504100 210700 504106 210764
rect 81525 210490 81591 210493
rect 82624 210490 82630 210492
rect 81525 210488 82630 210490
rect 81525 210432 81530 210488
rect 81586 210432 82630 210488
rect 81525 210430 82630 210432
rect 81525 210427 81591 210430
rect 82624 210428 82630 210430
rect 82694 210428 82700 210492
rect 82302 209340 82308 209404
rect 82372 209402 82378 209404
rect 82629 209402 82695 209405
rect 82372 209400 82695 209402
rect 82372 209344 82634 209400
rect 82690 209344 82695 209400
rect 82372 209342 82695 209344
rect 82372 209340 82378 209342
rect 82629 209339 82695 209342
rect 502006 209204 502012 209268
rect 502076 209266 502082 209268
rect 502149 209266 502215 209269
rect 502076 209264 502215 209266
rect 502076 209208 502154 209264
rect 502210 209208 502215 209264
rect 502076 209206 502215 209208
rect 502076 209204 502082 209206
rect 502149 209203 502215 209206
rect 80145 209130 80211 209133
rect 82486 209130 82492 209132
rect 80145 209128 82492 209130
rect 80145 209072 80150 209128
rect 80206 209072 82492 209128
rect 80145 209070 82492 209072
rect 80145 209067 80211 209070
rect 82486 209068 82492 209070
rect 82556 209068 82562 209132
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 81433 208042 81499 208045
rect 82302 208042 82308 208044
rect 81433 208040 82308 208042
rect 81433 207984 81438 208040
rect 81494 207984 82308 208040
rect 81433 207982 82308 207984
rect 81433 207979 81499 207982
rect 82302 207980 82308 207982
rect 82372 207980 82378 208044
rect 80237 207770 80303 207773
rect 82624 207770 82630 207772
rect 80237 207768 82630 207770
rect 80237 207712 80242 207768
rect 80298 207712 82630 207768
rect 80237 207710 82630 207712
rect 80237 207707 80303 207710
rect 82624 207708 82630 207710
rect 82694 207708 82700 207772
rect 503621 207770 503687 207773
rect 501860 207768 503687 207770
rect 501860 207712 503626 207768
rect 503682 207712 503687 207768
rect 501860 207710 503687 207712
rect 503621 207707 503687 207710
rect 81525 207226 81591 207229
rect 81525 207224 82156 207226
rect 81525 207168 81530 207224
rect 81586 207168 82156 207224
rect 81525 207166 82156 207168
rect 81525 207163 81591 207166
rect 77702 206212 77708 206276
rect 77772 206274 77778 206276
rect 78254 206274 78260 206276
rect 77772 206214 78260 206274
rect 77772 206212 77778 206214
rect 78254 206212 78260 206214
rect 78324 206212 78330 206276
rect 77518 206076 77524 206140
rect 77588 206138 77594 206140
rect 78254 206138 78260 206140
rect 77588 206078 78260 206138
rect 77588 206076 77594 206078
rect 78254 206076 78260 206078
rect 78324 206076 78330 206140
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect 501454 204852 501460 204916
rect 501524 204914 501530 204916
rect 503529 204914 503595 204917
rect 501524 204912 503595 204914
rect 501524 204856 503534 204912
rect 503590 204856 503595 204912
rect 501524 204854 503595 204856
rect 501524 204852 501530 204854
rect 503529 204851 503595 204854
rect 507025 204234 507091 204237
rect 501860 204232 507091 204234
rect 501860 204176 507030 204232
rect 507086 204176 507091 204232
rect 501860 204174 507091 204176
rect 507025 204171 507091 204174
rect 502144 204036 502150 204100
rect 502214 204098 502220 204100
rect 503529 204098 503595 204101
rect 502214 204096 503595 204098
rect 502214 204040 503534 204096
rect 503590 204040 503595 204096
rect 502214 204038 503595 204040
rect 502214 204036 502220 204038
rect 503529 204035 503595 204038
rect 80329 203690 80395 203693
rect 80329 203688 82156 203690
rect 80329 203632 80334 203688
rect 80390 203632 82156 203688
rect 80329 203630 82156 203632
rect 80329 203627 80395 203630
rect 501270 203628 501276 203692
rect 501340 203628 501346 203692
rect 501278 203148 501338 203628
rect 501454 203356 501460 203420
rect 501524 203418 501530 203420
rect 504582 203418 504588 203420
rect 501524 203358 504588 203418
rect 501524 203356 501530 203358
rect 504582 203356 504588 203358
rect 504652 203356 504658 203420
rect 501454 203220 501460 203284
rect 501524 203282 501530 203284
rect 502006 203282 502012 203284
rect 501524 203222 502012 203282
rect 501524 203220 501530 203222
rect 502006 203220 502012 203222
rect 502076 203220 502082 203284
rect 77886 203084 77892 203148
rect 77956 203146 77962 203148
rect 77956 203086 82370 203146
rect 77956 203084 77962 203086
rect 79133 203010 79199 203013
rect 80421 203010 80487 203013
rect 79133 203008 80487 203010
rect 79133 202952 79138 203008
rect 79194 202952 80426 203008
rect 80482 202952 80487 203008
rect 79133 202950 80487 202952
rect 82310 203010 82370 203086
rect 82486 203084 82492 203148
rect 82556 203146 82562 203148
rect 82556 203086 82738 203146
rect 82556 203084 82562 203086
rect 82486 203010 82492 203012
rect 82310 202950 82492 203010
rect 79133 202947 79199 202950
rect 80421 202947 80487 202950
rect 82486 202948 82492 202950
rect 82556 202948 82562 203012
rect 78070 202676 78076 202740
rect 78140 202738 78146 202740
rect 80145 202738 80211 202741
rect 78140 202736 80211 202738
rect 78140 202680 80150 202736
rect 80206 202680 80211 202736
rect 78140 202678 80211 202680
rect 78140 202676 78146 202678
rect 80145 202675 80211 202678
rect 80145 202058 80211 202061
rect 82486 202058 82492 202060
rect 80145 202056 82492 202058
rect 80145 202000 80150 202056
rect 80206 202000 82492 202056
rect 80145 201998 82492 202000
rect 80145 201995 80211 201998
rect 82486 201996 82492 201998
rect 82556 201996 82562 202060
rect 76373 201922 76439 201925
rect 77150 201922 77156 201924
rect 76373 201920 77156 201922
rect 76373 201864 76378 201920
rect 76434 201864 77156 201920
rect 76373 201862 77156 201864
rect 76373 201859 76439 201862
rect 77150 201860 77156 201862
rect 77220 201860 77226 201924
rect 81525 201922 81591 201925
rect 82486 201922 82492 201924
rect 81525 201920 82492 201922
rect 81525 201864 81530 201920
rect 81586 201864 82492 201920
rect 81525 201862 82492 201864
rect 81525 201859 81591 201862
rect 82486 201860 82492 201862
rect 82556 201860 82562 201924
rect 82486 201724 82492 201788
rect 82556 201786 82562 201788
rect 82678 201786 82738 203086
rect 501270 203084 501276 203148
rect 501340 203084 501346 203148
rect 501638 202132 501644 202196
rect 501708 202194 501714 202196
rect 502190 202194 502196 202196
rect 501708 202134 502196 202194
rect 501708 202132 501714 202134
rect 502190 202132 502196 202134
rect 502260 202132 502266 202196
rect 82556 201726 82738 201786
rect 82556 201724 82562 201726
rect 80237 201650 80303 201653
rect 82624 201650 82630 201652
rect 80237 201648 82630 201650
rect 80237 201592 80242 201648
rect 80298 201592 82630 201648
rect 80237 201590 82630 201592
rect 80237 201587 80303 201590
rect 82624 201588 82630 201590
rect 82694 201588 82700 201652
rect 82302 201452 82308 201516
rect 82372 201514 82378 201516
rect 82372 201454 82738 201514
rect 82372 201452 82378 201454
rect 81525 201242 81591 201245
rect 82302 201242 82308 201244
rect 81525 201240 82308 201242
rect 81525 201184 81530 201240
rect 81586 201184 82308 201240
rect 81525 201182 82308 201184
rect 81525 201179 81591 201182
rect 82302 201180 82308 201182
rect 82372 201180 82378 201244
rect 81525 201106 81591 201109
rect 82486 201106 82492 201108
rect 81525 201104 82492 201106
rect 81525 201048 81530 201104
rect 81586 201048 82492 201104
rect 81525 201046 82492 201048
rect 81525 201043 81591 201046
rect 82486 201044 82492 201046
rect 82556 201044 82562 201108
rect 76046 200908 76052 200972
rect 76116 200970 76122 200972
rect 77518 200970 77524 200972
rect 76116 200910 77524 200970
rect 76116 200908 76122 200910
rect 77518 200908 77524 200910
rect 77588 200908 77594 200972
rect 82302 200772 82308 200836
rect 82372 200834 82378 200836
rect 82678 200834 82738 201454
rect 501454 201180 501460 201244
rect 501524 201180 501530 201244
rect 82372 200774 82738 200834
rect 82372 200772 82378 200774
rect 501462 200668 501522 201180
rect 501270 200364 501276 200428
rect 501340 200426 501346 200428
rect 502006 200426 502012 200428
rect 501340 200366 502012 200426
rect 501340 200364 501346 200366
rect 502006 200364 502012 200366
rect 502076 200364 502082 200428
rect 2773 200290 2839 200293
rect 78254 200290 78260 200292
rect 2773 200288 78260 200290
rect 2773 200232 2778 200288
rect 2834 200232 78260 200288
rect 2773 200230 78260 200232
rect 2773 200227 2839 200230
rect 78254 200228 78260 200230
rect 78324 200228 78330 200292
rect 81433 200154 81499 200157
rect 81433 200152 82156 200154
rect 81433 200096 81438 200152
rect 81494 200096 82156 200152
rect 81433 200094 82156 200096
rect 81433 200091 81499 200094
rect 80145 199610 80211 199613
rect 82486 199610 82492 199612
rect 80145 199608 82492 199610
rect 80145 199552 80150 199608
rect 80206 199552 82492 199608
rect 80145 199550 82492 199552
rect 80145 199547 80211 199550
rect 82486 199548 82492 199550
rect 82556 199548 82562 199612
rect 501638 199412 501644 199476
rect 501708 199474 501714 199476
rect 504030 199474 504036 199476
rect 501708 199414 504036 199474
rect 501708 199412 501714 199414
rect 504030 199412 504036 199414
rect 504100 199412 504106 199476
rect 503621 199338 503687 199341
rect 504030 199338 504036 199340
rect 503621 199336 504036 199338
rect 503621 199280 503626 199336
rect 503682 199280 504036 199336
rect 503621 199278 504036 199280
rect 503621 199275 503687 199278
rect 504030 199276 504036 199278
rect 504100 199276 504106 199340
rect 76373 198114 76439 198117
rect 77150 198114 77156 198116
rect 76373 198112 77156 198114
rect 76373 198056 76378 198112
rect 76434 198056 77156 198112
rect 76373 198054 77156 198056
rect 76373 198051 76439 198054
rect 77150 198052 77156 198054
rect 77220 198052 77226 198116
rect 501822 198052 501828 198116
rect 501892 198114 501898 198116
rect 502149 198114 502215 198117
rect 501892 198112 502215 198114
rect 501892 198056 502154 198112
rect 502210 198056 502215 198112
rect 501892 198054 502215 198056
rect 501892 198052 501898 198054
rect 502149 198051 502215 198054
rect 502006 197372 502012 197436
rect 502076 197434 502082 197436
rect 503529 197434 503595 197437
rect 502076 197432 503595 197434
rect 502076 197376 503534 197432
rect 503590 197376 503595 197432
rect 502076 197374 503595 197376
rect 502076 197372 502082 197374
rect 503529 197371 503595 197374
rect 504817 197162 504883 197165
rect 501860 197160 504883 197162
rect 501860 197104 504822 197160
rect 504878 197104 504883 197160
rect 501860 197102 504883 197104
rect 504817 197099 504883 197102
rect 502006 196828 502012 196892
rect 502076 196890 502082 196892
rect 503621 196890 503687 196893
rect 502076 196888 503687 196890
rect 502076 196832 503626 196888
rect 503682 196832 503687 196888
rect 502076 196830 503687 196832
rect 502076 196828 502082 196830
rect 503621 196827 503687 196830
rect 501454 196692 501460 196756
rect 501524 196754 501530 196756
rect 502006 196754 502012 196756
rect 501524 196694 502012 196754
rect 501524 196692 501530 196694
rect 502006 196692 502012 196694
rect 502076 196692 502082 196756
rect 78857 196618 78923 196621
rect 78857 196616 82156 196618
rect 78857 196560 78862 196616
rect 78918 196560 82156 196616
rect 78857 196558 82156 196560
rect 78857 196555 78923 196558
rect 501454 196284 501460 196348
rect 501524 196346 501530 196348
rect 504582 196346 504588 196348
rect 501524 196286 504588 196346
rect 501524 196284 501530 196286
rect 504582 196284 504588 196286
rect 504652 196284 504658 196348
rect 501270 196148 501276 196212
rect 501340 196210 501346 196212
rect 503529 196210 503595 196213
rect 501340 196208 503595 196210
rect 501340 196152 503534 196208
rect 503590 196152 503595 196208
rect 501340 196150 503595 196152
rect 501340 196148 501346 196150
rect 503529 196147 503595 196150
rect 501454 195740 501460 195804
rect 501524 195740 501530 195804
rect 501462 195532 501522 195740
rect 501454 195468 501460 195532
rect 501524 195468 501530 195532
rect 82624 195394 82630 195396
rect 82310 195334 82630 195394
rect 82310 195122 82370 195334
rect 82624 195332 82630 195334
rect 82694 195332 82700 195396
rect 82486 195196 82492 195260
rect 82556 195258 82562 195260
rect 82629 195258 82695 195261
rect 82556 195256 82695 195258
rect 82556 195200 82634 195256
rect 82690 195200 82695 195256
rect 82556 195198 82695 195200
rect 82556 195196 82562 195198
rect 82629 195195 82695 195198
rect 82629 195122 82695 195125
rect 82310 195120 82695 195122
rect 82310 195064 82634 195120
rect 82690 195064 82695 195120
rect 82310 195062 82695 195064
rect 82629 195059 82695 195062
rect 82629 194988 82695 194989
rect 82624 194986 82630 194988
rect 82538 194926 82630 194986
rect 82624 194924 82630 194926
rect 82694 194924 82700 194988
rect 82629 194923 82695 194924
rect 82629 194852 82695 194853
rect 82624 194850 82630 194852
rect 82538 194790 82630 194850
rect 82624 194788 82630 194790
rect 82694 194788 82700 194852
rect 82629 194787 82695 194788
rect 77702 194652 77708 194716
rect 77772 194714 77778 194716
rect 82629 194714 82695 194717
rect 77772 194712 82695 194714
rect 77772 194656 82634 194712
rect 82690 194656 82695 194712
rect 77772 194654 82695 194656
rect 77772 194652 77778 194654
rect 82629 194651 82695 194654
rect 501454 194380 501460 194444
rect 501524 194442 501530 194444
rect 503529 194442 503595 194445
rect 501524 194440 503595 194442
rect 501524 194384 503534 194440
rect 503590 194384 503595 194440
rect 501524 194382 503595 194384
rect 501524 194380 501530 194382
rect 503529 194379 503595 194382
rect -960 193898 480 193988
rect 3417 193898 3483 193901
rect -960 193896 3483 193898
rect -960 193840 3422 193896
rect 3478 193840 3483 193896
rect -960 193838 3483 193840
rect -960 193748 480 193838
rect 3417 193835 3483 193838
rect 506974 193836 506980 193900
rect 507044 193898 507050 193900
rect 507342 193898 507348 193900
rect 507044 193838 507348 193898
rect 507044 193836 507050 193838
rect 507342 193836 507348 193838
rect 507412 193836 507418 193900
rect 503529 193626 503595 193629
rect 501860 193624 503595 193626
rect 501860 193568 503534 193624
rect 503590 193568 503595 193624
rect 501860 193566 503595 193568
rect 503529 193563 503595 193566
rect 583520 193476 584960 193716
rect 501454 193156 501460 193220
rect 501524 193218 501530 193220
rect 504582 193218 504588 193220
rect 501524 193158 504588 193218
rect 501524 193156 501530 193158
rect 504582 193156 504588 193158
rect 504652 193156 504658 193220
rect 503478 193082 503484 193084
rect 81525 192266 81591 192269
rect 82310 192266 82370 193052
rect 503118 193022 503484 193082
rect 503118 192541 503178 193022
rect 503478 193020 503484 193022
rect 503548 193020 503554 193084
rect 503478 192884 503484 192948
rect 503548 192946 503554 192948
rect 504030 192946 504036 192948
rect 503548 192886 504036 192946
rect 503548 192884 503554 192886
rect 504030 192884 504036 192886
rect 504100 192884 504106 192948
rect 503069 192536 503178 192541
rect 503069 192480 503074 192536
rect 503130 192480 503178 192536
rect 503069 192478 503178 192480
rect 503069 192475 503135 192478
rect 82486 192340 82492 192404
rect 82556 192340 82562 192404
rect 82624 192340 82630 192404
rect 82694 192340 82700 192404
rect 81525 192264 82370 192266
rect 81525 192208 81530 192264
rect 81586 192208 82370 192264
rect 81525 192206 82370 192208
rect 81525 192203 81591 192206
rect 82494 191996 82554 192340
rect 82486 191932 82492 191996
rect 82556 191932 82562 191996
rect 81525 191858 81591 191861
rect 82632 191858 82692 192340
rect 81525 191856 82692 191858
rect 81525 191800 81530 191856
rect 81586 191800 82692 191856
rect 81525 191798 82692 191800
rect 524413 191858 524479 191861
rect 524597 191858 524663 191861
rect 524413 191856 524663 191858
rect 524413 191800 524418 191856
rect 524474 191800 524602 191856
rect 524658 191800 524663 191856
rect 524413 191798 524663 191800
rect 81525 191795 81591 191798
rect 524413 191795 524479 191798
rect 524597 191795 524663 191798
rect 82624 191388 82630 191452
rect 82694 191388 82700 191452
rect 501270 191388 501276 191452
rect 501340 191450 501346 191452
rect 504582 191450 504588 191452
rect 501340 191390 504588 191450
rect 501340 191388 501346 191390
rect 504582 191388 504588 191390
rect 504652 191388 504658 191452
rect 82632 191314 82692 191388
rect 82126 191254 82692 191314
rect 82126 190770 82186 191254
rect 501270 191252 501276 191316
rect 501340 191314 501346 191316
rect 501638 191314 501644 191316
rect 501340 191254 501644 191314
rect 501340 191252 501346 191254
rect 501638 191252 501644 191254
rect 501708 191252 501714 191316
rect 82486 191116 82492 191180
rect 82556 191178 82562 191180
rect 82629 191178 82695 191181
rect 501454 191178 501460 191180
rect 82556 191176 82695 191178
rect 82556 191120 82634 191176
rect 82690 191120 82695 191176
rect 82556 191118 82695 191120
rect 82556 191116 82562 191118
rect 82629 191115 82695 191118
rect 501278 191118 501460 191178
rect 82486 190844 82492 190908
rect 82556 190906 82562 190908
rect 82629 190906 82695 190909
rect 82556 190904 82695 190906
rect 82556 190848 82634 190904
rect 82690 190848 82695 190904
rect 82556 190846 82695 190848
rect 82556 190844 82562 190846
rect 82629 190843 82695 190846
rect 82537 190770 82603 190773
rect 82126 190768 82603 190770
rect 82126 190712 82542 190768
rect 82598 190712 82603 190768
rect 82126 190710 82603 190712
rect 501278 190770 501338 191118
rect 501454 191116 501460 191118
rect 501524 191116 501530 191180
rect 501638 191116 501644 191180
rect 501708 191178 501714 191180
rect 502190 191178 502196 191180
rect 501708 191118 502196 191178
rect 501708 191116 501714 191118
rect 502190 191116 502196 191118
rect 502260 191116 502266 191180
rect 501454 190980 501460 191044
rect 501524 191042 501530 191044
rect 502006 191042 502012 191044
rect 501524 190982 502012 191042
rect 501524 190980 501530 190982
rect 502006 190980 502012 190982
rect 502076 190980 502082 191044
rect 502006 190844 502012 190908
rect 502076 190906 502082 190908
rect 503478 190906 503484 190908
rect 502076 190846 503484 190906
rect 502076 190844 502082 190846
rect 503478 190844 503484 190846
rect 503548 190844 503554 190908
rect 502190 190770 502196 190772
rect 501278 190710 502196 190770
rect 82537 190707 82603 190710
rect 502190 190708 502196 190710
rect 502260 190708 502266 190772
rect 82302 190436 82308 190500
rect 82372 190498 82378 190500
rect 82537 190498 82603 190501
rect 82372 190496 82603 190498
rect 82372 190440 82542 190496
rect 82598 190440 82603 190496
rect 82372 190438 82603 190440
rect 82372 190436 82378 190438
rect 82537 190435 82603 190438
rect 80145 190362 80211 190365
rect 82624 190362 82630 190364
rect 80145 190360 82630 190362
rect 80145 190304 80150 190360
rect 80206 190304 82630 190360
rect 80145 190302 82630 190304
rect 80145 190299 80211 190302
rect 82624 190300 82630 190302
rect 82694 190300 82700 190364
rect 506841 190090 506907 190093
rect 501860 190088 506907 190090
rect 501860 190032 506846 190088
rect 506902 190032 506907 190088
rect 501860 190030 506907 190032
rect 506841 190027 506907 190030
rect 82494 189277 82554 189788
rect 501270 189756 501276 189820
rect 501340 189818 501346 189820
rect 503069 189818 503135 189821
rect 501340 189816 503135 189818
rect 501340 189760 503074 189816
rect 503130 189760 503135 189816
rect 501340 189758 503135 189760
rect 501340 189756 501346 189758
rect 503069 189755 503135 189758
rect 82494 189272 82603 189277
rect 82494 189216 82542 189272
rect 82598 189216 82603 189272
rect 82494 189214 82603 189216
rect 82537 189211 82603 189214
rect 82486 188668 82492 188732
rect 82556 188730 82562 188732
rect 82629 188730 82695 188733
rect 82556 188728 82695 188730
rect 82556 188672 82634 188728
rect 82690 188672 82695 188728
rect 82556 188670 82695 188672
rect 82556 188668 82562 188670
rect 82629 188667 82695 188670
rect 78254 188396 78260 188460
rect 78324 188458 78330 188460
rect 80329 188458 80395 188461
rect 78324 188456 80395 188458
rect 78324 188400 80334 188456
rect 80390 188400 80395 188456
rect 78324 188398 80395 188400
rect 78324 188396 78330 188398
rect 80329 188395 80395 188398
rect 82486 187308 82492 187372
rect 82556 187370 82562 187372
rect 82629 187370 82695 187373
rect 82556 187368 82695 187370
rect 82556 187312 82634 187368
rect 82690 187312 82695 187368
rect 82556 187310 82695 187312
rect 82556 187308 82562 187310
rect 82629 187307 82695 187310
rect 82629 187100 82695 187101
rect 82624 187098 82630 187100
rect 82538 187038 82630 187098
rect 82624 187036 82630 187038
rect 82694 187036 82700 187100
rect 82629 187035 82695 187036
rect 82486 186900 82492 186964
rect 82556 186962 82562 186964
rect 82629 186962 82695 186965
rect 82556 186960 82695 186962
rect 82556 186904 82634 186960
rect 82690 186904 82695 186960
rect 82556 186902 82695 186904
rect 82556 186900 82562 186902
rect 82629 186899 82695 186902
rect 502006 186900 502012 186964
rect 502076 186962 502082 186964
rect 503478 186962 503484 186964
rect 502076 186902 503484 186962
rect 502076 186900 502082 186902
rect 503478 186900 503484 186902
rect 503548 186900 503554 186964
rect 503621 186826 503687 186829
rect 504214 186826 504220 186828
rect 503621 186824 504220 186826
rect 503621 186768 503626 186824
rect 503682 186768 504220 186824
rect 503621 186766 504220 186768
rect 503621 186763 503687 186766
rect 504214 186764 504220 186766
rect 504284 186764 504290 186828
rect 503069 186690 503135 186693
rect 503069 186688 503362 186690
rect 503069 186632 503074 186688
rect 503130 186632 503362 186688
rect 503069 186630 503362 186632
rect 503069 186627 503135 186630
rect 503069 186554 503135 186557
rect 501860 186552 503135 186554
rect 501860 186496 503074 186552
rect 503130 186496 503135 186552
rect 501860 186494 503135 186496
rect 503069 186491 503135 186494
rect 502190 186356 502196 186420
rect 502260 186418 502266 186420
rect 503302 186418 503362 186630
rect 502260 186358 503362 186418
rect 502260 186356 502266 186358
rect 80329 186282 80395 186285
rect 80329 186280 82156 186282
rect 80329 186224 80334 186280
rect 80390 186224 82156 186280
rect 80329 186222 82156 186224
rect 80329 186219 80395 186222
rect 501270 186220 501276 186284
rect 501340 186220 501346 186284
rect 77518 184588 77524 184652
rect 77588 184650 77594 184652
rect 78765 184650 78831 184653
rect 77588 184648 78831 184650
rect 77588 184592 78770 184648
rect 78826 184592 78831 184648
rect 77588 184590 78831 184592
rect 77588 184588 77594 184590
rect 78765 184587 78831 184590
rect 501278 184380 501338 186220
rect 503805 185874 503871 185877
rect 504398 185874 504404 185876
rect 503805 185872 504404 185874
rect 503805 185816 503810 185872
rect 503866 185816 504404 185872
rect 503805 185814 504404 185816
rect 503805 185811 503871 185814
rect 504398 185812 504404 185814
rect 504468 185812 504474 185876
rect 501454 184724 501460 184788
rect 501524 184724 501530 184788
rect 501638 184724 501644 184788
rect 501708 184724 501714 184788
rect 501822 184724 501828 184788
rect 501892 184724 501898 184788
rect 502006 184724 502012 184788
rect 502076 184724 502082 184788
rect 501462 184380 501522 184724
rect 501646 184380 501706 184724
rect 501830 184516 501890 184724
rect 502014 184516 502074 184724
rect 501822 184452 501828 184516
rect 501892 184452 501898 184516
rect 502006 184452 502012 184516
rect 502076 184452 502082 184516
rect 501270 184316 501276 184380
rect 501340 184316 501346 184380
rect 501454 184316 501460 184380
rect 501524 184316 501530 184380
rect 501638 184316 501644 184380
rect 501708 184316 501714 184380
rect 502190 183772 502196 183836
rect 502260 183834 502266 183836
rect 504214 183834 504220 183836
rect 502260 183774 504220 183834
rect 502260 183772 502266 183774
rect 504214 183772 504220 183774
rect 504284 183772 504290 183836
rect 502190 183636 502196 183700
rect 502260 183698 502266 183700
rect 503478 183698 503484 183700
rect 502260 183638 503484 183698
rect 502260 183636 502266 183638
rect 503478 183636 503484 183638
rect 503548 183636 503554 183700
rect 502006 183500 502012 183564
rect 502076 183562 502082 183564
rect 503805 183562 503871 183565
rect 502076 183560 503871 183562
rect 502076 183504 503810 183560
rect 503866 183504 503871 183560
rect 502076 183502 503871 183504
rect 502076 183500 502082 183502
rect 503805 183499 503871 183502
rect 532693 183562 532759 183565
rect 532877 183562 532943 183565
rect 532693 183560 532943 183562
rect 532693 183504 532698 183560
rect 532754 183504 532882 183560
rect 532938 183504 532943 183560
rect 532693 183502 532943 183504
rect 532693 183499 532759 183502
rect 532877 183499 532943 183502
rect 504817 183018 504883 183021
rect 501860 183016 504883 183018
rect 501860 182960 504822 183016
rect 504878 182960 504883 183016
rect 501860 182958 504883 182960
rect 504817 182955 504883 182958
rect 78765 182746 78831 182749
rect 78765 182744 82156 182746
rect 78765 182688 78770 182744
rect 78826 182688 82156 182744
rect 78765 182686 82156 182688
rect 78765 182683 78831 182686
rect 501454 182276 501460 182340
rect 501524 182338 501530 182340
rect 502006 182338 502012 182340
rect 501524 182278 502012 182338
rect 501524 182276 501530 182278
rect 502006 182276 502012 182278
rect 502076 182276 502082 182340
rect 502190 182066 502196 182068
rect 501278 182006 502196 182066
rect 501278 181794 501338 182006
rect 502190 182004 502196 182006
rect 502260 182004 502266 182068
rect 501454 181868 501460 181932
rect 501524 181930 501530 181932
rect 502190 181930 502196 181932
rect 501524 181870 502196 181930
rect 501524 181868 501530 181870
rect 502190 181868 502196 181870
rect 502260 181868 502266 181932
rect 579705 181930 579771 181933
rect 583520 181930 584960 182020
rect 579705 181928 584960 181930
rect 579705 181872 579710 181928
rect 579766 181872 584960 181928
rect 579705 181870 584960 181872
rect 579705 181867 579771 181870
rect 501454 181794 501460 181796
rect 501278 181734 501460 181794
rect 501454 181732 501460 181734
rect 501524 181732 501530 181796
rect 583520 181780 584960 181870
rect 82486 181324 82492 181388
rect 82556 181324 82562 181388
rect 82302 181052 82308 181116
rect 82372 181114 82378 181116
rect 82494 181114 82554 181324
rect 82372 181054 82554 181114
rect 82372 181052 82378 181054
rect 507526 181052 507532 181116
rect 507596 181114 507602 181116
rect 514661 181114 514727 181117
rect 507596 181112 514727 181114
rect 507596 181056 514666 181112
rect 514722 181056 514727 181112
rect 507596 181054 514727 181056
rect 507596 181052 507602 181054
rect 514661 181051 514727 181054
rect 521561 181114 521627 181117
rect 579705 181114 579771 181117
rect 521561 181112 524338 181114
rect 521561 181056 521566 181112
rect 521622 181056 524338 181112
rect 521561 181054 524338 181056
rect 521561 181051 521627 181054
rect 524278 180842 524338 181054
rect 547830 181112 579771 181114
rect 547830 181056 579710 181112
rect 579766 181056 579771 181112
rect 547830 181054 579771 181056
rect 533981 180978 534047 180981
rect 524462 180976 534047 180978
rect 524462 180920 533986 180976
rect 534042 180920 534047 180976
rect 524462 180918 534047 180920
rect 524462 180842 524522 180918
rect 533981 180915 534047 180918
rect 535453 180978 535519 180981
rect 535453 180976 543658 180978
rect 535453 180920 535458 180976
rect 535514 180920 543658 180976
rect 535453 180918 543658 180920
rect 535453 180915 535519 180918
rect 524278 180782 524522 180842
rect 543598 180842 543658 180918
rect 547830 180842 547890 181054
rect 579705 181051 579771 181054
rect 543598 180782 547890 180842
rect 503805 180298 503871 180301
rect 503302 180296 503871 180298
rect 503302 180240 503810 180296
rect 503866 180240 503871 180296
rect 503302 180238 503871 180240
rect 502190 180100 502196 180164
rect 502260 180162 502266 180164
rect 503069 180162 503135 180165
rect 502260 180160 503135 180162
rect 502260 180104 503074 180160
rect 503130 180104 503135 180160
rect 502260 180102 503135 180104
rect 502260 180100 502266 180102
rect 503069 180099 503135 180102
rect 77886 179964 77892 180028
rect 77956 180026 77962 180028
rect 80237 180026 80303 180029
rect 77956 180024 80303 180026
rect 77956 179968 80242 180024
rect 80298 179968 80303 180024
rect 77956 179966 80303 179968
rect 77956 179964 77962 179966
rect 80237 179963 80303 179966
rect 501454 179964 501460 180028
rect 501524 180026 501530 180028
rect 503302 180026 503362 180238
rect 503805 180235 503871 180238
rect 503478 180100 503484 180164
rect 503548 180162 503554 180164
rect 503805 180162 503871 180165
rect 503548 180160 503871 180162
rect 503548 180104 503810 180160
rect 503866 180104 503871 180160
rect 503548 180102 503871 180104
rect 503548 180100 503554 180102
rect 503805 180099 503871 180102
rect 501524 179966 503362 180026
rect 501524 179964 501530 179966
rect 80237 179890 80303 179893
rect 87321 179892 87387 179893
rect 88701 179892 88767 179893
rect 82486 179890 82492 179892
rect 80237 179888 82492 179890
rect 80237 179832 80242 179888
rect 80298 179832 82492 179888
rect 80237 179830 82492 179832
rect 80237 179827 80303 179830
rect 82486 179828 82492 179830
rect 82556 179828 82562 179892
rect 87316 179828 87322 179892
rect 87386 179890 87392 179892
rect 88701 179890 88748 179892
rect 87386 179830 87478 179890
rect 88656 179888 88748 179890
rect 88656 179832 88706 179888
rect 88656 179830 88748 179832
rect 87386 179828 87392 179830
rect 88701 179828 88748 179830
rect 88812 179828 88818 179892
rect 87321 179827 87387 179828
rect 88701 179827 88767 179828
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect 503805 179482 503871 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect 501860 179480 503871 179482
rect 501860 179424 503810 179480
rect 503866 179424 503871 179480
rect 501860 179422 503871 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 503805 179419 503871 179422
rect 82494 178668 82554 179180
rect 501270 179148 501276 179212
rect 501340 179148 501346 179212
rect 501278 178938 501338 179148
rect 502190 178938 502196 178940
rect 501278 178878 502196 178938
rect 502190 178876 502196 178878
rect 502260 178876 502266 178940
rect 82486 178604 82492 178668
rect 82556 178604 82562 178668
rect 501270 178468 501276 178532
rect 501340 178530 501346 178532
rect 504582 178530 504588 178532
rect 501340 178470 504588 178530
rect 501340 178468 501346 178470
rect 504582 178468 504588 178470
rect 504652 178468 504658 178532
rect 80145 178394 80211 178397
rect 82486 178394 82492 178396
rect 80145 178392 82492 178394
rect 80145 178336 80150 178392
rect 80206 178336 82492 178392
rect 80145 178334 82492 178336
rect 80145 178331 80211 178334
rect 82486 178332 82492 178334
rect 82556 178332 82562 178396
rect 501454 178394 501460 178396
rect 501278 178334 501460 178394
rect 501278 178122 501338 178334
rect 501454 178332 501460 178334
rect 501524 178332 501530 178396
rect 501454 178196 501460 178260
rect 501524 178258 501530 178260
rect 505829 178258 505895 178261
rect 501524 178256 505895 178258
rect 501524 178200 505834 178256
rect 505890 178200 505895 178256
rect 501524 178198 505895 178200
rect 501524 178196 501530 178198
rect 505829 178195 505895 178198
rect 501454 178122 501460 178124
rect 501278 178062 501460 178122
rect 501454 178060 501460 178062
rect 501524 178060 501530 178124
rect 502006 177244 502012 177308
rect 502076 177306 502082 177308
rect 502076 177246 502258 177306
rect 502076 177244 502082 177246
rect 501454 177108 501460 177172
rect 501524 177170 501530 177172
rect 502006 177170 502012 177172
rect 501524 177110 502012 177170
rect 501524 177108 501530 177110
rect 502006 177108 502012 177110
rect 502076 177108 502082 177172
rect 501454 176972 501460 177036
rect 501524 177034 501530 177036
rect 502198 177034 502258 177246
rect 501524 176974 502258 177034
rect 501524 176972 501530 176974
rect 501830 175946 501890 176188
rect 501830 175886 504466 175946
rect 501270 175748 501276 175812
rect 501340 175810 501346 175812
rect 504214 175810 504220 175812
rect 501340 175750 504220 175810
rect 501340 175748 501346 175750
rect 504214 175748 504220 175750
rect 504284 175748 504290 175812
rect 79961 175674 80027 175677
rect 79961 175672 82156 175674
rect 79961 175616 79966 175672
rect 80022 175616 82156 175672
rect 79961 175614 82156 175616
rect 79961 175611 80027 175614
rect 501270 175612 501276 175676
rect 501340 175612 501346 175676
rect 502006 175674 502012 175676
rect 501830 175614 502012 175674
rect 501278 175266 501338 175612
rect 501830 175402 501890 175614
rect 502006 175612 502012 175614
rect 502076 175612 502082 175676
rect 502006 175476 502012 175540
rect 502076 175538 502082 175540
rect 502190 175538 502196 175540
rect 502076 175478 502196 175538
rect 502076 175476 502082 175478
rect 502190 175476 502196 175478
rect 502260 175476 502266 175540
rect 502190 175402 502196 175404
rect 501830 175342 502196 175402
rect 502190 175340 502196 175342
rect 502260 175340 502266 175404
rect 504406 175266 504466 175886
rect 501278 175206 504466 175266
rect 82624 175130 82630 175132
rect 82494 175070 82630 175130
rect 82302 174524 82308 174588
rect 82372 174524 82378 174588
rect 82310 173770 82370 174524
rect 82494 173908 82554 175070
rect 82624 175068 82630 175070
rect 82694 175068 82700 175132
rect 502190 174042 502196 174044
rect 501278 173982 502196 174042
rect 82486 173844 82492 173908
rect 82556 173844 82562 173908
rect 82624 173770 82630 173772
rect 82310 173710 82630 173770
rect 82624 173708 82630 173710
rect 82694 173708 82700 173772
rect 501278 173226 501338 173982
rect 502190 173980 502196 173982
rect 502260 173980 502266 174044
rect 501638 173300 501644 173364
rect 501708 173362 501714 173364
rect 501708 173302 503362 173362
rect 501708 173300 501714 173302
rect 501638 173226 501644 173228
rect 501278 173166 501644 173226
rect 501638 173164 501644 173166
rect 501708 173164 501714 173228
rect 502190 173028 502196 173092
rect 502260 173090 502266 173092
rect 503069 173090 503135 173093
rect 502260 173088 503135 173090
rect 502260 173032 503074 173088
rect 503130 173032 503135 173088
rect 502260 173030 503135 173032
rect 503302 173090 503362 173302
rect 503621 173226 503687 173229
rect 504214 173226 504220 173228
rect 503621 173224 504220 173226
rect 503621 173168 503626 173224
rect 503682 173168 504220 173224
rect 503621 173166 504220 173168
rect 503621 173163 503687 173166
rect 504214 173164 504220 173166
rect 504284 173164 504290 173228
rect 506974 173164 506980 173228
rect 507044 173226 507050 173228
rect 507342 173226 507348 173228
rect 507044 173166 507348 173226
rect 507044 173164 507050 173166
rect 507342 173164 507348 173166
rect 507412 173164 507418 173228
rect 503621 173090 503687 173093
rect 503302 173088 503687 173090
rect 503302 173032 503626 173088
rect 503682 173032 503687 173088
rect 503302 173030 503687 173032
rect 502260 173028 502266 173030
rect 503069 173027 503135 173030
rect 503621 173027 503687 173030
rect 505001 172682 505067 172685
rect 501860 172680 505067 172682
rect 501860 172624 505006 172680
rect 505062 172624 505067 172680
rect 501860 172622 505067 172624
rect 505001 172619 505067 172622
rect 524413 172546 524479 172549
rect 524597 172546 524663 172549
rect 524413 172544 524663 172546
rect 524413 172488 524418 172544
rect 524474 172488 524602 172544
rect 524658 172488 524663 172544
rect 524413 172486 524663 172488
rect 524413 172483 524479 172486
rect 524597 172483 524663 172486
rect 532693 172546 532759 172549
rect 532877 172546 532943 172549
rect 532693 172544 532943 172546
rect 532693 172488 532698 172544
rect 532754 172488 532882 172544
rect 532938 172488 532943 172544
rect 532693 172486 532943 172488
rect 532693 172483 532759 172486
rect 532877 172483 532943 172486
rect 77886 172348 77892 172412
rect 77956 172410 77962 172412
rect 82624 172410 82630 172412
rect 77956 172350 82630 172410
rect 77956 172348 77962 172350
rect 82624 172348 82630 172350
rect 82694 172348 82700 172412
rect 501270 172348 501276 172412
rect 501340 172410 501346 172412
rect 504582 172410 504588 172412
rect 501340 172350 504588 172410
rect 501340 172348 501346 172350
rect 504582 172348 504588 172350
rect 504652 172348 504658 172412
rect 78673 172138 78739 172141
rect 78673 172136 82156 172138
rect 78673 172080 78678 172136
rect 78734 172080 82156 172136
rect 78673 172078 82156 172080
rect 78673 172075 78739 172078
rect 82486 171804 82492 171868
rect 82556 171804 82562 171868
rect 82494 171596 82554 171804
rect 87321 171596 87387 171597
rect 87597 171596 87663 171597
rect 82486 171532 82492 171596
rect 82556 171532 82562 171596
rect 87316 171532 87322 171596
rect 87386 171594 87392 171596
rect 87386 171534 87478 171594
rect 87597 171592 87644 171596
rect 87708 171594 87714 171596
rect 87597 171536 87602 171592
rect 87386 171532 87392 171534
rect 87597 171532 87644 171536
rect 87708 171534 87754 171594
rect 87708 171532 87714 171534
rect 87321 171531 87387 171532
rect 87597 171531 87663 171532
rect 80145 171458 80211 171461
rect 82624 171458 82630 171460
rect 80145 171456 82630 171458
rect 80145 171400 80150 171456
rect 80206 171400 82630 171456
rect 80145 171398 82630 171400
rect 80145 171395 80211 171398
rect 82624 171396 82630 171398
rect 82694 171396 82700 171460
rect 80237 171186 80303 171189
rect 80237 171184 82692 171186
rect 80237 171128 80242 171184
rect 80298 171128 82692 171184
rect 80237 171126 82692 171128
rect 80237 171123 80303 171126
rect 82632 171052 82692 171126
rect 501822 171124 501828 171188
rect 501892 171186 501898 171188
rect 501892 171126 502258 171186
rect 501892 171124 501898 171126
rect 82624 170988 82630 171052
rect 82694 170988 82700 171052
rect 81525 170778 81591 170781
rect 81525 170776 82692 170778
rect 81525 170720 81530 170776
rect 81586 170720 82692 170776
rect 81525 170718 82692 170720
rect 81525 170715 81591 170718
rect 82118 170642 82124 170644
rect 81942 170582 82124 170642
rect 81942 169826 82002 170582
rect 82118 170580 82124 170582
rect 82188 170580 82194 170644
rect 82632 170508 82692 170718
rect 82486 170506 82492 170508
rect 82310 170446 82492 170506
rect 82310 170234 82370 170446
rect 82486 170444 82492 170446
rect 82556 170444 82562 170508
rect 82624 170444 82630 170508
rect 82694 170444 82700 170508
rect 501638 170444 501644 170508
rect 501708 170506 501714 170508
rect 502006 170506 502012 170508
rect 501708 170446 502012 170506
rect 501708 170444 501714 170446
rect 502006 170444 502012 170446
rect 502076 170444 502082 170508
rect 82629 170234 82695 170237
rect 502198 170236 502258 171126
rect 82310 170232 82695 170234
rect 82310 170176 82634 170232
rect 82690 170176 82695 170232
rect 82310 170174 82695 170176
rect 82629 170171 82695 170174
rect 502190 170172 502196 170236
rect 502260 170172 502266 170236
rect 82486 170036 82492 170100
rect 82556 170098 82562 170100
rect 82629 170098 82695 170101
rect 82556 170096 82695 170098
rect 82556 170040 82634 170096
rect 82690 170040 82695 170096
rect 82556 170038 82695 170040
rect 82556 170036 82562 170038
rect 82629 170035 82695 170038
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 82118 169826 82124 169828
rect 81942 169766 82124 169826
rect 82118 169764 82124 169766
rect 82188 169764 82194 169828
rect 503621 169146 503687 169149
rect 501860 169144 503687 169146
rect 501860 169088 503626 169144
rect 503682 169088 503687 169144
rect 501860 169086 503687 169088
rect 503621 169083 503687 169086
rect 78673 168602 78739 168605
rect 78673 168600 82156 168602
rect 78673 168544 78678 168600
rect 78734 168544 82156 168600
rect 78673 168542 82156 168544
rect 78673 168539 78739 168542
rect 501822 166364 501828 166428
rect 501892 166426 501898 166428
rect 502977 166426 503043 166429
rect 501892 166424 503043 166426
rect 501892 166368 502982 166424
rect 503038 166368 503043 166424
rect 501892 166366 503043 166368
rect 501892 166364 501898 166366
rect 502977 166363 503043 166366
rect 501822 165956 501828 166020
rect 501892 166018 501898 166020
rect 502006 166018 502012 166020
rect 501892 165958 502012 166018
rect 501892 165956 501898 165958
rect 502006 165956 502012 165958
rect 502076 165956 502082 166020
rect 502006 165820 502012 165884
rect 502076 165882 502082 165884
rect 503897 165882 503963 165885
rect 502076 165880 503963 165882
rect 502076 165824 503902 165880
rect 503958 165824 503963 165880
rect 502076 165822 503963 165824
rect 502076 165820 502082 165822
rect 503897 165819 503963 165822
rect 78254 165548 78260 165612
rect 78324 165610 78330 165612
rect 80145 165610 80211 165613
rect 503897 165610 503963 165613
rect 78324 165608 80211 165610
rect 78324 165552 80150 165608
rect 80206 165552 80211 165608
rect 78324 165550 80211 165552
rect 501860 165608 503963 165610
rect 501860 165552 503902 165608
rect 503958 165552 503963 165608
rect 501860 165550 503963 165552
rect 78324 165548 78330 165550
rect 80145 165547 80211 165550
rect 503897 165547 503963 165550
rect 502977 165474 503043 165477
rect 504582 165474 504588 165476
rect 502977 165472 504588 165474
rect 502977 165416 502982 165472
rect 503038 165416 504588 165472
rect 502977 165414 504588 165416
rect 502977 165411 503043 165414
rect 504582 165412 504588 165414
rect 504652 165412 504658 165476
rect -960 165066 480 165156
rect 3417 165066 3483 165069
rect -960 165064 3483 165066
rect -960 165008 3422 165064
rect 3478 165008 3483 165064
rect -960 165006 3483 165008
rect -960 164916 480 165006
rect 3417 165003 3483 165006
rect 78673 165066 78739 165069
rect 502977 165066 503043 165069
rect 503478 165066 503484 165068
rect 78673 165064 82156 165066
rect 78673 165008 78678 165064
rect 78734 165008 82156 165064
rect 78673 165006 82156 165008
rect 502977 165064 503484 165066
rect 502977 165008 502982 165064
rect 503038 165008 503484 165064
rect 502977 165006 503484 165008
rect 78673 165003 78739 165006
rect 502977 165003 503043 165006
rect 503478 165004 503484 165006
rect 503548 165004 503554 165068
rect 503478 164868 503484 164932
rect 503548 164930 503554 164932
rect 504214 164930 504220 164932
rect 503548 164870 504220 164930
rect 503548 164868 503554 164870
rect 504214 164868 504220 164870
rect 504284 164868 504290 164932
rect 506974 164868 506980 164932
rect 507044 164930 507050 164932
rect 507342 164930 507348 164932
rect 507044 164870 507348 164930
rect 507044 164868 507050 164870
rect 507342 164868 507348 164870
rect 507412 164868 507418 164932
rect 501454 163780 501460 163844
rect 501524 163842 501530 163844
rect 502977 163842 503043 163845
rect 501524 163840 503043 163842
rect 501524 163784 502982 163840
rect 503038 163784 503043 163840
rect 501524 163782 503043 163784
rect 501524 163780 501530 163782
rect 502977 163779 503043 163782
rect 501454 163644 501460 163708
rect 501524 163706 501530 163708
rect 503897 163706 503963 163709
rect 501524 163704 503963 163706
rect 501524 163648 503902 163704
rect 503958 163648 503963 163704
rect 501524 163646 503963 163648
rect 501524 163644 501530 163646
rect 503897 163643 503963 163646
rect 501454 162828 501460 162892
rect 501524 162890 501530 162892
rect 502977 162890 503043 162893
rect 501524 162888 503043 162890
rect 501524 162832 502982 162888
rect 503038 162832 503043 162888
rect 501524 162830 503043 162832
rect 501524 162828 501530 162830
rect 502977 162827 503043 162830
rect 501454 162420 501460 162484
rect 501524 162482 501530 162484
rect 502977 162482 503043 162485
rect 501524 162480 503043 162482
rect 501524 162424 502982 162480
rect 503038 162424 503043 162480
rect 501524 162422 503043 162424
rect 501524 162420 501530 162422
rect 502977 162419 503043 162422
rect 501638 162284 501644 162348
rect 501708 162346 501714 162348
rect 502977 162346 503043 162349
rect 501708 162344 503043 162346
rect 501708 162288 502982 162344
rect 503038 162288 503043 162344
rect 501708 162286 503043 162288
rect 501708 162284 501714 162286
rect 502977 162283 503043 162286
rect 81525 162210 81591 162213
rect 82486 162210 82492 162212
rect 81525 162208 82492 162210
rect 81525 162152 81530 162208
rect 81586 162152 82492 162208
rect 81525 162150 82492 162152
rect 81525 162147 81591 162150
rect 82486 162148 82492 162150
rect 82556 162148 82562 162212
rect 502977 162074 503043 162077
rect 501860 162072 503043 162074
rect 501860 162016 502982 162072
rect 503038 162016 503043 162072
rect 501860 162014 503043 162016
rect 502977 162011 503043 162014
rect 501270 161740 501276 161804
rect 501340 161802 501346 161804
rect 503897 161802 503963 161805
rect 501340 161800 503963 161802
rect 501340 161744 503902 161800
rect 503958 161744 503963 161800
rect 501340 161742 503963 161744
rect 501340 161740 501346 161742
rect 503897 161739 503963 161742
rect 78673 161530 78739 161533
rect 78673 161528 82156 161530
rect 78673 161472 78678 161528
rect 78734 161472 82156 161528
rect 78673 161470 82156 161472
rect 78673 161467 78739 161470
rect 501270 161332 501276 161396
rect 501340 161394 501346 161396
rect 504030 161394 504036 161396
rect 501340 161334 504036 161394
rect 501340 161332 501346 161334
rect 504030 161332 504036 161334
rect 504100 161332 504106 161396
rect 81525 160850 81591 160853
rect 82486 160850 82492 160852
rect 81525 160848 82492 160850
rect 81525 160792 81530 160848
rect 81586 160792 82492 160848
rect 81525 160790 82492 160792
rect 81525 160787 81591 160790
rect 82486 160788 82492 160790
rect 82556 160788 82562 160852
rect 501638 160788 501644 160852
rect 501708 160850 501714 160852
rect 502006 160850 502012 160852
rect 501708 160790 502012 160850
rect 501708 160788 501714 160790
rect 502006 160788 502012 160790
rect 502076 160788 502082 160852
rect 77886 159020 77892 159084
rect 77956 159082 77962 159084
rect 82302 159082 82308 159084
rect 77956 159022 82308 159082
rect 77956 159020 77962 159022
rect 82302 159020 82308 159022
rect 82372 159020 82378 159084
rect 501689 158946 501755 158949
rect 501822 158946 501828 158948
rect 501689 158944 501828 158946
rect 501689 158888 501694 158944
rect 501750 158888 501828 158944
rect 501689 158886 501828 158888
rect 501689 158883 501755 158886
rect 501822 158884 501828 158886
rect 501892 158884 501898 158948
rect 502006 158748 502012 158812
rect 502076 158810 502082 158812
rect 504081 158810 504147 158813
rect 502076 158808 504147 158810
rect 502076 158752 504086 158808
rect 504142 158752 504147 158808
rect 502076 158750 504147 158752
rect 502076 158748 502082 158750
rect 504081 158747 504147 158750
rect 504081 158538 504147 158541
rect 501860 158536 504147 158538
rect 501860 158480 504086 158536
rect 504142 158480 504147 158536
rect 501860 158478 504147 158480
rect 504081 158475 504147 158478
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect 504582 158068 504588 158132
rect 504652 158130 504658 158132
rect 507761 158130 507827 158133
rect 504652 158128 507827 158130
rect 504652 158072 507766 158128
rect 507822 158072 507827 158128
rect 504652 158070 507827 158072
rect 504652 158068 504658 158070
rect 507761 158067 507827 158070
rect 82678 157453 82738 157964
rect 501270 157932 501276 157996
rect 501340 157994 501346 157996
rect 504030 157994 504036 157996
rect 501340 157934 504036 157994
rect 501340 157932 501346 157934
rect 504030 157932 504036 157934
rect 504100 157932 504106 157996
rect 82629 157448 82738 157453
rect 501597 157452 501663 157453
rect 501597 157450 501644 157452
rect 82629 157392 82634 157448
rect 82690 157392 82738 157448
rect 82629 157390 82738 157392
rect 501552 157448 501644 157450
rect 501552 157392 501602 157448
rect 501552 157390 501644 157392
rect 82629 157387 82695 157390
rect 501597 157388 501644 157390
rect 501708 157388 501714 157452
rect 503989 157450 504055 157453
rect 504582 157450 504588 157452
rect 503989 157448 504588 157450
rect 503989 157392 503994 157448
rect 504050 157392 504588 157448
rect 503989 157390 504588 157392
rect 501597 157387 501663 157388
rect 503989 157387 504055 157390
rect 504582 157388 504588 157390
rect 504652 157388 504658 157452
rect 81525 157314 81591 157317
rect 82486 157314 82492 157316
rect 81525 157312 82492 157314
rect 81525 157256 81530 157312
rect 81586 157256 82492 157312
rect 81525 157254 82492 157256
rect 81525 157251 81591 157254
rect 82486 157252 82492 157254
rect 82556 157252 82562 157316
rect 82302 156708 82308 156772
rect 82372 156770 82378 156772
rect 82624 156770 82630 156772
rect 82372 156710 82630 156770
rect 82372 156708 82378 156710
rect 82624 156708 82630 156710
rect 82694 156708 82700 156772
rect 501454 156572 501460 156636
rect 501524 156634 501530 156636
rect 501689 156634 501755 156637
rect 501524 156632 501755 156634
rect 501524 156576 501694 156632
rect 501750 156576 501755 156632
rect 501524 156574 501755 156576
rect 501524 156572 501530 156574
rect 501689 156571 501755 156574
rect 503478 155756 503484 155820
rect 503548 155818 503554 155820
rect 504214 155818 504220 155820
rect 503548 155758 504220 155818
rect 503548 155756 503554 155758
rect 504214 155756 504220 155758
rect 504284 155756 504290 155820
rect 502190 155620 502196 155684
rect 502260 155682 502266 155684
rect 503478 155682 503484 155684
rect 502260 155622 503484 155682
rect 502260 155620 502266 155622
rect 503478 155620 503484 155622
rect 503548 155620 503554 155684
rect 501873 155274 501939 155277
rect 502190 155274 502196 155276
rect 501873 155272 502196 155274
rect 501873 155216 501878 155272
rect 501934 155216 502196 155272
rect 501873 155214 502196 155216
rect 501873 155211 501939 155214
rect 502190 155212 502196 155214
rect 502260 155212 502266 155276
rect 506974 155212 506980 155276
rect 507044 155274 507050 155276
rect 507342 155274 507348 155276
rect 507044 155214 507348 155274
rect 507044 155212 507050 155214
rect 507342 155212 507348 155214
rect 507412 155212 507418 155276
rect 504081 155002 504147 155005
rect 501860 155000 504147 155002
rect 501860 154944 504086 155000
rect 504142 154944 504147 155000
rect 501860 154942 504147 154944
rect 504081 154939 504147 154942
rect 501689 154728 501755 154733
rect 501689 154672 501694 154728
rect 501750 154672 501755 154728
rect 501689 154667 501755 154672
rect 79961 154458 80027 154461
rect 79961 154456 82156 154458
rect 79961 154400 79966 154456
rect 80022 154400 82156 154456
rect 79961 154398 82156 154400
rect 79961 154395 80027 154398
rect 501692 153370 501752 154667
rect 501462 153310 501752 153370
rect 501462 153234 501522 153310
rect 501278 153174 501522 153234
rect 501278 152690 501338 153174
rect 505829 152690 505895 152693
rect 501278 152688 505895 152690
rect 501278 152632 505834 152688
rect 505890 152632 505895 152688
rect 501278 152630 505895 152632
rect 505829 152627 505895 152630
rect 501454 152084 501460 152148
rect 501524 152146 501530 152148
rect 505829 152146 505895 152149
rect 501524 152144 505895 152146
rect 501524 152088 505834 152144
rect 505890 152088 505895 152144
rect 501524 152086 505895 152088
rect 501524 152084 501530 152086
rect 505829 152083 505895 152086
rect 501505 151874 501571 151877
rect 505829 151874 505895 151877
rect 501505 151872 505895 151874
rect 501505 151816 501510 151872
rect 501566 151816 505834 151872
rect 505890 151816 505895 151872
rect 501505 151814 505895 151816
rect 501505 151811 501571 151814
rect 505829 151811 505895 151814
rect 78765 150922 78831 150925
rect 501462 150924 501522 151436
rect 78765 150920 82156 150922
rect -960 150786 480 150876
rect 78765 150864 78770 150920
rect 78826 150864 82156 150920
rect 78765 150862 82156 150864
rect 78765 150859 78831 150862
rect 501454 150860 501460 150924
rect 501524 150860 501530 150924
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 80145 149698 80211 149701
rect 82486 149698 82492 149700
rect 80145 149696 82492 149698
rect 80145 149640 80150 149696
rect 80206 149640 82492 149696
rect 80145 149638 82492 149640
rect 80145 149635 80211 149638
rect 82486 149636 82492 149638
rect 82556 149636 82562 149700
rect 501454 148820 501460 148884
rect 501524 148882 501530 148884
rect 502333 148882 502399 148885
rect 501524 148880 502399 148882
rect 501524 148824 502338 148880
rect 502394 148824 502399 148880
rect 501524 148822 502399 148824
rect 501524 148820 501530 148822
rect 502333 148819 502399 148822
rect 501454 148548 501460 148612
rect 501524 148610 501530 148612
rect 507342 148610 507348 148612
rect 501524 148550 507348 148610
rect 501524 148548 501530 148550
rect 507342 148548 507348 148550
rect 507412 148548 507418 148612
rect 503713 147930 503779 147933
rect 501860 147928 503779 147930
rect 501860 147872 503718 147928
rect 503774 147872 503779 147928
rect 501860 147870 503779 147872
rect 503713 147867 503779 147870
rect 504541 147658 504607 147661
rect 504406 147656 504607 147658
rect 504406 147600 504546 147656
rect 504602 147600 504607 147656
rect 504406 147598 504607 147600
rect 501270 147460 501276 147524
rect 501340 147522 501346 147524
rect 502333 147522 502399 147525
rect 501340 147520 502399 147522
rect 501340 147464 502338 147520
rect 502394 147464 502399 147520
rect 501340 147462 502399 147464
rect 501340 147460 501346 147462
rect 502333 147459 502399 147462
rect 504406 147386 504466 147598
rect 504541 147595 504607 147598
rect 507526 147386 507532 147388
rect 82310 146844 82370 147356
rect 504406 147326 507532 147386
rect 507526 147324 507532 147326
rect 507596 147324 507602 147388
rect 501454 147188 501460 147252
rect 501524 147250 501530 147252
rect 502333 147250 502399 147253
rect 501524 147248 502399 147250
rect 501524 147192 502338 147248
rect 502394 147192 502399 147248
rect 501524 147190 502399 147192
rect 501524 147188 501530 147190
rect 502333 147187 502399 147190
rect 502333 146978 502399 146981
rect 503478 146978 503484 146980
rect 502333 146976 503484 146978
rect 502333 146920 502338 146976
rect 502394 146920 503484 146976
rect 502333 146918 503484 146920
rect 502333 146915 502399 146918
rect 503478 146916 503484 146918
rect 503548 146916 503554 146980
rect 82302 146780 82308 146844
rect 82372 146780 82378 146844
rect 583520 146556 584960 146796
rect 504081 146162 504147 146165
rect 501278 146160 504147 146162
rect 501278 146104 504086 146160
rect 504142 146104 504147 146160
rect 501278 146102 504147 146104
rect 501278 145890 501338 146102
rect 504081 146099 504147 146102
rect 501454 145964 501460 146028
rect 501524 146026 501530 146028
rect 504081 146026 504147 146029
rect 501524 146024 504147 146026
rect 501524 145968 504086 146024
rect 504142 145968 504147 146024
rect 501524 145966 504147 145968
rect 501524 145964 501530 145966
rect 504081 145963 504147 145966
rect 501454 145890 501460 145892
rect 501278 145830 501460 145890
rect 501454 145828 501460 145830
rect 501524 145828 501530 145892
rect 504081 145890 504147 145893
rect 507342 145890 507348 145892
rect 504081 145888 507348 145890
rect 504081 145832 504086 145888
rect 504142 145832 507348 145888
rect 504081 145830 507348 145832
rect 504081 145827 504147 145830
rect 507342 145828 507348 145830
rect 507412 145828 507418 145892
rect 506974 145556 506980 145620
rect 507044 145618 507050 145620
rect 507342 145618 507348 145620
rect 507044 145558 507348 145618
rect 507044 145556 507050 145558
rect 507342 145556 507348 145558
rect 507412 145556 507418 145620
rect 82302 144468 82308 144532
rect 82372 144468 82378 144532
rect 80237 144122 80303 144125
rect 81525 144122 81591 144125
rect 82310 144122 82370 144468
rect 504081 144394 504147 144397
rect 501860 144392 504147 144394
rect 501860 144336 504086 144392
rect 504142 144336 504147 144392
rect 501860 144334 504147 144336
rect 504081 144331 504147 144334
rect 80237 144120 81591 144122
rect 80237 144064 80242 144120
rect 80298 144064 81530 144120
rect 81586 144064 81591 144120
rect 80237 144062 81591 144064
rect 80237 144059 80303 144062
rect 81525 144059 81591 144062
rect 81758 144062 82370 144122
rect 81525 143986 81591 143989
rect 81758 143986 81818 144062
rect 81525 143984 81818 143986
rect 81525 143928 81530 143984
rect 81586 143928 81818 143984
rect 81525 143926 81818 143928
rect 81525 143923 81591 143926
rect 503478 143924 503484 143988
rect 503548 143986 503554 143988
rect 504541 143986 504607 143989
rect 503548 143984 504607 143986
rect 503548 143928 504546 143984
rect 504602 143928 504607 143984
rect 503548 143926 504607 143928
rect 503548 143924 503554 143926
rect 504541 143923 504607 143926
rect 80237 143850 80303 143853
rect 507761 143850 507827 143853
rect 80237 143848 82156 143850
rect 80237 143792 80242 143848
rect 80298 143792 82156 143848
rect 80237 143790 82156 143792
rect 505694 143848 507827 143850
rect 505694 143792 507766 143848
rect 507822 143792 507827 143848
rect 505694 143790 507827 143792
rect 80237 143787 80303 143790
rect 504541 143578 504607 143581
rect 501278 143576 504607 143578
rect 501278 143520 504546 143576
rect 504602 143520 504607 143576
rect 501278 143518 504607 143520
rect 501278 143442 501338 143518
rect 504541 143515 504607 143518
rect 504541 143442 504607 143445
rect 501278 143440 504607 143442
rect 501278 143384 504546 143440
rect 504602 143384 504607 143440
rect 501278 143382 504607 143384
rect 505694 143442 505754 143790
rect 507761 143787 507827 143790
rect 505829 143442 505895 143445
rect 505694 143440 505895 143442
rect 505694 143384 505834 143440
rect 505890 143384 505895 143440
rect 505694 143382 505895 143384
rect 504541 143379 504607 143382
rect 505829 143379 505895 143382
rect 80145 143170 80211 143173
rect 82486 143170 82492 143172
rect 80145 143168 82492 143170
rect 80145 143112 80150 143168
rect 80206 143112 82492 143168
rect 80145 143110 82492 143112
rect 80145 143107 80211 143110
rect 82486 143108 82492 143110
rect 82556 143108 82562 143172
rect 80145 141946 80211 141949
rect 82486 141946 82492 141948
rect 80145 141944 82492 141946
rect 80145 141888 80150 141944
rect 80206 141888 82492 141944
rect 80145 141886 82492 141888
rect 80145 141883 80211 141886
rect 82486 141884 82492 141886
rect 82556 141884 82562 141948
rect 504541 140858 504607 140861
rect 501860 140856 504607 140858
rect 501860 140800 504546 140856
rect 504602 140800 504607 140856
rect 501860 140798 504607 140800
rect 504541 140795 504607 140798
rect 501270 140524 501276 140588
rect 501340 140586 501346 140588
rect 501873 140586 501939 140589
rect 501340 140584 501939 140586
rect 501340 140528 501878 140584
rect 501934 140528 501939 140584
rect 501340 140526 501939 140528
rect 501340 140524 501346 140526
rect 501873 140523 501939 140526
rect 501270 140388 501276 140452
rect 501340 140450 501346 140452
rect 501873 140450 501939 140453
rect 501340 140448 501939 140450
rect 501340 140392 501878 140448
rect 501934 140392 501939 140448
rect 501340 140390 501939 140392
rect 501340 140388 501346 140390
rect 501873 140387 501939 140390
rect 80145 140314 80211 140317
rect 80145 140312 82156 140314
rect 80145 140256 80150 140312
rect 80206 140256 82156 140312
rect 80145 140254 82156 140256
rect 80145 140251 80211 140254
rect 501270 140252 501276 140316
rect 501340 140314 501346 140316
rect 501873 140314 501939 140317
rect 501340 140312 501939 140314
rect 501340 140256 501878 140312
rect 501934 140256 501939 140312
rect 501340 140254 501939 140256
rect 501340 140252 501346 140254
rect 501873 140251 501939 140254
rect 501454 140116 501460 140180
rect 501524 140178 501530 140180
rect 501873 140178 501939 140181
rect 501524 140176 501939 140178
rect 501524 140120 501878 140176
rect 501934 140120 501939 140176
rect 501524 140118 501939 140120
rect 501524 140116 501530 140118
rect 501873 140115 501939 140118
rect 501873 140044 501939 140045
rect 501822 140042 501828 140044
rect 501782 139982 501828 140042
rect 501892 140040 501939 140044
rect 501934 139984 501939 140040
rect 501822 139980 501828 139982
rect 501892 139980 501939 139984
rect 501873 139979 501939 139980
rect 501822 139844 501828 139908
rect 501892 139906 501898 139908
rect 505829 139906 505895 139909
rect 501892 139904 505895 139906
rect 501892 139848 505834 139904
rect 505890 139848 505895 139904
rect 501892 139846 505895 139848
rect 501892 139844 501898 139846
rect 505829 139843 505895 139846
rect 506238 139300 506244 139364
rect 506308 139362 506314 139364
rect 506974 139362 506980 139364
rect 506308 139302 506980 139362
rect 506308 139300 506314 139302
rect 506974 139300 506980 139302
rect 507044 139300 507050 139364
rect 501873 138818 501939 138821
rect 503478 138818 503484 138820
rect 501873 138816 503484 138818
rect 501873 138760 501878 138816
rect 501934 138760 503484 138816
rect 501873 138758 503484 138760
rect 501873 138755 501939 138758
rect 503478 138756 503484 138758
rect 503548 138756 503554 138820
rect 501454 138620 501460 138684
rect 501524 138682 501530 138684
rect 501822 138682 501828 138684
rect 501524 138622 501828 138682
rect 501524 138620 501530 138622
rect 501822 138620 501828 138622
rect 501892 138620 501898 138684
rect 503478 138620 503484 138684
rect 503548 138682 503554 138684
rect 504030 138682 504036 138684
rect 503548 138622 504036 138682
rect 503548 138620 503554 138622
rect 504030 138620 504036 138622
rect 504100 138620 504106 138684
rect 501454 138546 501460 138548
rect 501278 138486 501460 138546
rect 501278 138274 501338 138486
rect 501454 138484 501460 138486
rect 501524 138484 501530 138548
rect 501454 138348 501460 138412
rect 501524 138410 501530 138412
rect 502333 138410 502399 138413
rect 501524 138408 502399 138410
rect 501524 138352 502338 138408
rect 502394 138352 502399 138408
rect 501524 138350 502399 138352
rect 501524 138348 501530 138350
rect 502333 138347 502399 138350
rect 502333 138274 502399 138277
rect 501278 138272 502399 138274
rect 501278 138216 502338 138272
rect 502394 138216 502399 138272
rect 501278 138214 502399 138216
rect 502333 138211 502399 138214
rect 502006 137940 502012 138004
rect 502076 137940 502082 138004
rect 501638 137804 501644 137868
rect 501708 137866 501714 137868
rect 501873 137866 501939 137869
rect 501708 137864 501939 137866
rect 501708 137808 501878 137864
rect 501934 137808 501939 137864
rect 501708 137806 501939 137808
rect 501708 137804 501714 137806
rect 501873 137803 501939 137806
rect 502014 137732 502074 137940
rect 502006 137668 502012 137732
rect 502076 137668 502082 137732
rect 80830 137458 80836 137460
rect 80286 137398 80836 137458
rect 80286 136778 80346 137398
rect 80830 137396 80836 137398
rect 80900 137396 80906 137460
rect 82486 137458 82492 137460
rect 81022 137398 82492 137458
rect 80421 137322 80487 137325
rect 80830 137322 80836 137324
rect 80421 137320 80836 137322
rect 80421 137264 80426 137320
rect 80482 137264 80836 137320
rect 80421 137262 80836 137264
rect 80421 137259 80487 137262
rect 80830 137260 80836 137262
rect 80900 137260 80906 137324
rect 80421 137186 80487 137189
rect 81022 137186 81082 137398
rect 82486 137396 82492 137398
rect 82556 137396 82562 137460
rect 502333 137458 502399 137461
rect 502333 137456 502626 137458
rect 502333 137400 502338 137456
rect 502394 137400 502626 137456
rect 502333 137398 502626 137400
rect 502333 137395 502399 137398
rect 82302 137322 82308 137324
rect 80421 137184 81082 137186
rect 80421 137128 80426 137184
rect 80482 137128 81082 137184
rect 80421 137126 81082 137128
rect 81206 137262 82308 137322
rect 80421 137123 80487 137126
rect 80421 136914 80487 136917
rect 81206 136914 81266 137262
rect 82302 137260 82308 137262
rect 82372 137260 82378 137324
rect 502333 137322 502399 137325
rect 501860 137320 502399 137322
rect 501860 137264 502338 137320
rect 502394 137264 502399 137320
rect 501860 137262 502399 137264
rect 502333 137259 502399 137262
rect 501270 136988 501276 137052
rect 501340 137050 501346 137052
rect 501873 137050 501939 137053
rect 501340 137048 501939 137050
rect 501340 136992 501878 137048
rect 501934 136992 501939 137048
rect 501340 136990 501939 136992
rect 501340 136988 501346 136990
rect 501873 136987 501939 136990
rect 80421 136912 81266 136914
rect 80421 136856 80426 136912
rect 80482 136856 81266 136912
rect 80421 136854 81266 136856
rect 80421 136851 80487 136854
rect 80421 136778 80487 136781
rect 80286 136776 80487 136778
rect 80286 136720 80426 136776
rect 80482 136720 80487 136776
rect 80286 136718 80487 136720
rect 80421 136715 80487 136718
rect 80973 136778 81039 136781
rect 80973 136776 82156 136778
rect 80973 136720 80978 136776
rect 81034 136720 82156 136776
rect 80973 136718 82156 136720
rect 80973 136715 81039 136718
rect 501270 136716 501276 136780
rect 501340 136778 501346 136780
rect 501873 136778 501939 136781
rect 501340 136776 501939 136778
rect 501340 136720 501878 136776
rect 501934 136720 501939 136776
rect 501340 136718 501939 136720
rect 501340 136716 501346 136718
rect 501873 136715 501939 136718
rect 501822 136580 501828 136644
rect 501892 136642 501898 136644
rect 502566 136642 502626 137398
rect 503713 137322 503779 137325
rect 504030 137322 504036 137324
rect 503713 137320 504036 137322
rect 503713 137264 503718 137320
rect 503774 137264 504036 137320
rect 503713 137262 504036 137264
rect 503713 137259 503779 137262
rect 504030 137260 504036 137262
rect 504100 137260 504106 137324
rect 501892 136582 502626 136642
rect 501892 136580 501898 136582
rect -960 136370 480 136460
rect 3417 136370 3483 136373
rect -960 136368 3483 136370
rect -960 136312 3422 136368
rect 3478 136312 3483 136368
rect -960 136310 3483 136312
rect -960 136220 480 136310
rect 3417 136307 3483 136310
rect 501454 136308 501460 136372
rect 501524 136370 501530 136372
rect 501689 136370 501755 136373
rect 501524 136368 501755 136370
rect 501524 136312 501694 136368
rect 501750 136312 501755 136368
rect 501524 136310 501755 136312
rect 501524 136308 501530 136310
rect 501689 136307 501755 136310
rect 82302 136036 82308 136100
rect 82372 136098 82378 136100
rect 82486 136098 82492 136100
rect 82372 136038 82492 136098
rect 82372 136036 82378 136038
rect 82486 136036 82492 136038
rect 82556 136036 82562 136100
rect 80421 135962 80487 135965
rect 82302 135962 82308 135964
rect 80421 135960 82308 135962
rect 80421 135904 80426 135960
rect 80482 135904 82308 135960
rect 80421 135902 82308 135904
rect 80421 135899 80487 135902
rect 82302 135900 82308 135902
rect 82372 135900 82378 135964
rect 501454 135084 501460 135148
rect 501524 135084 501530 135148
rect 504030 135084 504036 135148
rect 504100 135146 504106 135148
rect 504100 135086 504282 135146
rect 504100 135084 504106 135086
rect 501462 134876 501522 135084
rect 503713 135010 503779 135013
rect 504030 135010 504036 135012
rect 503713 135008 504036 135010
rect 503713 134952 503718 135008
rect 503774 134952 504036 135008
rect 503713 134950 504036 134952
rect 503713 134947 503779 134950
rect 504030 134948 504036 134950
rect 504100 134948 504106 135012
rect 501454 134812 501460 134876
rect 501524 134812 501530 134876
rect 501638 134812 501644 134876
rect 501708 134874 501714 134876
rect 504222 134874 504282 135086
rect 583520 134874 584960 134964
rect 501708 134814 504282 134874
rect 583342 134814 584960 134874
rect 501708 134812 501714 134814
rect 518942 134134 528570 134194
rect 503713 133922 503779 133925
rect 503713 133920 503914 133922
rect 503713 133864 503718 133920
rect 503774 133864 503914 133920
rect 503713 133862 503914 133864
rect 503713 133859 503779 133862
rect 503713 133786 503779 133789
rect 501860 133784 503779 133786
rect 501860 133728 503718 133784
rect 503774 133728 503779 133784
rect 501860 133726 503779 133728
rect 503713 133723 503779 133726
rect 501270 133452 501276 133516
rect 501340 133514 501346 133516
rect 503854 133514 503914 133862
rect 507342 133860 507348 133924
rect 507412 133922 507418 133924
rect 518942 133922 519002 134134
rect 528510 134058 528570 134134
rect 538262 134134 547890 134194
rect 528510 133998 538138 134058
rect 507412 133862 519002 133922
rect 538078 133922 538138 133998
rect 538262 133922 538322 134134
rect 547830 134058 547890 134134
rect 557582 134134 567210 134194
rect 547830 133998 557458 134058
rect 538078 133862 538322 133922
rect 557398 133922 557458 133998
rect 557582 133922 557642 134134
rect 567150 134058 567210 134134
rect 583342 134058 583402 134814
rect 583520 134724 584960 134814
rect 567150 133998 576778 134058
rect 557398 133862 557642 133922
rect 576718 133922 576778 133998
rect 576902 133998 583402 134058
rect 576902 133922 576962 133998
rect 576718 133862 576962 133922
rect 507412 133860 507418 133862
rect 501340 133454 503914 133514
rect 501340 133452 501346 133454
rect 78765 133242 78831 133245
rect 78765 133240 82156 133242
rect 78765 133184 78770 133240
rect 78826 133184 82156 133240
rect 78765 133182 82156 133184
rect 78765 133179 78831 133182
rect 506238 131956 506244 132020
rect 506308 132018 506314 132020
rect 506381 132018 506447 132021
rect 506308 132016 506447 132018
rect 506308 131960 506386 132016
rect 506442 131960 506447 132016
rect 506308 131958 506447 131960
rect 506308 131956 506314 131958
rect 506381 131955 506447 131958
rect 501270 130868 501276 130932
rect 501340 130930 501346 130932
rect 501340 130870 503546 130930
rect 501340 130868 501346 130870
rect 77518 130460 77524 130524
rect 77588 130522 77594 130524
rect 79593 130522 79659 130525
rect 77588 130520 79659 130522
rect 77588 130464 79598 130520
rect 79654 130464 79659 130520
rect 77588 130462 79659 130464
rect 503486 130522 503546 130870
rect 503713 130658 503779 130661
rect 504030 130658 504036 130660
rect 503713 130656 504036 130658
rect 503713 130600 503718 130656
rect 503774 130600 504036 130656
rect 503713 130598 504036 130600
rect 503713 130595 503779 130598
rect 504030 130596 504036 130598
rect 504100 130596 504106 130660
rect 504030 130522 504036 130524
rect 503486 130462 504036 130522
rect 77588 130460 77594 130462
rect 79593 130459 79659 130462
rect 504030 130460 504036 130462
rect 504100 130460 504106 130524
rect 503621 130250 503687 130253
rect 501860 130248 503687 130250
rect 501860 130192 503626 130248
rect 503682 130192 503687 130248
rect 501860 130190 503687 130192
rect 503621 130187 503687 130190
rect 77937 129706 78003 129709
rect 77937 129704 82156 129706
rect 77937 129648 77942 129704
rect 77998 129648 82156 129704
rect 77937 129646 82156 129648
rect 77937 129643 78003 129646
rect 82486 128964 82492 129028
rect 82556 129026 82562 129028
rect 82629 129026 82695 129029
rect 82556 129024 82695 129026
rect 82556 128968 82634 129024
rect 82690 128968 82695 129024
rect 82556 128966 82695 128968
rect 82556 128964 82562 128966
rect 82629 128963 82695 128966
rect 501646 126173 501706 126684
rect 79869 126170 79935 126173
rect 79869 126168 82156 126170
rect 79869 126112 79874 126168
rect 79930 126112 82156 126168
rect 79869 126110 82156 126112
rect 79869 126107 79935 126110
rect 501270 126108 501276 126172
rect 501340 126108 501346 126172
rect 501597 126168 501706 126173
rect 501597 126112 501602 126168
rect 501658 126112 501706 126168
rect 501597 126110 501706 126112
rect 501278 126034 501338 126108
rect 501597 126107 501663 126110
rect 504030 126034 504036 126036
rect 501278 125974 504036 126034
rect 504030 125972 504036 125974
rect 504100 125972 504106 126036
rect 503478 125156 503484 125220
rect 503548 125218 503554 125220
rect 504030 125218 504036 125220
rect 503548 125158 504036 125218
rect 503548 125156 503554 125158
rect 504030 125156 504036 125158
rect 504100 125156 504106 125220
rect 502190 125020 502196 125084
rect 502260 125082 502266 125084
rect 502260 125022 502442 125082
rect 502260 125020 502266 125022
rect 502057 124946 502123 124949
rect 502190 124946 502196 124948
rect 502057 124944 502196 124946
rect 502057 124888 502062 124944
rect 502118 124888 502196 124944
rect 502057 124886 502196 124888
rect 502057 124883 502123 124886
rect 502190 124884 502196 124886
rect 502260 124884 502266 124948
rect 502382 124674 502442 125022
rect 503478 124884 503484 124948
rect 503548 124946 503554 124948
rect 503621 124946 503687 124949
rect 503548 124944 503687 124946
rect 503548 124888 503626 124944
rect 503682 124888 503687 124944
rect 503548 124886 503687 124888
rect 503548 124884 503554 124886
rect 503621 124883 503687 124886
rect 502609 124674 502675 124677
rect 502382 124672 502675 124674
rect 502382 124616 502614 124672
rect 502670 124616 502675 124672
rect 502382 124614 502675 124616
rect 502609 124611 502675 124614
rect 77886 123932 77892 123996
rect 77956 123994 77962 123996
rect 83774 123994 83780 123996
rect 77956 123934 83780 123994
rect 77956 123932 77962 123934
rect 83774 123932 83780 123934
rect 83844 123932 83850 123996
rect 84326 123932 84332 123996
rect 84396 123994 84402 123996
rect 86718 123994 86724 123996
rect 84396 123934 86724 123994
rect 84396 123932 84402 123934
rect 86718 123932 86724 123934
rect 86788 123932 86794 123996
rect 88374 123932 88380 123996
rect 88444 123994 88450 123996
rect 90766 123994 90772 123996
rect 88444 123934 90772 123994
rect 88444 123932 88450 123934
rect 90766 123932 90772 123934
rect 90836 123932 90842 123996
rect 90950 123932 90956 123996
rect 91020 123994 91026 123996
rect 107694 123994 107700 123996
rect 91020 123934 107700 123994
rect 91020 123932 91026 123934
rect 107694 123932 107700 123934
rect 107764 123932 107770 123996
rect 463550 123932 463556 123996
rect 463620 123994 463626 123996
rect 491886 123994 491892 123996
rect 463620 123934 491892 123994
rect 463620 123932 463626 123934
rect 491886 123932 491892 123934
rect 491956 123932 491962 123996
rect 493542 123932 493548 123996
rect 493612 123994 493618 123996
rect 497958 123994 497964 123996
rect 493612 123934 497964 123994
rect 493612 123932 493618 123934
rect 497958 123932 497964 123934
rect 498028 123932 498034 123996
rect 498326 123932 498332 123996
rect 498396 123994 498402 123996
rect 499062 123994 499068 123996
rect 498396 123934 499068 123994
rect 498396 123932 498402 123934
rect 499062 123932 499068 123934
rect 499132 123932 499138 123996
rect 499614 123932 499620 123996
rect 499684 123994 499690 123996
rect 500718 123994 500724 123996
rect 499684 123934 500724 123994
rect 499684 123932 499690 123934
rect 500718 123932 500724 123934
rect 500788 123932 500794 123996
rect 503713 123994 503779 123997
rect 500910 123992 503779 123994
rect 500910 123936 503718 123992
rect 503774 123936 503779 123992
rect 500910 123934 503779 123936
rect 82997 123858 83063 123861
rect 83365 123858 83431 123861
rect 82997 123856 83431 123858
rect 82997 123800 83002 123856
rect 83058 123800 83370 123856
rect 83426 123800 83431 123856
rect 82997 123798 83431 123800
rect 82997 123795 83063 123798
rect 83365 123795 83431 123798
rect 83549 123858 83615 123861
rect 122782 123858 122788 123860
rect 83549 123856 122788 123858
rect 83549 123800 83554 123856
rect 83610 123800 122788 123856
rect 83549 123798 122788 123800
rect 83549 123795 83615 123798
rect 122782 123796 122788 123798
rect 122852 123796 122858 123860
rect 425462 123796 425468 123860
rect 425532 123858 425538 123860
rect 493174 123858 493180 123860
rect 425532 123798 493180 123858
rect 425532 123796 425538 123798
rect 493174 123796 493180 123798
rect 493244 123796 493250 123860
rect 497222 123796 497228 123860
rect 497292 123858 497298 123860
rect 499430 123858 499436 123860
rect 497292 123798 499436 123858
rect 497292 123796 497298 123798
rect 499430 123796 499436 123798
rect 499500 123796 499506 123860
rect 500910 123858 500970 123934
rect 503713 123931 503779 123934
rect 499622 123798 500970 123858
rect 83089 123722 83155 123725
rect 90950 123722 90956 123724
rect 83089 123720 90956 123722
rect 83089 123664 83094 123720
rect 83150 123664 90956 123720
rect 83089 123662 90956 123664
rect 83089 123659 83155 123662
rect 90950 123660 90956 123662
rect 91020 123660 91026 123724
rect 91134 123660 91140 123724
rect 91204 123722 91210 123724
rect 207054 123722 207060 123724
rect 91204 123662 207060 123722
rect 91204 123660 91210 123662
rect 207054 123660 207060 123662
rect 207124 123660 207130 123724
rect 320030 123660 320036 123724
rect 320100 123722 320106 123724
rect 320100 123662 499360 123722
rect 320100 123660 320106 123662
rect 82077 123586 82143 123589
rect 82670 123586 82676 123588
rect 82077 123584 82676 123586
rect 82077 123528 82082 123584
rect 82138 123528 82676 123584
rect 82077 123526 82676 123528
rect 82077 123523 82143 123526
rect 82670 123524 82676 123526
rect 82740 123524 82746 123588
rect 87454 123524 87460 123588
rect 87524 123586 87530 123588
rect 218094 123586 218100 123588
rect 87524 123526 218100 123586
rect 87524 123524 87530 123526
rect 218094 123524 218100 123526
rect 218164 123524 218170 123588
rect 234102 123524 234108 123588
rect 234172 123586 234178 123588
rect 235206 123586 235212 123588
rect 234172 123526 235212 123586
rect 234172 123524 234178 123526
rect 235206 123524 235212 123526
rect 235276 123524 235282 123588
rect 240174 123524 240180 123588
rect 240244 123586 240250 123588
rect 253054 123586 253060 123588
rect 240244 123526 253060 123586
rect 240244 123524 240250 123526
rect 253054 123524 253060 123526
rect 253124 123524 253130 123588
rect 275870 123524 275876 123588
rect 275940 123586 275946 123588
rect 498510 123586 498516 123588
rect 275940 123526 498516 123586
rect 275940 123524 275946 123526
rect 498510 123524 498516 123526
rect 498580 123524 498586 123588
rect 499300 123586 499360 123662
rect 499430 123660 499436 123724
rect 499500 123722 499506 123724
rect 499622 123722 499682 123798
rect 501270 123796 501276 123860
rect 501340 123858 501346 123860
rect 502149 123858 502215 123861
rect 501340 123856 502215 123858
rect 501340 123800 502154 123856
rect 502210 123800 502215 123856
rect 501340 123798 502215 123800
rect 501340 123796 501346 123798
rect 502149 123795 502215 123798
rect 499500 123662 499682 123722
rect 499500 123660 499506 123662
rect 500902 123660 500908 123724
rect 500972 123722 500978 123724
rect 502149 123722 502215 123725
rect 500972 123720 502215 123722
rect 500972 123664 502154 123720
rect 502210 123664 502215 123720
rect 500972 123662 502215 123664
rect 500972 123660 500978 123662
rect 502149 123659 502215 123662
rect 499798 123586 499804 123588
rect 499300 123526 499804 123586
rect 499798 123524 499804 123526
rect 499868 123524 499874 123588
rect 501597 123586 501663 123589
rect 499990 123584 501663 123586
rect 499990 123528 501602 123584
rect 501658 123528 501663 123584
rect 499990 123526 501663 123528
rect 80145 123450 80211 123453
rect 86166 123450 86172 123452
rect 80145 123448 86172 123450
rect 80145 123392 80150 123448
rect 80206 123392 86172 123448
rect 80145 123390 86172 123392
rect 80145 123387 80211 123390
rect 86166 123388 86172 123390
rect 86236 123388 86242 123452
rect 92606 123388 92612 123452
rect 92676 123450 92682 123452
rect 252502 123450 252508 123452
rect 92676 123390 252508 123450
rect 92676 123388 92682 123390
rect 252502 123388 252508 123390
rect 252572 123388 252578 123452
rect 258022 123388 258028 123452
rect 258092 123450 258098 123452
rect 260046 123450 260052 123452
rect 258092 123390 260052 123450
rect 258092 123388 258098 123390
rect 260046 123388 260052 123390
rect 260116 123388 260122 123452
rect 277342 123450 277348 123452
rect 275878 123390 277348 123450
rect 79593 123314 79659 123317
rect 83641 123314 83707 123317
rect 79593 123312 83707 123314
rect 79593 123256 79598 123312
rect 79654 123256 83646 123312
rect 83702 123256 83707 123312
rect 79593 123254 83707 123256
rect 79593 123251 79659 123254
rect 83641 123251 83707 123254
rect 88558 123252 88564 123316
rect 88628 123314 88634 123316
rect 93710 123314 93716 123316
rect 88628 123254 93716 123314
rect 88628 123252 88634 123254
rect 93710 123252 93716 123254
rect 93780 123252 93786 123316
rect 209814 123252 209820 123316
rect 209884 123314 209890 123316
rect 219198 123314 219204 123316
rect 209884 123254 219204 123314
rect 209884 123252 209890 123254
rect 219198 123252 219204 123254
rect 219268 123252 219274 123316
rect 79961 123178 80027 123181
rect 84694 123178 84700 123180
rect 79961 123176 84700 123178
rect 79961 123120 79966 123176
rect 80022 123120 84700 123176
rect 79961 123118 84700 123120
rect 79961 123115 80027 123118
rect 84694 123116 84700 123118
rect 84764 123116 84770 123180
rect 271638 123116 271644 123180
rect 271708 123178 271714 123180
rect 275878 123178 275938 123390
rect 277342 123388 277348 123390
rect 277412 123388 277418 123452
rect 295190 123388 295196 123452
rect 295260 123450 295266 123452
rect 296662 123450 296668 123452
rect 295260 123390 296668 123450
rect 295260 123388 295266 123390
rect 296662 123388 296668 123390
rect 296732 123388 296738 123452
rect 314510 123388 314516 123452
rect 314580 123450 314586 123452
rect 315982 123450 315988 123452
rect 314580 123390 315988 123450
rect 314580 123388 314586 123390
rect 315982 123388 315988 123390
rect 316052 123388 316058 123452
rect 333830 123388 333836 123452
rect 333900 123450 333906 123452
rect 335302 123450 335308 123452
rect 333900 123390 335308 123450
rect 333900 123388 333906 123390
rect 335302 123388 335308 123390
rect 335372 123388 335378 123452
rect 353150 123388 353156 123452
rect 353220 123450 353226 123452
rect 354622 123450 354628 123452
rect 353220 123390 354628 123450
rect 353220 123388 353226 123390
rect 354622 123388 354628 123390
rect 354692 123388 354698 123452
rect 372470 123388 372476 123452
rect 372540 123450 372546 123452
rect 373942 123450 373948 123452
rect 372540 123390 373948 123450
rect 372540 123388 372546 123390
rect 373942 123388 373948 123390
rect 374012 123388 374018 123452
rect 391790 123388 391796 123452
rect 391860 123450 391866 123452
rect 393262 123450 393268 123452
rect 391860 123390 393268 123450
rect 391860 123388 391866 123390
rect 393262 123388 393268 123390
rect 393332 123388 393338 123452
rect 411110 123388 411116 123452
rect 411180 123450 411186 123452
rect 412582 123450 412588 123452
rect 411180 123390 412588 123450
rect 411180 123388 411186 123390
rect 412582 123388 412588 123390
rect 412652 123388 412658 123452
rect 469254 123450 469260 123452
rect 422158 123390 469260 123450
rect 277526 123252 277532 123316
rect 277596 123314 277602 123316
rect 285622 123314 285628 123316
rect 277596 123254 285628 123314
rect 277596 123252 277602 123254
rect 285622 123252 285628 123254
rect 285692 123252 285698 123316
rect 296846 123252 296852 123316
rect 296916 123314 296922 123316
rect 304942 123314 304948 123316
rect 296916 123254 304948 123314
rect 296916 123252 296922 123254
rect 304942 123252 304948 123254
rect 305012 123252 305018 123316
rect 316166 123252 316172 123316
rect 316236 123314 316242 123316
rect 324262 123314 324268 123316
rect 316236 123254 324268 123314
rect 316236 123252 316242 123254
rect 324262 123252 324268 123254
rect 324332 123252 324338 123316
rect 335486 123252 335492 123316
rect 335556 123314 335562 123316
rect 343582 123314 343588 123316
rect 335556 123254 343588 123314
rect 335556 123252 335562 123254
rect 343582 123252 343588 123254
rect 343652 123252 343658 123316
rect 354806 123252 354812 123316
rect 354876 123314 354882 123316
rect 362902 123314 362908 123316
rect 354876 123254 362908 123314
rect 354876 123252 354882 123254
rect 362902 123252 362908 123254
rect 362972 123252 362978 123316
rect 374126 123252 374132 123316
rect 374196 123314 374202 123316
rect 382222 123314 382228 123316
rect 374196 123254 382228 123314
rect 374196 123252 374202 123254
rect 382222 123252 382228 123254
rect 382292 123252 382298 123316
rect 393446 123252 393452 123316
rect 393516 123314 393522 123316
rect 401542 123314 401548 123316
rect 393516 123254 401548 123314
rect 393516 123252 393522 123254
rect 401542 123252 401548 123254
rect 401612 123252 401618 123316
rect 412766 123252 412772 123316
rect 412836 123314 412842 123316
rect 422158 123314 422218 123390
rect 469254 123388 469260 123390
rect 469324 123388 469330 123452
rect 478638 123388 478644 123452
rect 478708 123450 478714 123452
rect 493358 123450 493364 123452
rect 478708 123390 493364 123450
rect 478708 123388 478714 123390
rect 493358 123388 493364 123390
rect 493428 123388 493434 123452
rect 412836 123254 422218 123314
rect 412836 123252 412842 123254
rect 466310 123252 466316 123316
rect 466380 123314 466386 123316
rect 474038 123314 474044 123316
rect 466380 123254 474044 123314
rect 466380 123252 466386 123254
rect 474038 123252 474044 123254
rect 474108 123252 474114 123316
rect 478270 123252 478276 123316
rect 478340 123314 478346 123316
rect 499990 123314 500050 123526
rect 501597 123523 501663 123526
rect 500534 123388 500540 123452
rect 500604 123450 500610 123452
rect 501597 123450 501663 123453
rect 500604 123448 501663 123450
rect 500604 123392 501602 123448
rect 501658 123392 501663 123448
rect 500604 123390 501663 123392
rect 500604 123388 500610 123390
rect 501597 123387 501663 123390
rect 478340 123254 500050 123314
rect 478340 123252 478346 123254
rect 500718 123252 500724 123316
rect 500788 123252 500794 123316
rect 271708 123118 275938 123178
rect 271708 123116 271714 123118
rect 493174 123116 493180 123180
rect 493244 123178 493250 123180
rect 499430 123178 499436 123180
rect 493244 123118 499436 123178
rect 493244 123116 493250 123118
rect 499430 123116 499436 123118
rect 499500 123116 499506 123180
rect 499798 123116 499804 123180
rect 499868 123178 499874 123180
rect 500726 123178 500786 123252
rect 499868 123118 500786 123178
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 499868 123116 499874 123118
rect 77518 122980 77524 123044
rect 77588 123042 77594 123044
rect 86902 123042 86908 123044
rect 77588 122982 86908 123042
rect 77588 122980 77594 122982
rect 86902 122980 86908 122982
rect 86972 122980 86978 123044
rect 88926 122980 88932 123044
rect 88996 123042 89002 123044
rect 92606 123042 92612 123044
rect 88996 122982 92612 123042
rect 88996 122980 89002 122982
rect 92606 122980 92612 122982
rect 92676 122980 92682 123044
rect 285622 122980 285628 123044
rect 285692 123042 285698 123044
rect 295190 123042 295196 123044
rect 285692 122982 295196 123042
rect 285692 122980 285698 122982
rect 295190 122980 295196 122982
rect 295260 122980 295266 123044
rect 304942 122980 304948 123044
rect 305012 123042 305018 123044
rect 314510 123042 314516 123044
rect 305012 122982 314516 123042
rect 305012 122980 305018 122982
rect 314510 122980 314516 122982
rect 314580 122980 314586 123044
rect 324262 122980 324268 123044
rect 324332 123042 324338 123044
rect 333830 123042 333836 123044
rect 324332 122982 333836 123042
rect 324332 122980 324338 122982
rect 333830 122980 333836 122982
rect 333900 122980 333906 123044
rect 343582 122980 343588 123044
rect 343652 123042 343658 123044
rect 353150 123042 353156 123044
rect 343652 122982 353156 123042
rect 343652 122980 343658 122982
rect 353150 122980 353156 122982
rect 353220 122980 353226 123044
rect 362902 122980 362908 123044
rect 362972 123042 362978 123044
rect 372470 123042 372476 123044
rect 362972 122982 372476 123042
rect 362972 122980 362978 122982
rect 372470 122980 372476 122982
rect 372540 122980 372546 123044
rect 382222 122980 382228 123044
rect 382292 123042 382298 123044
rect 391790 123042 391796 123044
rect 382292 122982 391796 123042
rect 382292 122980 382298 122982
rect 391790 122980 391796 122982
rect 391860 122980 391866 123044
rect 401542 122980 401548 123044
rect 401612 123042 401618 123044
rect 411110 123042 411116 123044
rect 401612 122982 411116 123042
rect 401612 122980 401618 122982
rect 411110 122980 411116 122982
rect 411180 122980 411186 123044
rect 493358 122980 493364 123044
rect 493428 123042 493434 123044
rect 500718 123042 500724 123044
rect 493428 122982 500724 123042
rect 493428 122980 493434 122982
rect 500718 122980 500724 122982
rect 500788 122980 500794 123044
rect 82629 122906 82695 122909
rect 99230 122906 99236 122908
rect 82629 122904 99236 122906
rect 82629 122848 82634 122904
rect 82690 122848 99236 122904
rect 82629 122846 99236 122848
rect 82629 122843 82695 122846
rect 99230 122844 99236 122846
rect 99300 122844 99306 122908
rect 369894 122844 369900 122908
rect 369964 122906 369970 122908
rect 379278 122906 379284 122908
rect 369964 122846 379284 122906
rect 369964 122844 369970 122846
rect 379278 122844 379284 122846
rect 379348 122844 379354 122908
rect 417550 122844 417556 122908
rect 417620 122906 417626 122908
rect 420126 122906 420132 122908
rect 417620 122846 420132 122906
rect 417620 122844 417626 122846
rect 420126 122844 420132 122846
rect 420196 122844 420202 122908
rect 425094 122844 425100 122908
rect 425164 122906 425170 122908
rect 434478 122906 434484 122908
rect 425164 122846 434484 122906
rect 425164 122844 425170 122846
rect 434478 122844 434484 122846
rect 434548 122844 434554 122908
rect 469438 122844 469444 122908
rect 469508 122906 469514 122908
rect 478638 122906 478644 122908
rect 469508 122846 478644 122906
rect 469508 122844 469514 122846
rect 478638 122844 478644 122846
rect 478708 122844 478714 122908
rect 486550 122844 486556 122908
rect 486620 122906 486626 122908
rect 501278 122906 501338 123148
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect 486620 122846 501338 122906
rect 486620 122844 486626 122846
rect 88926 122708 88932 122772
rect 88996 122708 89002 122772
rect 89294 122770 89300 122772
rect 89118 122710 89300 122770
rect 88934 122637 88994 122708
rect 87505 122634 87571 122637
rect 87822 122634 87828 122636
rect 87505 122632 87828 122634
rect 87505 122576 87510 122632
rect 87566 122576 87828 122632
rect 87505 122574 87828 122576
rect 87505 122571 87571 122574
rect 87822 122572 87828 122574
rect 87892 122572 87898 122636
rect 88934 122632 89043 122637
rect 88934 122576 88982 122632
rect 89038 122576 89043 122632
rect 88934 122574 89043 122576
rect 88977 122571 89043 122574
rect 78622 122300 78628 122364
rect 78692 122362 78698 122364
rect 86861 122362 86927 122365
rect 78692 122360 86927 122362
rect 78692 122304 86866 122360
rect 86922 122304 86927 122360
rect 78692 122302 86927 122304
rect 89118 122362 89178 122710
rect 89294 122708 89300 122710
rect 89364 122708 89370 122772
rect 91318 122708 91324 122772
rect 91388 122770 91394 122772
rect 91388 122710 149116 122770
rect 91388 122708 91394 122710
rect 149056 122637 149116 122710
rect 237230 122708 237236 122772
rect 237300 122770 237306 122772
rect 502057 122770 502123 122773
rect 237300 122768 502123 122770
rect 237300 122712 502062 122768
rect 502118 122712 502123 122768
rect 237300 122710 502123 122712
rect 237300 122708 237306 122710
rect 502057 122707 502123 122710
rect 89253 122634 89319 122637
rect 90633 122636 90699 122637
rect 89478 122634 89484 122636
rect 89253 122632 89484 122634
rect 89253 122576 89258 122632
rect 89314 122576 89484 122632
rect 89253 122574 89484 122576
rect 89253 122571 89319 122574
rect 89478 122572 89484 122574
rect 89548 122572 89554 122636
rect 90582 122634 90588 122636
rect 90542 122574 90588 122634
rect 90652 122632 90699 122636
rect 90694 122576 90699 122632
rect 90582 122572 90588 122574
rect 90652 122572 90699 122576
rect 91870 122572 91876 122636
rect 91940 122634 91946 122636
rect 92289 122634 92355 122637
rect 91940 122632 92355 122634
rect 91940 122576 92294 122632
rect 92350 122576 92355 122632
rect 91940 122574 92355 122576
rect 91940 122572 91946 122574
rect 90633 122571 90699 122572
rect 92289 122571 92355 122574
rect 101029 122634 101095 122637
rect 114318 122634 114324 122636
rect 101029 122632 114324 122634
rect 101029 122576 101034 122632
rect 101090 122576 114324 122632
rect 101029 122574 114324 122576
rect 101029 122571 101095 122574
rect 114318 122572 114324 122574
rect 114388 122572 114394 122636
rect 114686 122572 114692 122636
rect 114756 122634 114762 122636
rect 124213 122634 124279 122637
rect 114756 122632 124279 122634
rect 114756 122576 124218 122632
rect 124274 122576 124279 122632
rect 114756 122574 124279 122576
rect 114756 122572 114762 122574
rect 124213 122571 124279 122574
rect 133781 122634 133847 122637
rect 143533 122634 143599 122637
rect 133781 122632 143599 122634
rect 133781 122576 133786 122632
rect 133842 122576 143538 122632
rect 143594 122576 143599 122632
rect 133781 122574 143599 122576
rect 133781 122571 133847 122574
rect 143533 122571 143599 122574
rect 149053 122632 149119 122637
rect 149053 122576 149058 122632
rect 149114 122576 149119 122632
rect 149053 122571 149119 122576
rect 153101 122634 153167 122637
rect 172462 122634 172468 122636
rect 153101 122632 172468 122634
rect 153101 122576 153106 122632
rect 153162 122576 172468 122632
rect 153101 122574 172468 122576
rect 153101 122571 153167 122574
rect 172462 122572 172468 122574
rect 172532 122572 172538 122636
rect 191966 122572 191972 122636
rect 192036 122634 192042 122636
rect 201309 122634 201375 122637
rect 192036 122632 201375 122634
rect 192036 122576 201314 122632
rect 201370 122576 201375 122632
rect 192036 122574 201375 122576
rect 192036 122572 192042 122574
rect 201309 122571 201375 122574
rect 216581 122634 216647 122637
rect 500125 122634 500191 122637
rect 500309 122636 500375 122637
rect 500309 122634 500356 122636
rect 216581 122632 500191 122634
rect 216581 122576 216586 122632
rect 216642 122576 500130 122632
rect 500186 122576 500191 122632
rect 216581 122574 500191 122576
rect 500264 122632 500356 122634
rect 500264 122576 500314 122632
rect 500264 122574 500356 122576
rect 216581 122571 216647 122574
rect 500125 122571 500191 122574
rect 500309 122572 500356 122574
rect 500420 122572 500426 122636
rect 500493 122634 500559 122637
rect 507710 122634 507716 122636
rect 500493 122632 507716 122634
rect 500493 122576 500498 122632
rect 500554 122576 507716 122632
rect 500493 122574 507716 122576
rect 500309 122571 500375 122572
rect 500493 122571 500559 122574
rect 507710 122572 507716 122574
rect 507780 122572 507786 122636
rect 90030 122436 90036 122500
rect 90100 122498 90106 122500
rect 179413 122498 179479 122501
rect 90100 122496 179479 122498
rect 90100 122440 179418 122496
rect 179474 122440 179479 122496
rect 90100 122438 179479 122440
rect 90100 122436 90106 122438
rect 179413 122435 179479 122438
rect 209681 122498 209747 122501
rect 506606 122498 506612 122500
rect 209681 122496 506612 122498
rect 209681 122440 209686 122496
rect 209742 122440 506612 122496
rect 209681 122438 506612 122440
rect 209681 122435 209747 122438
rect 506606 122436 506612 122438
rect 506676 122436 506682 122500
rect 89294 122362 89300 122364
rect 89118 122302 89300 122362
rect 78692 122300 78698 122302
rect 86861 122299 86927 122302
rect 89294 122300 89300 122302
rect 89364 122300 89370 122364
rect 92790 122300 92796 122364
rect 92860 122362 92866 122364
rect 167085 122362 167151 122365
rect 92860 122360 167151 122362
rect 92860 122304 167090 122360
rect 167146 122304 167151 122360
rect 92860 122302 167151 122304
rect 92860 122300 92866 122302
rect 167085 122299 167151 122302
rect 169661 122362 169727 122365
rect 191782 122362 191788 122364
rect 169661 122360 191788 122362
rect 169661 122304 169666 122360
rect 169722 122304 191788 122360
rect 169661 122302 191788 122304
rect 169661 122299 169727 122302
rect 191782 122300 191788 122302
rect 191852 122300 191858 122364
rect 201401 122362 201467 122365
rect 212257 122362 212323 122365
rect 201401 122360 212323 122362
rect 201401 122304 201406 122360
rect 201462 122304 212262 122360
rect 212318 122304 212323 122360
rect 201401 122302 212323 122304
rect 201401 122299 201467 122302
rect 212257 122299 212323 122302
rect 212441 122362 212507 122365
rect 508078 122362 508084 122364
rect 212441 122360 508084 122362
rect 212441 122304 212446 122360
rect 212502 122304 508084 122360
rect 212441 122302 508084 122304
rect 212441 122299 212507 122302
rect 508078 122300 508084 122302
rect 508148 122300 508154 122364
rect 83825 122228 83891 122229
rect 83774 122226 83780 122228
rect -960 122090 480 122180
rect 83734 122166 83780 122226
rect 83844 122224 83891 122228
rect 83886 122168 83891 122224
rect 83774 122164 83780 122166
rect 83844 122164 83891 122168
rect 84878 122164 84884 122228
rect 84948 122226 84954 122228
rect 95325 122226 95391 122229
rect 84948 122224 95391 122226
rect 84948 122168 95330 122224
rect 95386 122168 95391 122224
rect 84948 122166 95391 122168
rect 84948 122164 84954 122166
rect 83825 122163 83891 122164
rect 95325 122163 95391 122166
rect 114686 122164 114692 122228
rect 114756 122226 114762 122228
rect 124213 122226 124279 122229
rect 114756 122224 124279 122226
rect 114756 122168 124218 122224
rect 124274 122168 124279 122224
rect 114756 122166 124279 122168
rect 114756 122164 114762 122166
rect 124213 122163 124279 122166
rect 133781 122226 133847 122229
rect 143533 122226 143599 122229
rect 133781 122224 143599 122226
rect 133781 122168 133786 122224
rect 133842 122168 143538 122224
rect 143594 122168 143599 122224
rect 133781 122166 143599 122168
rect 133781 122163 133847 122166
rect 143533 122163 143599 122166
rect 153101 122226 153167 122229
rect 162853 122226 162919 122229
rect 153101 122224 162919 122226
rect 153101 122168 153106 122224
rect 153162 122168 162858 122224
rect 162914 122168 162919 122224
rect 153101 122166 162919 122168
rect 153101 122163 153167 122166
rect 162853 122163 162919 122166
rect 172421 122226 172487 122229
rect 172605 122226 172671 122229
rect 172421 122224 172671 122226
rect 172421 122168 172426 122224
rect 172482 122168 172610 122224
rect 172666 122168 172671 122224
rect 172421 122166 172671 122168
rect 172421 122163 172487 122166
rect 172605 122163 172671 122166
rect 182081 122226 182147 122229
rect 182357 122226 182423 122229
rect 182081 122224 182423 122226
rect 182081 122168 182086 122224
rect 182142 122168 182362 122224
rect 182418 122168 182423 122224
rect 182081 122166 182423 122168
rect 182081 122163 182147 122166
rect 182357 122163 182423 122166
rect 191741 122226 191807 122229
rect 230422 122226 230428 122228
rect 191741 122224 230428 122226
rect 191741 122168 191746 122224
rect 191802 122168 230428 122224
rect 191741 122166 230428 122168
rect 191741 122163 191807 122166
rect 230422 122164 230428 122166
rect 230492 122164 230498 122228
rect 240041 122226 240107 122229
rect 240317 122226 240383 122229
rect 240041 122224 240383 122226
rect 240041 122168 240046 122224
rect 240102 122168 240322 122224
rect 240378 122168 240383 122224
rect 240041 122166 240383 122168
rect 240041 122163 240107 122166
rect 240317 122163 240383 122166
rect 241513 122226 241579 122229
rect 249793 122226 249859 122229
rect 241513 122224 249859 122226
rect 241513 122168 241518 122224
rect 241574 122168 249798 122224
rect 249854 122168 249859 122224
rect 241513 122166 249859 122168
rect 241513 122163 241579 122166
rect 249793 122163 249859 122166
rect 259361 122226 259427 122229
rect 269062 122226 269068 122228
rect 259361 122224 269068 122226
rect 259361 122168 259366 122224
rect 259422 122168 269068 122224
rect 259361 122166 269068 122168
rect 259361 122163 259427 122166
rect 269062 122164 269068 122166
rect 269132 122164 269138 122228
rect 278681 122226 278747 122229
rect 288382 122226 288388 122228
rect 278681 122224 288388 122226
rect 278681 122168 278686 122224
rect 278742 122168 288388 122224
rect 278681 122166 288388 122168
rect 278681 122163 278747 122166
rect 288382 122164 288388 122166
rect 288452 122164 288458 122228
rect 298001 122226 298067 122229
rect 299422 122226 299428 122228
rect 298001 122224 299428 122226
rect 298001 122168 298006 122224
rect 298062 122168 299428 122224
rect 298001 122166 299428 122168
rect 298001 122163 298067 122166
rect 299422 122164 299428 122166
rect 299492 122164 299498 122228
rect 299606 122164 299612 122228
rect 299676 122226 299682 122228
rect 318609 122226 318675 122229
rect 299676 122224 318675 122226
rect 299676 122168 318614 122224
rect 318670 122168 318675 122224
rect 299676 122166 318675 122168
rect 299676 122164 299682 122166
rect 318609 122163 318675 122166
rect 318793 122226 318859 122229
rect 327022 122226 327028 122228
rect 318793 122224 327028 122226
rect 318793 122168 318798 122224
rect 318854 122168 327028 122224
rect 318793 122166 327028 122168
rect 318793 122163 318859 122166
rect 327022 122164 327028 122166
rect 327092 122164 327098 122228
rect 336641 122226 336707 122229
rect 346342 122226 346348 122228
rect 336641 122224 346348 122226
rect 336641 122168 336646 122224
rect 336702 122168 346348 122224
rect 336641 122166 346348 122168
rect 336641 122163 336707 122166
rect 346342 122164 346348 122166
rect 346412 122164 346418 122228
rect 355961 122226 356027 122229
rect 365662 122226 365668 122228
rect 355961 122224 365668 122226
rect 355961 122168 355966 122224
rect 356022 122168 365668 122224
rect 355961 122166 365668 122168
rect 355961 122163 356027 122166
rect 365662 122164 365668 122166
rect 365732 122164 365738 122228
rect 375281 122226 375347 122229
rect 376753 122226 376819 122229
rect 375281 122224 376819 122226
rect 375281 122168 375286 122224
rect 375342 122168 376758 122224
rect 376814 122168 376819 122224
rect 375281 122166 376819 122168
rect 375281 122163 375347 122166
rect 376753 122163 376819 122166
rect 386137 122226 386203 122229
rect 404353 122226 404419 122229
rect 386137 122224 404419 122226
rect 386137 122168 386142 122224
rect 386198 122168 404358 122224
rect 404414 122168 404419 122224
rect 386137 122166 404419 122168
rect 386137 122163 386203 122166
rect 404353 122163 404419 122166
rect 413921 122226 413987 122229
rect 415485 122226 415551 122229
rect 413921 122224 415551 122226
rect 413921 122168 413926 122224
rect 413982 122168 415490 122224
rect 415546 122168 415551 122224
rect 413921 122166 415551 122168
rect 413921 122163 413987 122166
rect 415485 122163 415551 122166
rect 424961 122226 425027 122229
rect 426433 122226 426499 122229
rect 424961 122224 426499 122226
rect 424961 122168 424966 122224
rect 425022 122168 426438 122224
rect 426494 122168 426499 122224
rect 424961 122166 426499 122168
rect 424961 122163 425027 122166
rect 426433 122163 426499 122166
rect 434662 122164 434668 122228
rect 434732 122226 434738 122228
rect 444230 122226 444236 122228
rect 434732 122166 444236 122226
rect 434732 122164 434738 122166
rect 444230 122164 444236 122166
rect 444300 122164 444306 122228
rect 478270 122164 478276 122228
rect 478340 122226 478346 122228
rect 478638 122226 478644 122228
rect 478340 122166 478644 122226
rect 478340 122164 478346 122166
rect 478638 122164 478644 122166
rect 478708 122164 478714 122228
rect 491886 122164 491892 122228
rect 491956 122226 491962 122228
rect 495382 122226 495388 122228
rect 491956 122166 495388 122226
rect 491956 122164 491962 122166
rect 495382 122164 495388 122166
rect 495452 122164 495458 122228
rect 497406 122164 497412 122228
rect 497476 122226 497482 122228
rect 502609 122226 502675 122229
rect 497476 122224 502675 122226
rect 497476 122168 502614 122224
rect 502670 122168 502675 122224
rect 497476 122166 502675 122168
rect 497476 122164 497482 122166
rect 502609 122163 502675 122166
rect 3509 122090 3575 122093
rect -960 122088 3575 122090
rect -960 122032 3514 122088
rect 3570 122032 3575 122088
rect -960 122030 3575 122032
rect -960 121940 480 122030
rect 3509 122027 3575 122030
rect 84510 122028 84516 122092
rect 84580 122090 84586 122092
rect 87270 122090 87276 122092
rect 84580 122030 87276 122090
rect 84580 122028 84586 122030
rect 87270 122028 87276 122030
rect 87340 122028 87346 122092
rect 91502 122028 91508 122092
rect 91572 122090 91578 122092
rect 131205 122090 131271 122093
rect 91572 122088 131271 122090
rect 91572 122032 131210 122088
rect 131266 122032 131271 122088
rect 91572 122030 131271 122032
rect 91572 122028 91578 122030
rect 131205 122027 131271 122030
rect 140681 122090 140747 122093
rect 172513 122090 172579 122093
rect 140681 122088 172579 122090
rect 140681 122032 140686 122088
rect 140742 122032 172518 122088
rect 172574 122032 172579 122088
rect 140681 122030 172579 122032
rect 140681 122027 140747 122030
rect 172513 122027 172579 122030
rect 172789 122090 172855 122093
rect 196617 122090 196683 122093
rect 318742 122090 318748 122092
rect 172789 122088 191850 122090
rect 172789 122032 172794 122088
rect 172850 122032 191850 122088
rect 172789 122030 191850 122032
rect 172789 122027 172855 122030
rect 90582 121892 90588 121956
rect 90652 121954 90658 121956
rect 149053 121954 149119 121957
rect 153193 121954 153259 121957
rect 90652 121894 146586 121954
rect 90652 121892 90658 121894
rect 88977 121818 89043 121821
rect 146385 121818 146451 121821
rect 88977 121816 146451 121818
rect 88977 121760 88982 121816
rect 89038 121760 146390 121816
rect 146446 121760 146451 121816
rect 88977 121758 146451 121760
rect 146526 121818 146586 121894
rect 149053 121952 153259 121954
rect 149053 121896 149058 121952
rect 149114 121896 153198 121952
rect 153254 121896 153259 121952
rect 149053 121894 153259 121896
rect 149053 121891 149119 121894
rect 153193 121891 153259 121894
rect 149053 121818 149119 121821
rect 146526 121816 149119 121818
rect 146526 121760 149058 121816
rect 149114 121760 149119 121816
rect 146526 121758 149119 121760
rect 88977 121755 89043 121758
rect 146385 121755 146451 121758
rect 149053 121755 149119 121758
rect 172462 121756 172468 121820
rect 172532 121818 172538 121820
rect 173893 121818 173959 121821
rect 172532 121816 173959 121818
rect 172532 121760 173898 121816
rect 173954 121760 173959 121816
rect 172532 121758 173959 121760
rect 191790 121818 191850 122030
rect 196617 122088 318748 122090
rect 196617 122032 196622 122088
rect 196678 122032 318748 122088
rect 196617 122030 318748 122032
rect 196617 122027 196683 122030
rect 318742 122028 318748 122030
rect 318812 122028 318818 122092
rect 319110 122028 319116 122092
rect 319180 122090 319186 122092
rect 338062 122090 338068 122092
rect 319180 122030 338068 122090
rect 319180 122028 319186 122030
rect 338062 122028 338068 122030
rect 338132 122028 338138 122092
rect 338430 122028 338436 122092
rect 338500 122090 338506 122092
rect 504582 122090 504588 122092
rect 338500 122030 504588 122090
rect 338500 122028 338506 122030
rect 504582 122028 504588 122030
rect 504652 122028 504658 122092
rect 215150 121892 215156 121956
rect 215220 121954 215226 121956
rect 215518 121954 215524 121956
rect 215220 121894 215524 121954
rect 215220 121892 215226 121894
rect 215518 121892 215524 121894
rect 215588 121892 215594 121956
rect 237097 121954 237163 121957
rect 237230 121954 237236 121956
rect 237097 121952 237236 121954
rect 237097 121896 237102 121952
rect 237158 121896 237236 121952
rect 237097 121894 237236 121896
rect 237097 121891 237163 121894
rect 237230 121892 237236 121894
rect 237300 121892 237306 121956
rect 248321 121954 248387 121957
rect 318742 121954 318748 121956
rect 248321 121952 299490 121954
rect 248321 121896 248326 121952
rect 248382 121896 299490 121952
rect 248321 121894 299490 121896
rect 248321 121891 248387 121894
rect 196617 121818 196683 121821
rect 191790 121816 196683 121818
rect 191790 121760 196622 121816
rect 196678 121760 196683 121816
rect 191790 121758 196683 121760
rect 172532 121756 172538 121758
rect 173893 121755 173959 121758
rect 196617 121755 196683 121758
rect 243486 121756 243492 121820
rect 243556 121818 243562 121820
rect 259310 121818 259316 121820
rect 243556 121758 259316 121818
rect 243556 121756 243562 121758
rect 259310 121756 259316 121758
rect 259380 121756 259386 121820
rect 269062 121756 269068 121820
rect 269132 121818 269138 121820
rect 278681 121818 278747 121821
rect 269132 121816 278747 121818
rect 269132 121760 278686 121816
rect 278742 121760 278747 121816
rect 269132 121758 278747 121760
rect 269132 121756 269138 121758
rect 278681 121755 278747 121758
rect 281206 121756 281212 121820
rect 281276 121818 281282 121820
rect 293166 121818 293172 121820
rect 281276 121758 293172 121818
rect 281276 121756 281282 121758
rect 293166 121756 293172 121758
rect 293236 121756 293242 121820
rect 299430 121818 299490 121894
rect 299614 121894 318748 121954
rect 299614 121818 299674 121894
rect 318742 121892 318748 121894
rect 318812 121892 318818 121956
rect 319110 121892 319116 121956
rect 319180 121954 319186 121956
rect 338062 121954 338068 121956
rect 319180 121894 338068 121954
rect 319180 121892 319186 121894
rect 338062 121892 338068 121894
rect 338132 121892 338138 121956
rect 338614 121892 338620 121956
rect 338684 121954 338690 121956
rect 506790 121954 506796 121956
rect 338684 121894 506796 121954
rect 338684 121892 338690 121894
rect 506790 121892 506796 121894
rect 506860 121892 506866 121956
rect 299430 121758 299674 121818
rect 301446 121756 301452 121820
rect 301516 121818 301522 121820
rect 322606 121818 322612 121820
rect 301516 121758 322612 121818
rect 301516 121756 301522 121758
rect 322606 121756 322612 121758
rect 322676 121756 322682 121820
rect 322841 121818 322907 121821
rect 338113 121818 338179 121821
rect 322841 121816 338179 121818
rect 322841 121760 322846 121816
rect 322902 121760 338118 121816
rect 338174 121760 338179 121816
rect 322841 121758 338179 121760
rect 322841 121755 322907 121758
rect 338113 121755 338179 121758
rect 342989 121818 343055 121821
rect 509785 121818 509851 121821
rect 342989 121816 509851 121818
rect 342989 121760 342994 121816
rect 343050 121760 509790 121816
rect 509846 121760 509851 121816
rect 342989 121758 509851 121760
rect 342989 121755 343055 121758
rect 509785 121755 509851 121758
rect 93710 121620 93716 121684
rect 93780 121682 93786 121684
rect 142153 121682 142219 121685
rect 93780 121680 142219 121682
rect 93780 121624 142158 121680
rect 142214 121624 142219 121680
rect 93780 121622 142219 121624
rect 93780 121620 93786 121622
rect 142153 121619 142219 121622
rect 230606 121620 230612 121684
rect 230676 121682 230682 121684
rect 239857 121682 239923 121685
rect 230676 121680 239923 121682
rect 230676 121624 239862 121680
rect 239918 121624 239923 121680
rect 230676 121622 239923 121624
rect 230676 121620 230682 121622
rect 239857 121619 239923 121622
rect 288382 121620 288388 121684
rect 288452 121682 288458 121684
rect 298001 121682 298067 121685
rect 288452 121680 298067 121682
rect 288452 121624 298006 121680
rect 298062 121624 298067 121680
rect 288452 121622 298067 121624
rect 288452 121620 288458 121622
rect 298001 121619 298067 121622
rect 327022 121620 327028 121684
rect 327092 121682 327098 121684
rect 330937 121682 331003 121685
rect 327092 121680 331003 121682
rect 327092 121624 330942 121680
rect 330998 121624 331003 121680
rect 327092 121622 331003 121624
rect 327092 121620 327098 121622
rect 330937 121619 331003 121622
rect 331070 121620 331076 121684
rect 331140 121682 331146 121684
rect 344870 121682 344876 121684
rect 331140 121622 344876 121682
rect 331140 121620 331146 121622
rect 344870 121620 344876 121622
rect 344940 121620 344946 121684
rect 347078 121620 347084 121684
rect 347148 121682 347154 121684
rect 355961 121682 356027 121685
rect 347148 121680 356027 121682
rect 347148 121624 355966 121680
rect 356022 121624 356027 121680
rect 347148 121622 356027 121624
rect 347148 121620 347154 121622
rect 355961 121619 356027 121622
rect 365662 121620 365668 121684
rect 365732 121682 365738 121684
rect 375281 121682 375347 121685
rect 365732 121680 375347 121682
rect 365732 121624 375286 121680
rect 375342 121624 375347 121680
rect 365732 121622 375347 121624
rect 365732 121620 365738 121622
rect 375281 121619 375347 121622
rect 419441 121682 419507 121685
rect 502926 121682 502932 121684
rect 419441 121680 502932 121682
rect 419441 121624 419446 121680
rect 419502 121624 502932 121680
rect 419441 121622 502932 121624
rect 419441 121619 419507 121622
rect 502926 121620 502932 121622
rect 502996 121620 503002 121684
rect 89662 121484 89668 121548
rect 89732 121546 89738 121548
rect 117773 121546 117839 121549
rect 89732 121544 117839 121546
rect 89732 121488 117778 121544
rect 117834 121488 117839 121544
rect 89732 121486 117839 121488
rect 89732 121484 89738 121486
rect 117773 121483 117839 121486
rect 168281 121546 168347 121549
rect 508405 121546 508471 121549
rect 168281 121544 508471 121546
rect 168281 121488 168286 121544
rect 168342 121488 508410 121544
rect 508466 121488 508471 121544
rect 168281 121486 508471 121488
rect 168281 121483 168347 121486
rect 508405 121483 508471 121486
rect 85062 121348 85068 121412
rect 85132 121410 85138 121412
rect 116710 121410 116716 121412
rect 85132 121350 116716 121410
rect 85132 121348 85138 121350
rect 116710 121348 116716 121350
rect 116780 121348 116786 121412
rect 158713 121410 158779 121413
rect 499205 121410 499271 121413
rect 499389 121412 499455 121413
rect 499389 121410 499436 121412
rect 158713 121408 499271 121410
rect 158713 121352 158718 121408
rect 158774 121352 499210 121408
rect 499266 121352 499271 121408
rect 158713 121350 499271 121352
rect 499344 121408 499436 121410
rect 499344 121352 499394 121408
rect 499344 121350 499436 121352
rect 158713 121347 158779 121350
rect 499205 121347 499271 121350
rect 499389 121348 499436 121350
rect 499500 121348 499506 121412
rect 499849 121410 499915 121413
rect 503621 121410 503687 121413
rect 499849 121408 503687 121410
rect 499849 121352 499854 121408
rect 499910 121352 503626 121408
rect 503682 121352 503687 121408
rect 499849 121350 503687 121352
rect 499389 121347 499455 121348
rect 499849 121347 499915 121350
rect 503621 121347 503687 121350
rect 90214 121212 90220 121276
rect 90284 121274 90290 121276
rect 182449 121274 182515 121277
rect 90284 121272 182515 121274
rect 90284 121216 182454 121272
rect 182510 121216 182515 121272
rect 90284 121214 182515 121216
rect 90284 121212 90290 121214
rect 182449 121211 182515 121214
rect 187233 121274 187299 121277
rect 499113 121274 499179 121277
rect 187233 121272 499179 121274
rect 187233 121216 187238 121272
rect 187294 121216 499118 121272
rect 499174 121216 499179 121272
rect 187233 121214 499179 121216
rect 187233 121211 187299 121214
rect 499113 121211 499179 121214
rect 499297 121274 499363 121277
rect 505686 121274 505692 121276
rect 499297 121272 505692 121274
rect 499297 121216 499302 121272
rect 499358 121216 505692 121272
rect 499297 121214 505692 121216
rect 499297 121211 499363 121214
rect 505686 121212 505692 121214
rect 505756 121212 505762 121276
rect 105353 121138 105419 121141
rect 114318 121138 114324 121140
rect 105353 121136 114324 121138
rect 105353 121080 105358 121136
rect 105414 121080 114324 121136
rect 105353 121078 114324 121080
rect 105353 121075 105419 121078
rect 114318 121076 114324 121078
rect 114388 121076 114394 121140
rect 495382 121076 495388 121140
rect 495452 121138 495458 121140
rect 496077 121138 496143 121141
rect 495452 121136 496143 121138
rect 495452 121080 496082 121136
rect 496138 121080 496143 121136
rect 495452 121078 496143 121080
rect 495452 121076 495458 121078
rect 496077 121075 496143 121078
rect 496486 121076 496492 121140
rect 496556 121138 496562 121140
rect 501454 121138 501460 121140
rect 496556 121078 501460 121138
rect 496556 121076 496562 121078
rect 501454 121076 501460 121078
rect 501524 121076 501530 121140
rect 328361 121002 328427 121005
rect 498377 121004 498443 121005
rect 498561 121004 498627 121005
rect 495934 121002 495940 121004
rect 328361 121000 495940 121002
rect 328361 120944 328366 121000
rect 328422 120944 495940 121000
rect 328361 120942 495940 120944
rect 328361 120939 328427 120942
rect 495934 120940 495940 120942
rect 496004 120940 496010 121004
rect 498326 121002 498332 121004
rect 498286 120942 498332 121002
rect 498396 121000 498443 121004
rect 498438 120944 498443 121000
rect 498326 120940 498332 120942
rect 498396 120940 498443 120944
rect 498510 120940 498516 121004
rect 498580 121002 498627 121004
rect 500401 121002 500467 121005
rect 501086 121002 501092 121004
rect 498580 121000 498672 121002
rect 498622 120944 498672 121000
rect 498580 120942 498672 120944
rect 500401 121000 501092 121002
rect 500401 120944 500406 121000
rect 500462 120944 501092 121000
rect 500401 120942 501092 120944
rect 498580 120940 498627 120942
rect 498377 120939 498443 120940
rect 498561 120939 498627 120940
rect 500401 120939 500467 120942
rect 501086 120940 501092 120942
rect 501156 120940 501162 121004
rect 502057 121002 502123 121005
rect 508589 121002 508655 121005
rect 502057 121000 508655 121002
rect 502057 120944 502062 121000
rect 502118 120944 508594 121000
rect 508650 120944 508655 121000
rect 502057 120942 508655 120944
rect 502057 120939 502123 120942
rect 508589 120939 508655 120942
rect 273161 120866 273227 120869
rect 501638 120866 501644 120868
rect 273161 120864 501644 120866
rect 273161 120808 273166 120864
rect 273222 120808 501644 120864
rect 273161 120806 501644 120808
rect 273161 120803 273227 120806
rect 501638 120804 501644 120806
rect 501708 120804 501714 120868
rect 82854 120668 82860 120732
rect 82924 120730 82930 120732
rect 84101 120730 84167 120733
rect 82924 120728 84167 120730
rect 82924 120672 84106 120728
rect 84162 120672 84167 120728
rect 82924 120670 84167 120672
rect 82924 120668 82930 120670
rect 84101 120667 84167 120670
rect 88190 120668 88196 120732
rect 88260 120730 88266 120732
rect 88425 120730 88491 120733
rect 88260 120728 88491 120730
rect 88260 120672 88430 120728
rect 88486 120672 88491 120728
rect 88260 120670 88491 120672
rect 88260 120668 88266 120670
rect 88425 120667 88491 120670
rect 242801 120730 242867 120733
rect 499941 120730 500007 120733
rect 242801 120728 500007 120730
rect 242801 120672 242806 120728
rect 242862 120672 499946 120728
rect 500002 120672 500007 120728
rect 242801 120670 500007 120672
rect 242801 120667 242867 120670
rect 499941 120667 500007 120670
rect 501086 120668 501092 120732
rect 501156 120730 501162 120732
rect 501873 120730 501939 120733
rect 501156 120728 501939 120730
rect 501156 120672 501878 120728
rect 501934 120672 501939 120728
rect 501156 120670 501939 120672
rect 501156 120668 501162 120670
rect 501873 120667 501939 120670
rect 498377 120594 498443 120597
rect 498510 120594 498516 120596
rect 498377 120592 498516 120594
rect 498377 120536 498382 120592
rect 498438 120536 498516 120592
rect 498377 120534 498516 120536
rect 498377 120531 498443 120534
rect 498510 120532 498516 120534
rect 498580 120532 498586 120596
rect 498929 120594 498995 120597
rect 507577 120594 507643 120597
rect 498929 120592 507643 120594
rect 498929 120536 498934 120592
rect 498990 120536 507582 120592
rect 507638 120536 507643 120592
rect 498929 120534 507643 120536
rect 498929 120531 498995 120534
rect 507577 120531 507643 120534
rect 499113 120458 499179 120461
rect 507158 120458 507164 120460
rect 499113 120456 507164 120458
rect 499113 120400 499118 120456
rect 499174 120400 507164 120456
rect 499113 120398 507164 120400
rect 499113 120395 499179 120398
rect 507158 120396 507164 120398
rect 507228 120396 507234 120460
rect 500033 120324 500099 120325
rect 498694 120260 498700 120324
rect 498764 120322 498770 120324
rect 499614 120322 499620 120324
rect 498764 120262 499620 120322
rect 498764 120260 498770 120262
rect 499614 120260 499620 120262
rect 499684 120260 499690 120324
rect 499982 120322 499988 120324
rect 499942 120262 499988 120322
rect 500052 120320 500099 120324
rect 500094 120264 500099 120320
rect 499982 120260 499988 120262
rect 500052 120260 500099 120264
rect 500033 120259 500099 120260
rect 193254 120124 193260 120188
rect 193324 120186 193330 120188
rect 196566 120186 196572 120188
rect 193324 120126 196572 120186
rect 193324 120124 193330 120126
rect 196566 120124 196572 120126
rect 196636 120124 196642 120188
rect 408534 120124 408540 120188
rect 408604 120186 408610 120188
rect 422886 120186 422892 120188
rect 408604 120126 422892 120186
rect 408604 120124 408610 120126
rect 422886 120124 422892 120126
rect 422956 120124 422962 120188
rect 446622 120124 446628 120188
rect 446692 120186 446698 120188
rect 453614 120186 453620 120188
rect 446692 120126 453620 120186
rect 446692 120124 446698 120126
rect 453614 120124 453620 120126
rect 453684 120124 453690 120188
rect 89253 120050 89319 120053
rect 320633 120050 320699 120053
rect 89253 120048 320699 120050
rect 89253 119992 89258 120048
rect 89314 119992 320638 120048
rect 320694 119992 320699 120048
rect 89253 119990 320699 119992
rect 89253 119987 89319 119990
rect 320633 119987 320699 119990
rect 331254 119988 331260 120052
rect 331324 120050 331330 120052
rect 340638 120050 340644 120052
rect 331324 119990 340644 120050
rect 331324 119988 331330 119990
rect 340638 119988 340644 119990
rect 340708 119988 340714 120052
rect 376702 119988 376708 120052
rect 376772 120050 376778 120052
rect 389633 120050 389699 120053
rect 376772 120048 389699 120050
rect 376772 119992 389638 120048
rect 389694 119992 389699 120048
rect 376772 119990 389699 119992
rect 376772 119988 376778 119990
rect 389633 119987 389699 119990
rect 389817 120050 389883 120053
rect 507485 120050 507551 120053
rect 389817 120048 507551 120050
rect 389817 119992 389822 120048
rect 389878 119992 507490 120048
rect 507546 119992 507551 120048
rect 389817 119990 507551 119992
rect 389817 119987 389883 119990
rect 507485 119987 507551 119990
rect 85246 119852 85252 119916
rect 85316 119914 85322 119916
rect 201493 119914 201559 119917
rect 85316 119912 201559 119914
rect 85316 119856 201498 119912
rect 201554 119856 201559 119912
rect 85316 119854 201559 119856
rect 85316 119852 85322 119854
rect 201493 119851 201559 119854
rect 289721 119914 289787 119917
rect 511349 119914 511415 119917
rect 289721 119912 511415 119914
rect 289721 119856 289726 119912
rect 289782 119856 511354 119912
rect 511410 119856 511415 119912
rect 289721 119854 511415 119856
rect 289721 119851 289787 119854
rect 511349 119851 511415 119854
rect 93342 119716 93348 119780
rect 93412 119778 93418 119780
rect 139577 119778 139643 119781
rect 93412 119776 139643 119778
rect 93412 119720 139582 119776
rect 139638 119720 139643 119776
rect 93412 119718 139643 119720
rect 93412 119716 93418 119718
rect 139577 119715 139643 119718
rect 153101 119778 153167 119781
rect 508865 119778 508931 119781
rect 153101 119776 508931 119778
rect 153101 119720 153106 119776
rect 153162 119720 508870 119776
rect 508926 119720 508931 119776
rect 153101 119718 508931 119720
rect 153101 119715 153167 119718
rect 508865 119715 508931 119718
rect 92238 119580 92244 119644
rect 92308 119642 92314 119644
rect 130009 119642 130075 119645
rect 92308 119640 130075 119642
rect 92308 119584 130014 119640
rect 130070 119584 130075 119640
rect 92308 119582 130075 119584
rect 92308 119580 92314 119582
rect 130009 119579 130075 119582
rect 146201 119642 146267 119645
rect 509734 119642 509740 119644
rect 146201 119640 509740 119642
rect 146201 119584 146206 119640
rect 146262 119584 509740 119640
rect 146201 119582 509740 119584
rect 146201 119579 146267 119582
rect 509734 119580 509740 119582
rect 509804 119580 509810 119644
rect 141969 119506 142035 119509
rect 540329 119506 540395 119509
rect 141969 119504 540395 119506
rect 141969 119448 141974 119504
rect 142030 119448 540334 119504
rect 540390 119448 540395 119504
rect 141969 119446 540395 119448
rect 141969 119443 142035 119446
rect 540329 119443 540395 119446
rect 96705 119370 96771 119373
rect 506657 119370 506723 119373
rect 96705 119368 506723 119370
rect 96705 119312 96710 119368
rect 96766 119312 506662 119368
rect 506718 119312 506723 119368
rect 96705 119310 506723 119312
rect 96705 119307 96771 119310
rect 506657 119307 506723 119310
rect 87822 119172 87828 119236
rect 87892 119234 87898 119236
rect 190453 119234 190519 119237
rect 87892 119232 190519 119234
rect 87892 119176 190458 119232
rect 190514 119176 190519 119232
rect 87892 119174 190519 119176
rect 87892 119172 87898 119174
rect 190453 119171 190519 119174
rect 296621 119234 296687 119237
rect 509366 119234 509372 119236
rect 296621 119232 509372 119234
rect 296621 119176 296626 119232
rect 296682 119176 509372 119232
rect 296621 119174 509372 119176
rect 296621 119171 296687 119174
rect 509366 119172 509372 119174
rect 509436 119172 509442 119236
rect 89846 119036 89852 119100
rect 89916 119098 89922 119100
rect 193213 119098 193279 119101
rect 89916 119096 193279 119098
rect 89916 119040 193218 119096
rect 193274 119040 193279 119096
rect 89916 119038 193279 119040
rect 89916 119036 89922 119038
rect 193213 119035 193279 119038
rect 317321 119098 317387 119101
rect 510245 119098 510311 119101
rect 317321 119096 510311 119098
rect 317321 119040 317326 119096
rect 317382 119040 510250 119096
rect 510306 119040 510311 119096
rect 317321 119038 510311 119040
rect 317321 119035 317387 119038
rect 510245 119035 510311 119038
rect 85614 118900 85620 118964
rect 85684 118962 85690 118964
rect 187693 118962 187759 118965
rect 85684 118960 187759 118962
rect 85684 118904 187698 118960
rect 187754 118904 187759 118960
rect 85684 118902 187759 118904
rect 85684 118900 85690 118902
rect 187693 118899 187759 118902
rect 394734 118900 394740 118964
rect 394804 118962 394810 118964
rect 399518 118962 399524 118964
rect 394804 118902 399524 118962
rect 394804 118900 394810 118902
rect 399518 118900 399524 118902
rect 399588 118900 399594 118964
rect 453982 118900 453988 118964
rect 454052 118962 454058 118964
rect 457294 118962 457300 118964
rect 454052 118902 457300 118962
rect 454052 118900 454058 118902
rect 457294 118900 457300 118902
rect 457364 118900 457370 118964
rect 496721 118962 496787 118965
rect 497406 118962 497412 118964
rect 496721 118960 497412 118962
rect 496721 118904 496726 118960
rect 496782 118904 497412 118960
rect 496721 118902 497412 118904
rect 496721 118899 496787 118902
rect 497406 118900 497412 118902
rect 497476 118900 497482 118964
rect 92606 118764 92612 118828
rect 92676 118826 92682 118828
rect 176653 118826 176719 118829
rect 92676 118824 176719 118826
rect 92676 118768 176658 118824
rect 176714 118768 176719 118824
rect 92676 118766 176719 118768
rect 92676 118764 92682 118766
rect 176653 118763 176719 118766
rect 174486 118628 174492 118692
rect 174556 118690 174562 118692
rect 183318 118690 183324 118692
rect 174556 118630 183324 118690
rect 174556 118628 174562 118630
rect 183318 118628 183324 118630
rect 183388 118628 183394 118692
rect 186262 118628 186268 118692
rect 186332 118690 186338 118692
rect 190494 118690 190500 118692
rect 186332 118630 190500 118690
rect 186332 118628 186338 118630
rect 190494 118628 190500 118630
rect 190564 118628 190570 118692
rect 251214 118628 251220 118692
rect 251284 118690 251290 118692
rect 265566 118690 265572 118692
rect 251284 118630 265572 118690
rect 251284 118628 251290 118630
rect 265566 118628 265572 118630
rect 265636 118628 265642 118692
rect 269798 118628 269804 118692
rect 269868 118690 269874 118692
rect 273662 118690 273668 118692
rect 269868 118630 273668 118690
rect 269868 118628 269874 118630
rect 273662 118628 273668 118630
rect 273732 118628 273738 118692
rect 315982 118628 315988 118692
rect 316052 118690 316058 118692
rect 326838 118690 326844 118692
rect 316052 118630 326844 118690
rect 316052 118628 316058 118630
rect 326838 118628 326844 118630
rect 326908 118628 326914 118692
rect 389633 118690 389699 118693
rect 394550 118690 394556 118692
rect 389633 118688 394556 118690
rect 389633 118632 389638 118688
rect 389694 118632 394556 118688
rect 389633 118630 394556 118632
rect 389633 118627 389699 118630
rect 394550 118628 394556 118630
rect 394620 118628 394626 118692
rect 425094 118628 425100 118692
rect 425164 118690 425170 118692
rect 434294 118690 434300 118692
rect 425164 118630 434300 118690
rect 425164 118628 425170 118630
rect 434294 118628 434300 118630
rect 434364 118628 434370 118692
rect 495934 118220 495940 118284
rect 496004 118282 496010 118284
rect 502057 118282 502123 118285
rect 496004 118280 502123 118282
rect 496004 118224 502062 118280
rect 502118 118224 502123 118280
rect 496004 118222 502123 118224
rect 496004 118220 496010 118222
rect 502057 118219 502123 118222
rect 504030 118220 504036 118284
rect 504100 118282 504106 118284
rect 504541 118282 504607 118285
rect 504100 118280 504607 118282
rect 504100 118224 504546 118280
rect 504602 118224 504607 118280
rect 504100 118222 504607 118224
rect 504100 118220 504106 118222
rect 504541 118219 504607 118222
rect 83181 118012 83247 118013
rect 83181 118010 83228 118012
rect 83136 118008 83228 118010
rect 83136 117952 83186 118008
rect 83136 117950 83228 117952
rect 83181 117948 83228 117950
rect 83292 117948 83298 118012
rect 499798 117948 499804 118012
rect 499868 118010 499874 118012
rect 500309 118010 500375 118013
rect 499868 118008 500375 118010
rect 499868 117952 500314 118008
rect 500370 117952 500375 118008
rect 499868 117950 500375 117952
rect 499868 117948 499874 117950
rect 83181 117947 83247 117948
rect 500309 117947 500375 117950
rect 493501 117196 493567 117197
rect 493501 117194 493548 117196
rect 493456 117192 493548 117194
rect 493456 117136 493506 117192
rect 493456 117134 493548 117136
rect 493501 117132 493548 117134
rect 493612 117132 493618 117196
rect 493501 117131 493567 117132
rect 86033 116924 86099 116925
rect 85982 116922 85988 116924
rect 85942 116862 85988 116922
rect 86052 116920 86099 116924
rect 86094 116864 86099 116920
rect 85982 116860 85988 116862
rect 86052 116860 86099 116864
rect 86033 116859 86099 116860
rect 86902 116724 86908 116788
rect 86972 116786 86978 116788
rect 87137 116786 87203 116789
rect 86972 116784 87203 116786
rect 86972 116728 87142 116784
rect 87198 116728 87203 116784
rect 86972 116726 87203 116728
rect 86972 116724 86978 116726
rect 87137 116723 87203 116726
rect 87321 116786 87387 116789
rect 371325 116786 371391 116789
rect 87321 116784 371391 116786
rect 87321 116728 87326 116784
rect 87382 116728 371330 116784
rect 371386 116728 371391 116784
rect 87321 116726 371391 116728
rect 87321 116723 87387 116726
rect 371325 116723 371391 116726
rect 498326 116724 498332 116788
rect 498396 116786 498402 116788
rect 498561 116786 498627 116789
rect 498396 116784 498627 116786
rect 498396 116728 498566 116784
rect 498622 116728 498627 116784
rect 498396 116726 498627 116728
rect 498396 116724 498402 116726
rect 498561 116723 498627 116726
rect 505686 116724 505692 116788
rect 505756 116786 505762 116788
rect 506238 116786 506244 116788
rect 505756 116726 506244 116786
rect 505756 116724 505762 116726
rect 506238 116724 506244 116726
rect 506308 116724 506314 116788
rect 78990 116588 78996 116652
rect 79060 116650 79066 116652
rect 529933 116650 529999 116653
rect 79060 116648 529999 116650
rect 79060 116592 529938 116648
rect 529994 116592 529999 116648
rect 79060 116590 529999 116592
rect 79060 116588 79066 116590
rect 529933 116587 529999 116590
rect 82302 116452 82308 116516
rect 82372 116514 82378 116516
rect 563145 116514 563211 116517
rect 82372 116512 563211 116514
rect 82372 116456 563150 116512
rect 563206 116456 563211 116512
rect 82372 116454 563211 116456
rect 82372 116452 82378 116454
rect 563145 116451 563211 116454
rect 500718 116180 500724 116244
rect 500788 116242 500794 116244
rect 503478 116242 503484 116244
rect 500788 116182 503484 116242
rect 500788 116180 500794 116182
rect 503478 116180 503484 116182
rect 503548 116180 503554 116244
rect 499062 116044 499068 116108
rect 499132 116106 499138 116108
rect 503989 116106 504055 116109
rect 499132 116104 504055 116106
rect 499132 116048 503994 116104
rect 504050 116048 504055 116104
rect 499132 116046 504055 116048
rect 499132 116044 499138 116046
rect 503989 116043 504055 116046
rect 118417 115970 118483 115973
rect 118417 115968 121562 115970
rect 118417 115912 118422 115968
rect 118478 115912 121562 115968
rect 118417 115910 121562 115912
rect 118417 115907 118483 115910
rect 121361 115834 121427 115837
rect 121502 115834 121562 115910
rect 121361 115832 121562 115834
rect 121361 115776 121366 115832
rect 121422 115776 121562 115832
rect 121361 115774 121562 115776
rect 121361 115771 121427 115774
rect 88006 115364 88012 115428
rect 88076 115426 88082 115428
rect 88374 115426 88380 115428
rect 88076 115366 88380 115426
rect 88076 115364 88082 115366
rect 88374 115364 88380 115366
rect 88444 115364 88450 115428
rect 375281 115426 375347 115429
rect 501270 115426 501276 115428
rect 375281 115424 501276 115426
rect 375281 115368 375286 115424
rect 375342 115368 501276 115424
rect 375281 115366 501276 115368
rect 375281 115363 375347 115366
rect 501270 115364 501276 115366
rect 501340 115364 501346 115428
rect 217961 115290 218027 115293
rect 504398 115290 504404 115292
rect 217961 115288 504404 115290
rect 217961 115232 217966 115288
rect 218022 115232 504404 115288
rect 217961 115230 504404 115232
rect 217961 115227 218027 115230
rect 504398 115228 504404 115230
rect 504468 115228 504474 115292
rect 78806 115092 78812 115156
rect 78876 115154 78882 115156
rect 458173 115154 458239 115157
rect 78876 115152 458239 115154
rect 78876 115096 458178 115152
rect 458234 115096 458239 115152
rect 78876 115094 458239 115096
rect 78876 115092 78882 115094
rect 458173 115091 458239 115094
rect 500401 114612 500467 114613
rect 500350 114610 500356 114612
rect 500310 114550 500356 114610
rect 500420 114608 500467 114612
rect 500462 114552 500467 114608
rect 500350 114548 500356 114550
rect 500420 114548 500467 114552
rect 500401 114547 500467 114548
rect 500125 113386 500191 113389
rect 500125 113384 500234 113386
rect 500125 113328 500130 113384
rect 500186 113328 500234 113384
rect 500125 113323 500234 113328
rect 500174 113252 500234 113323
rect 500166 113188 500172 113252
rect 500236 113188 500242 113252
rect 328453 111482 328519 111485
rect 338062 111482 338068 111484
rect 328453 111480 338068 111482
rect 328453 111424 328458 111480
rect 328514 111424 338068 111480
rect 328453 111422 338068 111424
rect 328453 111419 328519 111422
rect 338062 111420 338068 111422
rect 338132 111420 338138 111484
rect 469213 111482 469279 111485
rect 473302 111482 473308 111484
rect 469213 111480 473308 111482
rect 469213 111424 469218 111480
rect 469274 111424 473308 111480
rect 469213 111422 473308 111424
rect 469213 111419 469279 111422
rect 473302 111420 473308 111422
rect 473372 111420 473378 111484
rect 580349 111482 580415 111485
rect 583520 111482 584960 111572
rect 580349 111480 584960 111482
rect 580349 111424 580354 111480
rect 580410 111424 584960 111480
rect 580349 111422 584960 111424
rect 580349 111419 580415 111422
rect 488533 111346 488599 111349
rect 501086 111346 501092 111348
rect 488533 111344 501092 111346
rect 488533 111288 488538 111344
rect 488594 111288 501092 111344
rect 488533 111286 501092 111288
rect 488533 111283 488599 111286
rect 501086 111284 501092 111286
rect 501156 111284 501162 111348
rect 583520 111332 584960 111422
rect 86585 111210 86651 111213
rect 87270 111210 87276 111212
rect 86585 111208 87276 111210
rect 86585 111152 86590 111208
rect 86646 111152 87276 111208
rect 86585 111150 87276 111152
rect 86585 111147 86651 111150
rect 87270 111148 87276 111150
rect 87340 111148 87346 111212
rect 266077 111210 266143 111213
rect 276013 111210 276079 111213
rect 266077 111208 276079 111210
rect 266077 111152 266082 111208
rect 266138 111152 276018 111208
rect 276074 111152 276079 111208
rect 266077 111150 276079 111152
rect 266077 111147 266143 111150
rect 276013 111147 276079 111150
rect 285489 111210 285555 111213
rect 295333 111210 295399 111213
rect 285489 111208 295399 111210
rect 285489 111152 285494 111208
rect 285550 111152 295338 111208
rect 295394 111152 295399 111208
rect 285489 111150 295399 111152
rect 285489 111147 285555 111150
rect 295333 111147 295399 111150
rect 304901 111210 304967 111213
rect 314653 111210 314719 111213
rect 304901 111208 314719 111210
rect 304901 111152 304906 111208
rect 304962 111152 314658 111208
rect 314714 111152 314719 111208
rect 304901 111150 314719 111152
rect 304901 111147 304967 111150
rect 314653 111147 314719 111150
rect 323577 111210 323643 111213
rect 328453 111210 328519 111213
rect 323577 111208 328519 111210
rect 323577 111152 323582 111208
rect 323638 111152 328458 111208
rect 328514 111152 328519 111208
rect 323577 111150 328519 111152
rect 323577 111147 323643 111150
rect 328453 111147 328519 111150
rect 338062 111148 338068 111212
rect 338132 111210 338138 111212
rect 343541 111210 343607 111213
rect 338132 111208 343607 111210
rect 338132 111152 343546 111208
rect 343602 111152 343607 111208
rect 338132 111150 343607 111152
rect 338132 111148 338138 111150
rect 343541 111147 343607 111150
rect 343725 111210 343791 111213
rect 353293 111210 353359 111213
rect 343725 111208 353359 111210
rect 343725 111152 343730 111208
rect 343786 111152 353298 111208
rect 353354 111152 353359 111208
rect 343725 111150 353359 111152
rect 343725 111147 343791 111150
rect 353293 111147 353359 111150
rect 362769 111210 362835 111213
rect 372705 111210 372771 111213
rect 362769 111208 372771 111210
rect 362769 111152 362774 111208
rect 362830 111152 372710 111208
rect 372766 111152 372771 111208
rect 362769 111150 372771 111152
rect 362769 111147 362835 111150
rect 372705 111147 372771 111150
rect 382089 111210 382155 111213
rect 386505 111210 386571 111213
rect 382089 111208 386571 111210
rect 382089 111152 382094 111208
rect 382150 111152 386510 111208
rect 386566 111152 386571 111208
rect 382089 111150 386571 111152
rect 382089 111147 382155 111150
rect 386505 111147 386571 111150
rect 401685 111210 401751 111213
rect 411253 111210 411319 111213
rect 401685 111208 411319 111210
rect 401685 111152 401690 111208
rect 401746 111152 411258 111208
rect 411314 111152 411319 111208
rect 401685 111150 411319 111152
rect 401685 111147 401751 111150
rect 411253 111147 411319 111150
rect 420729 111210 420795 111213
rect 430573 111210 430639 111213
rect 420729 111208 430639 111210
rect 420729 111152 420734 111208
rect 420790 111152 430578 111208
rect 430634 111152 430639 111208
rect 420729 111150 430639 111152
rect 420729 111147 420795 111150
rect 430573 111147 430639 111150
rect 440141 111210 440207 111213
rect 444465 111210 444531 111213
rect 440141 111208 444531 111210
rect 440141 111152 440146 111208
rect 440202 111152 444470 111208
rect 444526 111152 444531 111208
rect 440141 111150 444531 111152
rect 440141 111147 440207 111150
rect 444465 111147 444531 111150
rect 459645 111210 459711 111213
rect 469213 111210 469279 111213
rect 459645 111208 469279 111210
rect 459645 111152 459650 111208
rect 459706 111152 469218 111208
rect 469274 111152 469279 111208
rect 459645 111150 469279 111152
rect 459645 111147 459711 111150
rect 469213 111147 469279 111150
rect 473302 111148 473308 111212
rect 473372 111210 473378 111212
rect 478781 111210 478847 111213
rect 473372 111208 478847 111210
rect 473372 111152 478786 111208
rect 478842 111152 478847 111208
rect 473372 111150 478847 111152
rect 473372 111148 473378 111150
rect 478781 111147 478847 111150
rect 478965 111210 479031 111213
rect 488533 111210 488599 111213
rect 478965 111208 488599 111210
rect 478965 111152 478970 111208
rect 479026 111152 488538 111208
rect 488594 111152 488599 111208
rect 478965 111150 488599 111152
rect 478965 111147 479031 111150
rect 488533 111147 488599 111150
rect 81198 111012 81204 111076
rect 81268 111074 81274 111076
rect 378133 111074 378199 111077
rect 81268 111072 378199 111074
rect 81268 111016 378138 111072
rect 378194 111016 378199 111072
rect 81268 111014 378199 111016
rect 81268 111012 81274 111014
rect 378133 111011 378199 111014
rect 386505 110938 386571 110941
rect 396022 110938 396028 110940
rect 386505 110936 396028 110938
rect 386505 110880 386510 110936
rect 386566 110880 396028 110936
rect 386505 110878 396028 110880
rect 386505 110875 386571 110878
rect 396022 110876 396028 110878
rect 396092 110876 396098 110940
rect 444465 110938 444531 110941
rect 453982 110938 453988 110940
rect 444465 110936 453988 110938
rect 444465 110880 444470 110936
rect 444526 110880 453988 110936
rect 444465 110878 453988 110880
rect 444465 110875 444531 110878
rect 453982 110876 453988 110878
rect 454052 110876 454058 110940
rect 396022 110604 396028 110668
rect 396092 110666 396098 110668
rect 401685 110666 401751 110669
rect 396092 110664 401751 110666
rect 396092 110608 401690 110664
rect 401746 110608 401751 110664
rect 396092 110606 401751 110608
rect 396092 110604 396098 110606
rect 401685 110603 401751 110606
rect 453982 110604 453988 110668
rect 454052 110666 454058 110668
rect 459645 110666 459711 110669
rect 454052 110664 459711 110666
rect 454052 110608 459650 110664
rect 459706 110608 459711 110664
rect 454052 110606 459711 110608
rect 454052 110604 454058 110606
rect 459645 110603 459711 110606
rect 500125 109716 500191 109717
rect 500125 109714 500172 109716
rect 500080 109712 500172 109714
rect 500080 109656 500130 109712
rect 500080 109654 500172 109656
rect 500125 109652 500172 109654
rect 500236 109652 500242 109716
rect 500125 109651 500191 109652
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 84285 106996 84351 106997
rect 82854 106932 82860 106996
rect 82924 106994 82930 106996
rect 83406 106994 83412 106996
rect 82924 106934 83412 106994
rect 82924 106932 82930 106934
rect 83406 106932 83412 106934
rect 83476 106932 83482 106996
rect 84285 106994 84332 106996
rect 84240 106992 84332 106994
rect 84240 106936 84290 106992
rect 84240 106934 84332 106936
rect 84285 106932 84332 106934
rect 84396 106932 84402 106996
rect 86585 106994 86651 106997
rect 86718 106994 86724 106996
rect 86585 106992 86724 106994
rect 86585 106936 86590 106992
rect 86646 106936 86724 106992
rect 86585 106934 86724 106936
rect 84285 106931 84351 106932
rect 86585 106931 86651 106934
rect 86718 106932 86724 106934
rect 86788 106932 86794 106996
rect 498510 106932 498516 106996
rect 498580 106994 498586 106996
rect 499430 106994 499436 106996
rect 498580 106934 499436 106994
rect 498580 106932 498586 106934
rect 499430 106932 499436 106934
rect 499500 106932 499506 106996
rect 86033 106452 86099 106453
rect 85982 106450 85988 106452
rect 85942 106390 85988 106450
rect 86052 106448 86099 106452
rect 86094 106392 86099 106448
rect 85982 106388 85988 106390
rect 86052 106388 86099 106392
rect 86033 106387 86099 106388
rect 83181 106316 83247 106317
rect 83181 106312 83228 106316
rect 83292 106314 83298 106316
rect 88241 106314 88307 106317
rect 88425 106314 88491 106317
rect 83181 106256 83186 106312
rect 83181 106252 83228 106256
rect 83292 106254 83338 106314
rect 88241 106312 88491 106314
rect 88241 106256 88246 106312
rect 88302 106256 88430 106312
rect 88486 106256 88491 106312
rect 88241 106254 88491 106256
rect 83292 106252 83298 106254
rect 83181 106251 83247 106252
rect 88241 106251 88307 106254
rect 88425 106251 88491 106254
rect 272609 106178 272675 106181
rect 272885 106178 272951 106181
rect 272609 106176 272951 106178
rect 272609 106120 272614 106176
rect 272670 106120 272890 106176
rect 272946 106120 272951 106176
rect 272609 106118 272951 106120
rect 272609 106115 272675 106118
rect 272885 106115 272951 106118
rect 504398 105980 504404 106044
rect 504468 106042 504474 106044
rect 504541 106042 504607 106045
rect 504468 106040 504607 106042
rect 504468 105984 504546 106040
rect 504602 105984 504607 106040
rect 504468 105982 504607 105984
rect 504468 105980 504474 105982
rect 504541 105979 504607 105982
rect 87137 105908 87203 105909
rect 85982 105844 85988 105908
rect 86052 105844 86058 105908
rect 87086 105906 87092 105908
rect 87046 105846 87092 105906
rect 87156 105904 87203 105908
rect 87198 105848 87203 105904
rect 87086 105844 87092 105846
rect 87156 105844 87203 105848
rect 85990 105772 86050 105844
rect 87137 105843 87203 105844
rect 85982 105708 85988 105772
rect 86052 105708 86058 105772
rect 83273 104820 83339 104821
rect 83222 104756 83228 104820
rect 83292 104818 83339 104820
rect 83292 104816 83384 104818
rect 83334 104760 83384 104816
rect 83292 104758 83384 104760
rect 83292 104756 83339 104758
rect 500350 104756 500356 104820
rect 500420 104756 500426 104820
rect 83273 104755 83339 104756
rect 500358 104682 500418 104756
rect 500769 104682 500835 104685
rect 500358 104680 500835 104682
rect 500358 104624 500774 104680
rect 500830 104624 500835 104680
rect 500358 104622 500835 104624
rect 500769 104619 500835 104622
rect 498878 104484 498884 104548
rect 498948 104546 498954 104548
rect 499246 104546 499252 104548
rect 498948 104486 499252 104546
rect 498948 104484 498954 104486
rect 499246 104484 499252 104486
rect 499316 104484 499322 104548
rect 496854 102172 496860 102236
rect 496924 102234 496930 102236
rect 497038 102234 497044 102236
rect 496924 102174 497044 102234
rect 496924 102172 496930 102174
rect 497038 102172 497044 102174
rect 497108 102172 497114 102236
rect 88241 101556 88307 101557
rect 88190 101554 88196 101556
rect 88150 101494 88196 101554
rect 88260 101552 88307 101556
rect 88302 101496 88307 101552
rect 88190 101492 88196 101494
rect 88260 101492 88307 101496
rect 88241 101491 88307 101492
rect 13629 101418 13695 101421
rect 505686 101418 505692 101420
rect 13629 101416 505692 101418
rect 13629 101360 13634 101416
rect 13690 101360 505692 101416
rect 13629 101358 505692 101360
rect 13629 101355 13695 101358
rect 505686 101356 505692 101358
rect 505756 101356 505762 101420
rect 583520 99636 584960 99876
rect 84285 98700 84351 98701
rect 84285 98698 84332 98700
rect 84240 98696 84332 98698
rect 84240 98640 84290 98696
rect 84240 98638 84332 98640
rect 84285 98636 84332 98638
rect 84396 98636 84402 98700
rect 504030 98636 504036 98700
rect 504100 98698 504106 98700
rect 504398 98698 504404 98700
rect 504100 98638 504404 98698
rect 504100 98636 504106 98638
rect 504398 98636 504404 98638
rect 504468 98636 504474 98700
rect 84285 98635 84351 98636
rect 82854 97956 82860 98020
rect 82924 98018 82930 98020
rect 83406 98018 83412 98020
rect 82924 97958 83412 98018
rect 82924 97956 82930 97958
rect 83406 97956 83412 97958
rect 83476 97956 83482 98020
rect 289721 97068 289787 97069
rect 289670 97066 289676 97068
rect 289630 97006 289676 97066
rect 289740 97064 289787 97068
rect 289782 97008 289787 97064
rect 289670 97004 289676 97006
rect 289740 97004 289787 97008
rect 289721 97003 289787 97004
rect 500125 96796 500191 96797
rect 500125 96794 500172 96796
rect 500080 96792 500172 96794
rect 500080 96736 500130 96792
rect 500080 96734 500172 96736
rect 500125 96732 500172 96734
rect 500236 96732 500242 96796
rect 504214 96732 504220 96796
rect 504284 96732 504290 96796
rect 500125 96731 500191 96732
rect 289721 96660 289787 96661
rect 289670 96658 289676 96660
rect 289630 96598 289676 96658
rect 289740 96656 289787 96660
rect 289782 96600 289787 96656
rect 289670 96596 289676 96598
rect 289740 96596 289787 96600
rect 289721 96595 289787 96596
rect 88149 96524 88215 96525
rect 504222 96524 504282 96732
rect 88149 96522 88196 96524
rect 88104 96520 88196 96522
rect 88104 96464 88154 96520
rect 88104 96462 88196 96464
rect 88149 96460 88196 96462
rect 88260 96460 88266 96524
rect 504214 96460 504220 96524
rect 504284 96460 504290 96524
rect 88149 96459 88215 96460
rect 87965 96388 88031 96389
rect 87965 96386 88012 96388
rect 87920 96384 88012 96386
rect 87920 96328 87970 96384
rect 87920 96326 88012 96328
rect 87965 96324 88012 96326
rect 88076 96324 88082 96388
rect 87965 96323 88031 96324
rect 83273 95300 83339 95301
rect 83222 95298 83228 95300
rect 83182 95238 83228 95298
rect 83292 95296 83339 95300
rect 83334 95240 83339 95296
rect 83222 95236 83228 95238
rect 83292 95236 83339 95240
rect 83273 95235 83339 95236
rect 499941 95164 500007 95165
rect 499941 95162 499988 95164
rect 499896 95160 499988 95162
rect 499896 95104 499946 95160
rect 499896 95102 499988 95104
rect 499941 95100 499988 95102
rect 500052 95100 500058 95164
rect 499941 95099 500007 95100
rect 88149 94620 88215 94621
rect 88149 94616 88196 94620
rect 88260 94618 88266 94620
rect 88149 94560 88154 94616
rect 88149 94556 88196 94560
rect 88260 94558 88306 94618
rect 88260 94556 88266 94558
rect 88149 94555 88215 94556
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 500585 92852 500651 92853
rect 500534 92788 500540 92852
rect 500604 92850 500651 92852
rect 500604 92848 500696 92850
rect 500646 92792 500696 92848
rect 500604 92790 500696 92792
rect 500604 92788 500651 92790
rect 500585 92787 500651 92788
rect 87965 92716 88031 92717
rect 500677 92716 500743 92717
rect 87965 92712 88012 92716
rect 88076 92714 88082 92716
rect 500677 92714 500724 92716
rect 87965 92656 87970 92712
rect 87965 92652 88012 92656
rect 88076 92654 88122 92714
rect 500632 92712 500724 92714
rect 500632 92656 500682 92712
rect 500632 92654 500724 92656
rect 88076 92652 88082 92654
rect 500677 92652 500724 92654
rect 500788 92652 500794 92716
rect 87965 92651 88031 92652
rect 500677 92651 500743 92652
rect 88006 92380 88012 92444
rect 88076 92380 88082 92444
rect 499430 92442 499436 92444
rect 499254 92382 499436 92442
rect 88014 92036 88074 92380
rect 499254 92308 499314 92382
rect 499430 92380 499436 92382
rect 499500 92380 499506 92444
rect 499246 92244 499252 92308
rect 499316 92244 499322 92308
rect 88006 91972 88012 92036
rect 88076 91972 88082 92036
rect 500585 91764 500651 91765
rect 500534 91762 500540 91764
rect 500494 91702 500540 91762
rect 500604 91760 500651 91764
rect 500646 91704 500651 91760
rect 500534 91700 500540 91702
rect 500604 91700 500651 91704
rect 500585 91699 500651 91700
rect 87638 88300 87644 88364
rect 87708 88362 87714 88364
rect 88190 88362 88196 88364
rect 87708 88302 88196 88362
rect 87708 88300 87714 88302
rect 88190 88300 88196 88302
rect 88260 88300 88266 88364
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 503989 87684 504055 87685
rect 503989 87682 504036 87684
rect 503944 87680 504036 87682
rect 503944 87624 503994 87680
rect 503944 87622 504036 87624
rect 503989 87620 504036 87622
rect 504100 87620 504106 87684
rect 503989 87619 504055 87620
rect 518942 87214 528570 87274
rect 289537 87002 289603 87005
rect 289721 87002 289787 87005
rect 289537 87000 289787 87002
rect 289537 86944 289542 87000
rect 289598 86944 289726 87000
rect 289782 86944 289787 87000
rect 289537 86942 289787 86944
rect 289537 86939 289603 86942
rect 289721 86939 289787 86942
rect 436093 87002 436159 87005
rect 436277 87002 436343 87005
rect 436093 87000 436343 87002
rect 436093 86944 436098 87000
rect 436154 86944 436282 87000
rect 436338 86944 436343 87000
rect 436093 86942 436343 86944
rect 436093 86939 436159 86942
rect 436277 86939 436343 86942
rect 500769 87002 500835 87005
rect 501086 87002 501092 87004
rect 500769 87000 501092 87002
rect 500769 86944 500774 87000
rect 500830 86944 501092 87000
rect 500769 86942 501092 86944
rect 500769 86939 500835 86942
rect 501086 86940 501092 86942
rect 501156 86940 501162 87004
rect 506054 86940 506060 87004
rect 506124 87002 506130 87004
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 557582 87214 567210 87274
rect 528510 87078 538138 87138
rect 506124 86942 519002 87002
rect 538078 87002 538138 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 538078 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 506124 86940 506130 86942
rect 83273 86868 83339 86869
rect 83222 86804 83228 86868
rect 83292 86866 83339 86868
rect 83292 86864 83384 86866
rect 83334 86808 83384 86864
rect 83292 86806 83384 86808
rect 83292 86804 83339 86806
rect 83273 86803 83339 86804
rect 84377 86324 84443 86325
rect 87137 86324 87203 86325
rect 84326 86322 84332 86324
rect 84286 86262 84332 86322
rect 84396 86320 84443 86324
rect 87086 86322 87092 86324
rect 84438 86264 84443 86320
rect 84326 86260 84332 86262
rect 84396 86260 84443 86264
rect 87046 86262 87092 86322
rect 87156 86320 87203 86324
rect 87198 86264 87203 86320
rect 87086 86260 87092 86262
rect 87156 86260 87203 86264
rect 84377 86259 84443 86260
rect 87137 86259 87203 86260
rect 82854 84900 82860 84964
rect 82924 84962 82930 84964
rect 83406 84962 83412 84964
rect 82924 84902 83412 84962
rect 82924 84900 82930 84902
rect 83406 84900 83412 84902
rect 83476 84900 83482 84964
rect 331121 84826 331187 84829
rect 502558 84826 502564 84828
rect 331121 84824 502564 84826
rect 331121 84768 331126 84824
rect 331182 84768 502564 84824
rect 331121 84766 502564 84768
rect 331121 84763 331187 84766
rect 502558 84764 502564 84766
rect 502628 84764 502634 84828
rect 87454 84220 87460 84284
rect 87524 84282 87530 84284
rect 87638 84282 87644 84284
rect 87524 84222 87644 84282
rect 87524 84220 87530 84222
rect 87638 84220 87644 84222
rect 87708 84220 87714 84284
rect 88006 84084 88012 84148
rect 88076 84084 88082 84148
rect 88014 83876 88074 84084
rect 88006 83812 88012 83876
rect 88076 83812 88082 83876
rect 501086 83058 501092 83060
rect 500358 82998 501092 83058
rect 500358 82924 500418 82998
rect 501086 82996 501092 82998
rect 501156 82996 501162 83060
rect 500350 82860 500356 82924
rect 500420 82860 500426 82924
rect 504265 80204 504331 80205
rect 504214 80140 504220 80204
rect 504284 80202 504331 80204
rect 504284 80200 504376 80202
rect 504326 80144 504376 80200
rect 504284 80142 504376 80144
rect 504284 80140 504331 80142
rect 504265 80139 504331 80140
rect 3417 80066 3483 80069
rect 508262 80066 508268 80068
rect 3417 80064 508268 80066
rect 3417 80008 3422 80064
rect 3478 80008 508268 80064
rect 3417 80006 508268 80008
rect 3417 80003 3483 80006
rect 508262 80004 508268 80006
rect 508332 80004 508338 80068
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 82854 78644 82860 78708
rect 82924 78706 82930 78708
rect 83406 78706 83412 78708
rect 82924 78646 83412 78706
rect 82924 78644 82930 78646
rect 83406 78644 83412 78646
rect 83476 78644 83482 78708
rect 84377 78028 84443 78029
rect 87137 78028 87203 78029
rect 84326 78026 84332 78028
rect 84286 77966 84332 78026
rect 84396 78024 84443 78028
rect 87086 78026 87092 78028
rect 84438 77968 84443 78024
rect 84326 77964 84332 77966
rect 84396 77964 84443 77968
rect 87046 77966 87092 78026
rect 87156 78024 87203 78028
rect 87597 78028 87663 78029
rect 88241 78028 88307 78029
rect 87597 78026 87644 78028
rect 87198 77968 87203 78024
rect 87086 77964 87092 77966
rect 87156 77964 87203 77968
rect 87552 78024 87644 78026
rect 87552 77968 87602 78024
rect 87552 77966 87644 77968
rect 84377 77963 84443 77964
rect 87137 77963 87203 77964
rect 87597 77964 87644 77966
rect 87708 77964 87714 78028
rect 88190 78026 88196 78028
rect 88150 77966 88196 78026
rect 88260 78024 88307 78028
rect 88302 77968 88307 78024
rect 88190 77964 88196 77966
rect 88260 77964 88307 77968
rect 87597 77963 87663 77964
rect 88241 77963 88307 77964
rect 83273 77348 83339 77349
rect 83222 77346 83228 77348
rect 83182 77286 83228 77346
rect 83292 77344 83339 77348
rect 503989 77348 504055 77349
rect 504265 77348 504331 77349
rect 503989 77346 504036 77348
rect 83334 77288 83339 77344
rect 83222 77284 83228 77286
rect 83292 77284 83339 77288
rect 503944 77344 504036 77346
rect 503944 77288 503994 77344
rect 503944 77286 504036 77288
rect 83273 77283 83339 77284
rect 503989 77284 504036 77286
rect 504100 77284 504106 77348
rect 504214 77346 504220 77348
rect 504174 77286 504220 77346
rect 504284 77344 504331 77348
rect 504326 77288 504331 77344
rect 504214 77284 504220 77286
rect 504284 77284 504331 77288
rect 503989 77283 504055 77284
rect 504265 77283 504331 77284
rect 435817 77210 435883 77213
rect 436093 77210 436159 77213
rect 500401 77212 500467 77213
rect 435817 77208 436159 77210
rect 435817 77152 435822 77208
rect 435878 77152 436098 77208
rect 436154 77152 436159 77208
rect 435817 77150 436159 77152
rect 435817 77147 435883 77150
rect 436093 77147 436159 77150
rect 500350 77148 500356 77212
rect 500420 77210 500467 77212
rect 500420 77208 500512 77210
rect 500462 77152 500512 77208
rect 500420 77150 500512 77152
rect 500420 77148 500467 77150
rect 500401 77147 500467 77148
rect 83273 77076 83339 77077
rect 83268 77074 83274 77076
rect 83182 77014 83274 77074
rect 83268 77012 83274 77014
rect 83338 77012 83344 77076
rect 83273 77011 83339 77012
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 499246 72932 499252 72996
rect 499316 72994 499322 72996
rect 499389 72994 499455 72997
rect 499316 72992 499455 72994
rect 499316 72936 499394 72992
rect 499450 72936 499455 72992
rect 499316 72934 499455 72936
rect 499316 72932 499322 72934
rect 499389 72931 499455 72934
rect 117313 71770 117379 71773
rect 117497 71770 117563 71773
rect 117313 71768 117563 71770
rect 117313 71712 117318 71768
rect 117374 71712 117502 71768
rect 117558 71712 117563 71768
rect 117313 71710 117563 71712
rect 117313 71707 117379 71710
rect 117497 71707 117563 71710
rect 120073 71770 120139 71773
rect 120257 71770 120323 71773
rect 120073 71768 120323 71770
rect 120073 71712 120078 71768
rect 120134 71712 120262 71768
rect 120318 71712 120323 71768
rect 120073 71710 120323 71712
rect 120073 71707 120139 71710
rect 120257 71707 120323 71710
rect 152774 70348 152780 70412
rect 152844 70410 152850 70412
rect 152917 70410 152983 70413
rect 152844 70408 152983 70410
rect 152844 70352 152922 70408
rect 152978 70352 152983 70408
rect 152844 70350 152983 70352
rect 152844 70348 152850 70350
rect 152917 70347 152983 70350
rect 88241 69188 88307 69189
rect 88190 69186 88196 69188
rect 88150 69126 88196 69186
rect 88260 69184 88307 69188
rect 88302 69128 88307 69184
rect 88190 69124 88196 69126
rect 88260 69124 88307 69128
rect 88241 69123 88307 69124
rect 500401 68372 500467 68373
rect 500350 68370 500356 68372
rect 500310 68310 500356 68370
rect 500420 68368 500467 68372
rect 500462 68312 500467 68368
rect 500350 68308 500356 68310
rect 500420 68308 500467 68312
rect 500401 68307 500467 68308
rect 179321 67826 179387 67829
rect 179321 67824 179522 67826
rect 179321 67768 179326 67824
rect 179382 67768 179522 67824
rect 179321 67766 179522 67768
rect 179321 67763 179387 67766
rect 83273 67692 83339 67693
rect 83222 67690 83228 67692
rect 83182 67630 83228 67690
rect 83292 67688 83339 67692
rect 83334 67632 83339 67688
rect 83222 67628 83228 67630
rect 83292 67628 83339 67632
rect 83273 67627 83339 67628
rect 87597 67692 87663 67693
rect 152825 67692 152891 67693
rect 87597 67688 87644 67692
rect 87708 67690 87714 67692
rect 87597 67632 87602 67688
rect 87597 67628 87644 67632
rect 87708 67630 87754 67690
rect 87708 67628 87714 67630
rect 152774 67628 152780 67692
rect 152844 67690 152891 67692
rect 179321 67690 179387 67693
rect 179462 67690 179522 67766
rect 152844 67688 152936 67690
rect 152886 67632 152936 67688
rect 152844 67630 152936 67632
rect 179321 67688 179522 67690
rect 179321 67632 179326 67688
rect 179382 67632 179522 67688
rect 179321 67630 179522 67632
rect 435817 67690 435883 67693
rect 436093 67690 436159 67693
rect 435817 67688 436159 67690
rect 435817 67632 435822 67688
rect 435878 67632 436098 67688
rect 436154 67632 436159 67688
rect 435817 67630 436159 67632
rect 152844 67628 152891 67630
rect 87597 67627 87663 67628
rect 152825 67627 152891 67628
rect 179321 67627 179387 67630
rect 435817 67627 435883 67630
rect 436093 67627 436159 67630
rect 498377 67554 498443 67557
rect 498510 67554 498516 67556
rect 498377 67552 498516 67554
rect 498377 67496 498382 67552
rect 498438 67496 498516 67552
rect 498377 67494 498516 67496
rect 498377 67491 498443 67494
rect 498510 67492 498516 67494
rect 498580 67492 498586 67556
rect 85982 67220 85988 67284
rect 86052 67220 86058 67284
rect 85990 67148 86050 67220
rect 85982 67084 85988 67148
rect 86052 67084 86058 67148
rect 82854 65452 82860 65516
rect 82924 65514 82930 65516
rect 83406 65514 83412 65516
rect 82924 65454 83412 65514
rect 82924 65452 82930 65454
rect 83406 65452 83412 65454
rect 83476 65452 83482 65516
rect -960 64562 480 64652
rect 2773 64562 2839 64565
rect -960 64560 2839 64562
rect -960 64504 2778 64560
rect 2834 64504 2839 64560
rect -960 64502 2839 64504
rect -960 64412 480 64502
rect 2773 64499 2839 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 85757 62796 85823 62797
rect 498377 62796 498443 62797
rect 85757 62794 85804 62796
rect 85712 62792 85804 62794
rect 85712 62736 85762 62792
rect 85712 62734 85804 62736
rect 85757 62732 85804 62734
rect 85868 62732 85874 62796
rect 498326 62794 498332 62796
rect 498286 62734 498332 62794
rect 498396 62792 498443 62796
rect 498438 62736 498443 62792
rect 498326 62732 498332 62734
rect 498396 62732 498443 62736
rect 85757 62731 85823 62732
rect 498377 62731 498443 62732
rect 87638 62250 87644 62252
rect 87462 62190 87644 62250
rect 87462 61980 87522 62190
rect 87638 62188 87644 62190
rect 87708 62188 87714 62252
rect 87454 61916 87460 61980
rect 87524 61916 87530 61980
rect 152917 61436 152983 61437
rect 152917 61434 152964 61436
rect 152872 61432 152964 61434
rect 152872 61376 152922 61432
rect 152872 61374 152964 61376
rect 152917 61372 152964 61374
rect 153028 61372 153034 61436
rect 152917 61371 152983 61372
rect 501638 60692 501644 60756
rect 501708 60754 501714 60756
rect 501822 60754 501828 60756
rect 501708 60694 501828 60754
rect 501708 60692 501714 60694
rect 501822 60692 501828 60694
rect 501892 60692 501898 60756
rect 83273 57900 83339 57901
rect 87505 57900 87571 57901
rect 83222 57836 83228 57900
rect 83292 57898 83339 57900
rect 83292 57896 83384 57898
rect 83334 57840 83384 57896
rect 83292 57838 83384 57840
rect 83292 57836 83339 57838
rect 87454 57836 87460 57900
rect 87524 57898 87571 57900
rect 87524 57896 87616 57898
rect 87566 57840 87616 57896
rect 87524 57838 87616 57840
rect 87524 57836 87571 57838
rect 498326 57836 498332 57900
rect 498396 57836 498402 57900
rect 83273 57835 83339 57836
rect 87505 57835 87571 57836
rect 498334 57765 498394 57836
rect 498334 57760 498443 57765
rect 498334 57704 498382 57760
rect 498438 57704 498443 57760
rect 498334 57702 498443 57704
rect 498377 57699 498443 57702
rect 504030 57564 504036 57628
rect 504100 57626 504106 57628
rect 504582 57626 504588 57628
rect 504100 57566 504588 57626
rect 504100 57564 504106 57566
rect 504582 57564 504588 57566
rect 504652 57564 504658 57628
rect 500033 56810 500099 56813
rect 499990 56808 500099 56810
rect 499990 56752 500038 56808
rect 500094 56752 500099 56808
rect 499990 56747 500099 56752
rect 499990 56676 500050 56747
rect 499982 56612 499988 56676
rect 500052 56612 500058 56676
rect 500493 56540 500559 56541
rect 500493 56538 500540 56540
rect 500448 56536 500540 56538
rect 500448 56480 500498 56536
rect 500448 56478 500540 56480
rect 500493 56476 500540 56478
rect 500604 56476 500610 56540
rect 500493 56475 500559 56476
rect 82854 55796 82860 55860
rect 82924 55858 82930 55860
rect 83406 55858 83412 55860
rect 82924 55798 83412 55858
rect 82924 55796 82930 55798
rect 83406 55796 83412 55798
rect 83476 55796 83482 55860
rect 499389 55450 499455 55453
rect 499389 55448 499498 55450
rect 499389 55392 499394 55448
rect 499450 55392 499498 55448
rect 499389 55387 499498 55392
rect 499438 55316 499498 55387
rect 499430 55252 499436 55316
rect 499500 55252 499506 55316
rect 583520 52716 584960 52956
rect 117497 52458 117563 52461
rect 117681 52458 117747 52461
rect 117497 52456 117747 52458
rect 117497 52400 117502 52456
rect 117558 52400 117686 52456
rect 117742 52400 117747 52456
rect 117497 52398 117747 52400
rect 117497 52395 117563 52398
rect 117681 52395 117747 52398
rect 120257 52458 120323 52461
rect 120441 52458 120507 52461
rect 120257 52456 120507 52458
rect 120257 52400 120262 52456
rect 120318 52400 120446 52456
rect 120502 52400 120507 52456
rect 120257 52398 120507 52400
rect 120257 52395 120323 52398
rect 120441 52395 120507 52398
rect 153009 50964 153075 50965
rect 152958 50962 152964 50964
rect 152918 50902 152964 50962
rect 153028 50960 153075 50964
rect 153070 50904 153075 50960
rect 152958 50900 152964 50902
rect 153028 50900 153075 50904
rect 153009 50899 153075 50900
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 499941 49060 500007 49061
rect 500401 49060 500467 49061
rect 499941 49058 499988 49060
rect 499896 49056 499988 49058
rect 499896 49000 499946 49056
rect 499896 48998 499988 49000
rect 499941 48996 499988 48998
rect 500052 48996 500058 49060
rect 500350 49058 500356 49060
rect 500310 48998 500356 49058
rect 500420 49056 500467 49060
rect 500462 49000 500467 49056
rect 500350 48996 500356 48998
rect 500420 48996 500467 49000
rect 499941 48995 500007 48996
rect 500401 48995 500467 48996
rect 503989 49058 504055 49061
rect 504214 49058 504220 49060
rect 503989 49056 504220 49058
rect 503989 49000 503994 49056
rect 504050 49000 504220 49056
rect 503989 48998 504220 49000
rect 503989 48995 504055 48998
rect 504214 48996 504220 48998
rect 504284 48996 504290 49060
rect 504449 49058 504515 49061
rect 504582 49058 504588 49060
rect 504449 49056 504588 49058
rect 504449 49000 504454 49056
rect 504510 49000 504588 49056
rect 504449 48998 504588 49000
rect 504449 48995 504515 48998
rect 504582 48996 504588 48998
rect 504652 48996 504658 49060
rect 500493 48924 500559 48925
rect 500493 48922 500540 48924
rect 500448 48920 500540 48922
rect 500448 48864 500498 48920
rect 500448 48862 500540 48864
rect 500493 48860 500540 48862
rect 500604 48860 500610 48924
rect 500493 48859 500559 48860
rect 85757 48514 85823 48517
rect 85757 48512 85866 48514
rect 85757 48456 85762 48512
rect 85818 48456 85866 48512
rect 85757 48451 85866 48456
rect 83273 48380 83339 48381
rect 85806 48380 85866 48451
rect 87505 48380 87571 48381
rect 83222 48378 83228 48380
rect 83182 48318 83228 48378
rect 83292 48376 83339 48380
rect 83334 48320 83339 48376
rect 83222 48316 83228 48318
rect 83292 48316 83339 48320
rect 85798 48316 85804 48380
rect 85868 48316 85874 48380
rect 87454 48378 87460 48380
rect 87414 48318 87460 48378
rect 87524 48376 87571 48380
rect 87566 48320 87571 48376
rect 87454 48316 87460 48318
rect 87524 48316 87571 48320
rect 83273 48315 83339 48316
rect 87505 48315 87571 48316
rect 498377 48378 498443 48381
rect 498510 48378 498516 48380
rect 498377 48376 498516 48378
rect 498377 48320 498382 48376
rect 498438 48320 498516 48376
rect 498377 48318 498516 48320
rect 498377 48315 498443 48318
rect 498510 48316 498516 48318
rect 498580 48316 498586 48380
rect 85982 48044 85988 48108
rect 86052 48044 86058 48108
rect 85990 47836 86050 48044
rect 85982 47772 85988 47836
rect 86052 47772 86058 47836
rect 498510 44434 498516 44436
rect 498334 44374 498516 44434
rect 498334 44300 498394 44374
rect 498510 44372 498516 44374
rect 498580 44372 498586 44436
rect 498326 44236 498332 44300
rect 498396 44236 498402 44300
rect 85849 43484 85915 43485
rect 85798 43482 85804 43484
rect 85758 43422 85804 43482
rect 85868 43480 85915 43484
rect 85910 43424 85915 43480
rect 85798 43420 85804 43422
rect 85868 43420 85915 43424
rect 85849 43419 85915 43420
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 86718 40218 86724 40220
rect 86542 40158 86724 40218
rect 86542 39948 86602 40158
rect 86718 40156 86724 40158
rect 86788 40156 86794 40220
rect 87454 40218 87460 40220
rect 87278 40158 87460 40218
rect 87278 39948 87338 40158
rect 87454 40156 87460 40158
rect 87524 40156 87530 40220
rect 84326 39884 84332 39948
rect 84396 39946 84402 39948
rect 84510 39946 84516 39948
rect 84396 39886 84516 39946
rect 84396 39884 84402 39886
rect 84510 39884 84516 39886
rect 84580 39884 84586 39948
rect 86534 39884 86540 39948
rect 86604 39884 86610 39948
rect 87270 39884 87276 39948
rect 87340 39884 87346 39948
rect 453941 39266 454007 39269
rect 500401 39266 500467 39269
rect 453941 39264 500467 39266
rect 453941 39208 453946 39264
rect 454002 39208 500406 39264
rect 500462 39208 500467 39264
rect 453941 39206 500467 39208
rect 453941 39203 454007 39206
rect 500401 39203 500467 39206
rect 499941 38858 500007 38861
rect 503989 38858 504055 38861
rect 499941 38856 500050 38858
rect 499941 38800 499946 38856
rect 500002 38800 500050 38856
rect 499941 38795 500050 38800
rect 503989 38856 504282 38858
rect 503989 38800 503994 38856
rect 504050 38800 504282 38856
rect 503989 38798 504282 38800
rect 503989 38795 504055 38798
rect 499990 38724 500050 38795
rect 504222 38724 504282 38798
rect 504449 38724 504515 38725
rect 499982 38660 499988 38724
rect 500052 38660 500058 38724
rect 504214 38660 504220 38724
rect 504284 38660 504290 38724
rect 504398 38660 504404 38724
rect 504468 38722 504515 38724
rect 504468 38720 504560 38722
rect 504510 38664 504560 38720
rect 504468 38662 504560 38664
rect 504468 38660 504515 38662
rect 504449 38659 504515 38660
rect 83273 38588 83339 38589
rect 83222 38524 83228 38588
rect 83292 38586 83339 38588
rect 83292 38584 83384 38586
rect 83334 38528 83384 38584
rect 83292 38526 83384 38528
rect 83292 38524 83339 38526
rect 83273 38523 83339 38524
rect 85849 37498 85915 37501
rect 85806 37496 85915 37498
rect 85806 37440 85854 37496
rect 85910 37440 85915 37496
rect 85806 37435 85915 37440
rect 85806 37364 85866 37435
rect 85798 37300 85804 37364
rect 85868 37300 85874 37364
rect 220261 37362 220327 37365
rect 220445 37362 220511 37365
rect 220261 37360 220511 37362
rect 220261 37304 220266 37360
rect 220322 37304 220450 37360
rect 220506 37304 220511 37360
rect 220261 37302 220511 37304
rect 220261 37299 220327 37302
rect 220445 37299 220511 37302
rect 499430 37300 499436 37364
rect 499500 37300 499506 37364
rect 499438 37090 499498 37300
rect 500585 37228 500651 37229
rect 500534 37164 500540 37228
rect 500604 37226 500651 37228
rect 500604 37224 500696 37226
rect 500646 37168 500696 37224
rect 500604 37166 500696 37168
rect 500604 37164 500651 37166
rect 500585 37163 500651 37164
rect 499614 37090 499620 37092
rect 499438 37030 499620 37090
rect 499614 37028 499620 37030
rect 499684 37028 499690 37092
rect -960 35866 480 35956
rect 3141 35866 3207 35869
rect -960 35864 3207 35866
rect -960 35808 3146 35864
rect 3202 35808 3207 35864
rect -960 35806 3207 35808
rect -960 35716 480 35806
rect 3141 35803 3207 35806
rect 87270 35260 87276 35324
rect 87340 35322 87346 35324
rect 87505 35322 87571 35325
rect 87340 35320 87571 35322
rect 87340 35264 87510 35320
rect 87566 35264 87571 35320
rect 87340 35262 87571 35264
rect 87340 35260 87346 35262
rect 87505 35259 87571 35262
rect 83406 35124 83412 35188
rect 83476 35186 83482 35188
rect 425605 35186 425671 35189
rect 83476 35184 425671 35186
rect 83476 35128 425610 35184
rect 425666 35128 425671 35184
rect 83476 35126 425671 35128
rect 83476 35124 83482 35126
rect 425605 35123 425671 35126
rect 498285 34372 498351 34373
rect 498285 34370 498332 34372
rect 498240 34368 498332 34370
rect 498240 34312 498290 34368
rect 498240 34310 498332 34312
rect 498285 34308 498332 34310
rect 498396 34308 498402 34372
rect 498285 34307 498351 34308
rect 500585 29748 500651 29749
rect 499982 29684 499988 29748
rect 500052 29746 500058 29748
rect 500350 29746 500356 29748
rect 500052 29686 500356 29746
rect 500052 29684 500058 29686
rect 500350 29684 500356 29686
rect 500420 29684 500426 29748
rect 500534 29746 500540 29748
rect 500494 29686 500540 29746
rect 500604 29744 500651 29748
rect 500646 29688 500651 29744
rect 500534 29684 500540 29686
rect 500604 29684 500651 29688
rect 500585 29683 500651 29684
rect 583520 29338 584960 29428
rect 518942 29278 528570 29338
rect 83273 29202 83339 29205
rect 83230 29200 83339 29202
rect 83230 29144 83278 29200
rect 83334 29144 83339 29200
rect 83230 29139 83339 29144
rect 83230 29068 83290 29139
rect 83222 29004 83228 29068
rect 83292 29004 83298 29068
rect 505870 29004 505876 29068
rect 505940 29066 505946 29068
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 557582 29278 567210 29338
rect 528510 29142 538138 29202
rect 505940 29006 519002 29066
rect 538078 29066 538138 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 538078 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 505940 29004 505946 29006
rect 85849 27572 85915 27573
rect 85798 27508 85804 27572
rect 85868 27570 85915 27572
rect 85868 27568 85960 27570
rect 85910 27512 85960 27568
rect 85868 27510 85960 27512
rect 85868 27508 85915 27510
rect 85849 27507 85915 27508
rect 497038 26346 497044 26348
rect 496862 26286 497044 26346
rect 496862 26076 496922 26286
rect 497038 26284 497044 26286
rect 497108 26284 497114 26348
rect 496854 26012 496860 26076
rect 496924 26012 496930 26076
rect 498285 25122 498351 25125
rect 498285 25120 498394 25122
rect 498285 25064 498290 25120
rect 498346 25064 498394 25120
rect 498285 25059 498394 25064
rect 498334 24988 498394 25059
rect 498326 24924 498332 24988
rect 498396 24924 498402 24988
rect 120073 24850 120139 24853
rect 120349 24850 120415 24853
rect 120073 24848 120415 24850
rect 120073 24792 120078 24848
rect 120134 24792 120354 24848
rect 120410 24792 120415 24848
rect 120073 24790 120415 24792
rect 120073 24787 120139 24790
rect 120349 24787 120415 24790
rect 87505 23492 87571 23493
rect 84326 23428 84332 23492
rect 84396 23490 84402 23492
rect 84510 23490 84516 23492
rect 84396 23430 84516 23490
rect 84396 23428 84402 23430
rect 84510 23428 84516 23430
rect 84580 23428 84586 23492
rect 87454 23490 87460 23492
rect 87414 23430 87460 23490
rect 87524 23488 87571 23492
rect 87566 23432 87571 23488
rect 87454 23428 87460 23430
rect 87524 23428 87571 23432
rect 87505 23427 87571 23428
rect 84377 23356 84443 23357
rect 84326 23292 84332 23356
rect 84396 23354 84443 23356
rect 84396 23352 84488 23354
rect 84438 23296 84488 23352
rect 84396 23294 84488 23296
rect 84396 23292 84443 23294
rect 84377 23291 84443 23292
rect 86401 22810 86467 22813
rect 86534 22810 86540 22812
rect 86401 22808 86540 22810
rect 86401 22752 86406 22808
rect 86462 22752 86540 22808
rect 86401 22750 86540 22752
rect 86401 22747 86467 22750
rect 86534 22748 86540 22750
rect 86604 22748 86610 22812
rect 507894 21994 507900 21996
rect 614 21934 507900 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 507894 21932 507900 21934
rect 507964 21932 507970 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 85941 19276 86007 19277
rect 83222 19212 83228 19276
rect 83292 19212 83298 19276
rect 85941 19274 85988 19276
rect 85896 19272 85988 19274
rect 85896 19216 85946 19272
rect 85896 19214 85988 19216
rect 85941 19212 85988 19214
rect 86052 19212 86058 19276
rect 83230 19141 83290 19212
rect 85941 19211 86007 19212
rect 83230 19136 83339 19141
rect 83230 19080 83278 19136
rect 83334 19080 83339 19136
rect 83230 19078 83339 19080
rect 83273 19075 83339 19078
rect 297909 19138 297975 19141
rect 315941 19138 316007 19141
rect 297909 19136 316007 19138
rect 297909 19080 297914 19136
rect 297970 19080 315946 19136
rect 316002 19080 316007 19136
rect 297909 19078 316007 19080
rect 297909 19075 297975 19078
rect 315941 19075 316007 19078
rect 325693 19138 325759 19141
rect 335905 19138 335971 19141
rect 325693 19136 335971 19138
rect 325693 19080 325698 19136
rect 325754 19080 335910 19136
rect 335966 19080 335971 19136
rect 325693 19078 335971 19080
rect 325693 19075 325759 19078
rect 335905 19075 335971 19078
rect 345013 19138 345079 19141
rect 355317 19138 355383 19141
rect 345013 19136 355383 19138
rect 345013 19080 345018 19136
rect 345074 19080 355322 19136
rect 355378 19080 355383 19136
rect 345013 19078 355383 19080
rect 345013 19075 345079 19078
rect 355317 19075 355383 19078
rect 364333 19138 364399 19141
rect 378777 19138 378843 19141
rect 364333 19136 378843 19138
rect 364333 19080 364338 19136
rect 364394 19080 378782 19136
rect 378838 19080 378843 19136
rect 364333 19078 378843 19080
rect 364333 19075 364399 19078
rect 378777 19075 378843 19078
rect 383653 19138 383719 19141
rect 412541 19138 412607 19141
rect 383653 19136 412607 19138
rect 383653 19080 383658 19136
rect 383714 19080 412546 19136
rect 412602 19080 412607 19136
rect 383653 19078 412607 19080
rect 383653 19075 383719 19078
rect 412541 19075 412607 19078
rect 422293 19138 422359 19141
rect 432045 19138 432111 19141
rect 422293 19136 432111 19138
rect 422293 19080 422298 19136
rect 422354 19080 432050 19136
rect 432106 19080 432111 19136
rect 422293 19078 432111 19080
rect 422293 19075 422359 19078
rect 432045 19075 432111 19078
rect 441613 19138 441679 19141
rect 447133 19138 447199 19141
rect 441613 19136 447199 19138
rect 441613 19080 441618 19136
rect 441674 19080 447138 19136
rect 447194 19080 447199 19136
rect 441613 19078 447199 19080
rect 441613 19075 441679 19078
rect 447133 19075 447199 19078
rect 478137 19138 478203 19141
rect 485681 19138 485747 19141
rect 478137 19136 485747 19138
rect 478137 19080 478142 19136
rect 478198 19080 485686 19136
rect 485742 19080 485747 19136
rect 478137 19078 485747 19080
rect 478137 19075 478203 19078
rect 485681 19075 485747 19078
rect 314561 19002 314627 19005
rect 498878 19002 498884 19004
rect 314561 19000 498884 19002
rect 314561 18944 314566 19000
rect 314622 18944 498884 19000
rect 314561 18942 498884 18944
rect 314561 18939 314627 18942
rect 498878 18940 498884 18942
rect 498948 18940 498954 19004
rect 315941 18866 316007 18869
rect 325693 18866 325759 18869
rect 315941 18864 325759 18866
rect 315941 18808 315946 18864
rect 316002 18808 325698 18864
rect 325754 18808 325759 18864
rect 315941 18806 325759 18808
rect 315941 18803 316007 18806
rect 325693 18803 325759 18806
rect 335905 18866 335971 18869
rect 345013 18866 345079 18869
rect 335905 18864 345079 18866
rect 335905 18808 335910 18864
rect 335966 18808 345018 18864
rect 345074 18808 345079 18864
rect 335905 18806 345079 18808
rect 335905 18803 335971 18806
rect 345013 18803 345079 18806
rect 355317 18866 355383 18869
rect 364333 18866 364399 18869
rect 355317 18864 364399 18866
rect 355317 18808 355322 18864
rect 355378 18808 364338 18864
rect 364394 18808 364399 18864
rect 355317 18806 364399 18808
rect 355317 18803 355383 18806
rect 364333 18803 364399 18806
rect 378777 18866 378843 18869
rect 383653 18866 383719 18869
rect 378777 18864 383719 18866
rect 378777 18808 378782 18864
rect 378838 18808 383658 18864
rect 383714 18808 383719 18864
rect 378777 18806 383719 18808
rect 378777 18803 378843 18806
rect 383653 18803 383719 18806
rect 412541 18866 412607 18869
rect 422293 18866 422359 18869
rect 412541 18864 422359 18866
rect 412541 18808 412546 18864
rect 412602 18808 422298 18864
rect 422354 18808 422359 18864
rect 412541 18806 422359 18808
rect 412541 18803 412607 18806
rect 422293 18803 422359 18806
rect 432045 18866 432111 18869
rect 441613 18866 441679 18869
rect 432045 18864 441679 18866
rect 432045 18808 432050 18864
rect 432106 18808 441618 18864
rect 441674 18808 441679 18864
rect 432045 18806 441679 18808
rect 432045 18803 432111 18806
rect 441613 18803 441679 18806
rect 447133 18866 447199 18869
rect 462589 18866 462655 18869
rect 447133 18864 462655 18866
rect 447133 18808 447138 18864
rect 447194 18808 462594 18864
rect 462650 18808 462655 18864
rect 447133 18806 462655 18808
rect 447133 18803 447199 18806
rect 462589 18803 462655 18806
rect 87454 18668 87460 18732
rect 87524 18730 87530 18732
rect 448513 18730 448579 18733
rect 87524 18728 448579 18730
rect 87524 18672 448518 18728
rect 448574 18672 448579 18728
rect 87524 18670 448579 18672
rect 87524 18668 87530 18670
rect 448513 18667 448579 18670
rect 485681 18730 485747 18733
rect 499614 18730 499620 18732
rect 485681 18728 499620 18730
rect 485681 18672 485686 18728
rect 485742 18672 499620 18728
rect 485681 18670 499620 18672
rect 485681 18667 485747 18670
rect 499614 18668 499620 18670
rect 499684 18668 499690 18732
rect 64689 18594 64755 18597
rect 505502 18594 505508 18596
rect 64689 18592 505508 18594
rect 64689 18536 64694 18592
rect 64750 18536 505508 18592
rect 64689 18534 505508 18536
rect 64689 18531 64755 18534
rect 505502 18532 505508 18534
rect 505572 18532 505578 18596
rect 462589 18458 462655 18461
rect 478137 18458 478203 18461
rect 462589 18456 478203 18458
rect 462589 18400 462594 18456
rect 462650 18400 478142 18456
rect 478198 18400 478203 18456
rect 462589 18398 478203 18400
rect 462589 18395 462655 18398
rect 478137 18395 478203 18398
rect 85849 18186 85915 18189
rect 85622 18184 85915 18186
rect 85622 18128 85854 18184
rect 85910 18128 85915 18184
rect 85622 18126 85915 18128
rect 85622 18052 85682 18126
rect 85849 18123 85915 18126
rect 85614 17988 85620 18052
rect 85684 17988 85690 18052
rect 580257 17642 580323 17645
rect 583520 17642 584960 17732
rect 580257 17640 584960 17642
rect 580257 17584 580262 17640
rect 580318 17584 584960 17640
rect 580257 17582 584960 17584
rect 580257 17579 580323 17582
rect 190361 17506 190427 17509
rect 503662 17506 503668 17508
rect 190361 17504 503668 17506
rect 190361 17448 190366 17504
rect 190422 17448 503668 17504
rect 190361 17446 503668 17448
rect 190361 17443 190427 17446
rect 503662 17444 503668 17446
rect 503732 17444 503738 17508
rect 583520 17492 584960 17582
rect 165521 17370 165587 17373
rect 503846 17370 503852 17372
rect 165521 17368 503852 17370
rect 165521 17312 165526 17368
rect 165582 17312 503852 17368
rect 165521 17310 503852 17312
rect 165521 17307 165587 17310
rect 503846 17308 503852 17310
rect 503916 17308 503922 17372
rect 79174 17172 79180 17236
rect 79244 17234 79250 17236
rect 481725 17234 481791 17237
rect 79244 17232 481791 17234
rect 79244 17176 481730 17232
rect 481786 17176 481791 17232
rect 79244 17174 481791 17176
rect 79244 17172 79250 17174
rect 481725 17171 481791 17174
rect 204161 16418 204227 16421
rect 503110 16418 503116 16420
rect 204161 16416 503116 16418
rect 204161 16360 204166 16416
rect 204222 16360 503116 16416
rect 204161 16358 503116 16360
rect 204161 16355 204227 16358
rect 503110 16356 503116 16358
rect 503180 16356 503186 16420
rect 199929 16282 199995 16285
rect 502374 16282 502380 16284
rect 199929 16280 502380 16282
rect 199929 16224 199934 16280
rect 199990 16224 502380 16280
rect 199929 16222 502380 16224
rect 199929 16219 199995 16222
rect 502374 16220 502380 16222
rect 502444 16220 502450 16284
rect 99097 16146 99163 16149
rect 504214 16146 504220 16148
rect 99097 16144 504220 16146
rect 99097 16088 99102 16144
rect 99158 16088 504220 16144
rect 99097 16086 504220 16088
rect 99097 16083 99163 16086
rect 504214 16084 504220 16086
rect 504284 16084 504290 16148
rect 83917 16010 83983 16013
rect 500534 16010 500540 16012
rect 83917 16008 500540 16010
rect 83917 15952 83922 16008
rect 83978 15952 500540 16008
rect 83917 15950 500540 15952
rect 83917 15947 83983 15950
rect 500534 15948 500540 15950
rect 500604 15948 500610 16012
rect 83273 15874 83339 15877
rect 560293 15874 560359 15877
rect 83273 15872 560359 15874
rect 83273 15816 83278 15872
rect 83334 15816 560298 15872
rect 560354 15816 560359 15872
rect 83273 15814 560359 15816
rect 83273 15811 83339 15814
rect 560293 15811 560359 15814
rect 498326 15268 498332 15332
rect 498396 15330 498402 15332
rect 498469 15330 498535 15333
rect 498396 15328 498535 15330
rect 498396 15272 498474 15328
rect 498530 15272 498535 15328
rect 498396 15270 498535 15272
rect 498396 15268 498402 15270
rect 498469 15267 498535 15270
rect 499941 15194 500007 15197
rect 500217 15194 500283 15197
rect 499941 15192 500283 15194
rect 499941 15136 499946 15192
rect 500002 15136 500222 15192
rect 500278 15136 500283 15192
rect 499941 15134 500283 15136
rect 499941 15131 500007 15134
rect 500217 15131 500283 15134
rect 195421 14650 195487 14653
rect 502742 14650 502748 14652
rect 195421 14648 502748 14650
rect 195421 14592 195426 14648
rect 195482 14592 502748 14648
rect 195421 14590 502748 14592
rect 195421 14587 195487 14590
rect 502742 14588 502748 14590
rect 502812 14588 502818 14652
rect 81014 14452 81020 14516
rect 81084 14514 81090 14516
rect 553393 14514 553459 14517
rect 81084 14512 553459 14514
rect 81084 14456 553398 14512
rect 553454 14456 553459 14512
rect 81084 14454 553459 14456
rect 81084 14452 81090 14454
rect 553393 14451 553459 14454
rect 82721 13970 82787 13973
rect 82678 13968 82787 13970
rect 82678 13912 82726 13968
rect 82782 13912 82787 13968
rect 82678 13907 82787 13912
rect 82678 13837 82738 13907
rect 82629 13832 82738 13837
rect 84377 13836 84443 13837
rect 84326 13834 84332 13836
rect 82629 13776 82634 13832
rect 82690 13776 82738 13832
rect 82629 13774 82738 13776
rect 84286 13774 84332 13834
rect 84396 13832 84443 13836
rect 84438 13776 84443 13832
rect 82629 13771 82695 13774
rect 84326 13772 84332 13774
rect 84396 13772 84443 13776
rect 84377 13771 84443 13772
rect 84377 13700 84443 13701
rect 84326 13636 84332 13700
rect 84396 13698 84443 13700
rect 84396 13696 84488 13698
rect 84438 13640 84488 13696
rect 84396 13638 84488 13640
rect 84396 13636 84443 13638
rect 84377 13635 84443 13636
rect 83038 12956 83044 13020
rect 83108 13018 83114 13020
rect 538213 13018 538279 13021
rect 83108 13016 538279 13018
rect 83108 12960 538218 13016
rect 538274 12960 538279 13016
rect 83108 12958 538279 12960
rect 83108 12956 83114 12958
rect 538213 12955 538279 12958
rect 82118 11732 82124 11796
rect 82188 11794 82194 11796
rect 437473 11794 437539 11797
rect 82188 11792 437539 11794
rect 82188 11736 437478 11792
rect 437534 11736 437539 11792
rect 82188 11734 437539 11736
rect 82188 11732 82194 11734
rect 437473 11731 437539 11734
rect 81750 11596 81756 11660
rect 81820 11658 81826 11660
rect 512085 11658 512151 11661
rect 81820 11656 512151 11658
rect 81820 11600 512090 11656
rect 512146 11600 512151 11656
rect 81820 11598 512151 11600
rect 81820 11596 81826 11598
rect 512085 11595 512151 11598
rect 79726 10508 79732 10572
rect 79796 10570 79802 10572
rect 369209 10570 369275 10573
rect 79796 10568 369275 10570
rect 79796 10512 369214 10568
rect 369270 10512 369275 10568
rect 79796 10510 369275 10512
rect 79796 10508 79802 10510
rect 369209 10507 369275 10510
rect 81566 10372 81572 10436
rect 81636 10434 81642 10436
rect 433517 10434 433583 10437
rect 81636 10432 433583 10434
rect 81636 10376 433522 10432
rect 433578 10376 433583 10432
rect 81636 10374 433583 10376
rect 81636 10372 81642 10374
rect 433517 10371 433583 10374
rect 151721 10298 151787 10301
rect 504398 10298 504404 10300
rect 151721 10296 504404 10298
rect 151721 10240 151726 10296
rect 151782 10240 504404 10296
rect 151721 10238 504404 10240
rect 151721 10235 151787 10238
rect 504398 10236 504404 10238
rect 504468 10236 504474 10300
rect 85614 9828 85620 9892
rect 85684 9890 85690 9892
rect 85941 9890 86007 9893
rect 223573 9890 223639 9893
rect 85684 9830 85866 9890
rect 85684 9828 85690 9830
rect 85806 9756 85866 9830
rect 85941 9888 86050 9890
rect 85941 9832 85946 9888
rect 86002 9832 86050 9888
rect 85941 9827 86050 9832
rect 85990 9756 86050 9827
rect 223438 9888 223639 9890
rect 223438 9832 223578 9888
rect 223634 9832 223639 9888
rect 223438 9830 223639 9832
rect 85798 9692 85804 9756
rect 85868 9692 85874 9756
rect 85982 9692 85988 9756
rect 86052 9692 86058 9756
rect 195421 9754 195487 9757
rect 195605 9754 195671 9757
rect 195421 9752 195671 9754
rect 195421 9696 195426 9752
rect 195482 9696 195610 9752
rect 195666 9696 195671 9752
rect 195421 9694 195671 9696
rect 195421 9691 195487 9694
rect 195605 9691 195671 9694
rect 223438 9720 223498 9830
rect 223573 9827 223639 9830
rect 258073 9754 258139 9757
rect 258257 9754 258323 9757
rect 258073 9752 258323 9754
rect 223573 9720 223639 9723
rect 223438 9718 223639 9720
rect 223438 9662 223578 9718
rect 223634 9662 223639 9718
rect 258073 9696 258078 9752
rect 258134 9696 258262 9752
rect 258318 9696 258323 9752
rect 258073 9694 258323 9696
rect 258073 9691 258139 9694
rect 258257 9691 258323 9694
rect 427629 9754 427695 9757
rect 427813 9754 427879 9757
rect 498469 9756 498535 9757
rect 498469 9754 498516 9756
rect 427629 9752 427879 9754
rect 427629 9696 427634 9752
rect 427690 9696 427818 9752
rect 427874 9696 427879 9752
rect 427629 9694 427879 9696
rect 498424 9752 498516 9754
rect 498424 9696 498474 9752
rect 498424 9694 498516 9696
rect 427629 9691 427695 9694
rect 427813 9691 427879 9694
rect 498469 9692 498516 9694
rect 498580 9692 498586 9756
rect 498469 9691 498535 9692
rect 223438 9660 223639 9662
rect 223573 9657 223639 9660
rect 85982 9420 85988 9484
rect 86052 9482 86058 9484
rect 86217 9482 86283 9485
rect 86052 9480 86283 9482
rect 86052 9424 86222 9480
rect 86278 9424 86283 9480
rect 86052 9422 86283 9424
rect 86052 9420 86058 9422
rect 86217 9419 86283 9422
rect 91686 8876 91692 8940
rect 91756 8938 91762 8940
rect 290733 8938 290799 8941
rect 91756 8936 290799 8938
rect 91756 8880 290738 8936
rect 290794 8880 290799 8936
rect 91756 8878 290799 8880
rect 91756 8876 91762 8878
rect 290733 8875 290799 8878
rect 353753 8938 353819 8941
rect 500350 8938 500356 8940
rect 353753 8936 500356 8938
rect 353753 8880 353758 8936
rect 353814 8880 500356 8936
rect 353753 8878 500356 8880
rect 353753 8875 353819 8878
rect 500350 8876 500356 8878
rect 500420 8876 500426 8940
rect 85798 8196 85804 8260
rect 85868 8196 85874 8260
rect 223573 8258 223639 8261
rect 223438 8256 223639 8258
rect 223438 8200 223578 8256
rect 223634 8200 223639 8256
rect 223438 8198 223639 8200
rect 85806 8122 85866 8196
rect 87781 8122 87847 8125
rect 85806 8120 87847 8122
rect 85806 8064 87786 8120
rect 87842 8064 87847 8120
rect 85806 8062 87847 8064
rect 223438 8122 223498 8198
rect 223573 8195 223639 8198
rect 289721 8258 289787 8261
rect 289905 8258 289971 8261
rect 289721 8256 289971 8258
rect 289721 8200 289726 8256
rect 289782 8200 289910 8256
rect 289966 8200 289971 8256
rect 289721 8198 289971 8200
rect 289721 8195 289787 8198
rect 289905 8195 289971 8198
rect 224217 8122 224283 8125
rect 223438 8120 224283 8122
rect 223438 8064 224222 8120
rect 224278 8064 224283 8120
rect 223438 8062 224283 8064
rect 87781 8059 87847 8062
rect 224217 8059 224283 8062
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 80053 6898 80119 6901
rect 80329 6898 80395 6901
rect 80053 6896 80395 6898
rect 80053 6840 80058 6896
rect 80114 6840 80334 6896
rect 80390 6840 80395 6896
rect 80053 6838 80395 6840
rect 80053 6835 80119 6838
rect 80329 6835 80395 6838
rect 93158 6836 93164 6900
rect 93228 6898 93234 6900
rect 387057 6898 387123 6901
rect 93228 6896 387123 6898
rect 93228 6840 387062 6896
rect 387118 6840 387123 6896
rect 93228 6838 387123 6840
rect 93228 6836 93234 6838
rect 387057 6835 387123 6838
rect 465625 6898 465691 6901
rect 510654 6898 510660 6900
rect 465625 6896 510660 6898
rect 465625 6840 465630 6896
rect 465686 6840 510660 6896
rect 465625 6838 510660 6840
rect 465625 6835 465691 6838
rect 510654 6836 510660 6838
rect 510724 6836 510730 6900
rect 85430 6700 85436 6764
rect 85500 6762 85506 6764
rect 390645 6762 390711 6765
rect 85500 6760 390711 6762
rect 85500 6704 390650 6760
rect 390706 6704 390711 6760
rect 85500 6702 390711 6704
rect 85500 6700 85506 6702
rect 390645 6699 390711 6702
rect 407297 6762 407363 6765
rect 496854 6762 496860 6764
rect 407297 6760 496860 6762
rect 407297 6704 407302 6760
rect 407358 6704 496860 6760
rect 407297 6702 496860 6704
rect 407297 6699 407363 6702
rect 496854 6700 496860 6702
rect 496924 6700 496930 6764
rect 79358 6564 79364 6628
rect 79428 6626 79434 6628
rect 389449 6626 389515 6629
rect 79428 6624 389515 6626
rect 79428 6568 389454 6624
rect 389510 6568 389515 6624
rect 79428 6566 389515 6568
rect 79428 6564 79434 6566
rect 389449 6563 389515 6566
rect 403709 6626 403775 6629
rect 507526 6626 507532 6628
rect 403709 6624 507532 6626
rect 403709 6568 403714 6624
rect 403770 6568 507532 6624
rect 403709 6566 507532 6568
rect 403709 6563 403775 6566
rect 507526 6564 507532 6566
rect 507596 6564 507602 6628
rect 81382 6428 81388 6492
rect 81452 6490 81458 6492
rect 414473 6490 414539 6493
rect 81452 6488 414539 6490
rect 81452 6432 414478 6488
rect 414534 6432 414539 6488
rect 81452 6430 414539 6432
rect 81452 6428 81458 6430
rect 414473 6427 414539 6430
rect 422753 6490 422819 6493
rect 497406 6490 497412 6492
rect 422753 6488 497412 6490
rect 422753 6432 422758 6488
rect 422814 6432 497412 6488
rect 422753 6430 497412 6432
rect 422753 6427 422819 6430
rect 497406 6428 497412 6430
rect 497476 6428 497482 6492
rect 79542 6292 79548 6356
rect 79612 6354 79618 6356
rect 535729 6354 535795 6357
rect 79612 6352 535795 6354
rect 79612 6296 535734 6352
rect 535790 6296 535795 6352
rect 79612 6294 535795 6296
rect 79612 6292 79618 6294
rect 535729 6291 535795 6294
rect 81934 6156 81940 6220
rect 82004 6218 82010 6220
rect 561949 6218 562015 6221
rect 82004 6216 562015 6218
rect 82004 6160 561954 6216
rect 562010 6160 562015 6216
rect 82004 6158 562015 6160
rect 82004 6156 82010 6158
rect 561949 6155 562015 6158
rect 88006 6020 88012 6084
rect 88076 6082 88082 6084
rect 325233 6082 325299 6085
rect 88076 6080 325299 6082
rect 88076 6024 325238 6080
rect 325294 6024 325299 6080
rect 88076 6022 325299 6024
rect 88076 6020 88082 6022
rect 325233 6019 325299 6022
rect 470317 6082 470383 6085
rect 509182 6082 509188 6084
rect 470317 6080 509188 6082
rect 470317 6024 470322 6080
rect 470378 6024 509188 6080
rect 470317 6022 509188 6024
rect 470317 6019 470383 6022
rect 509182 6020 509188 6022
rect 509252 6020 509258 6084
rect 92054 5884 92060 5948
rect 92124 5946 92130 5948
rect 318057 5946 318123 5949
rect 92124 5944 318123 5946
rect 92124 5888 318062 5944
rect 318118 5888 318123 5944
rect 92124 5886 318123 5888
rect 92124 5884 92130 5886
rect 318057 5883 318123 5886
rect 87781 5810 87847 5813
rect 230105 5810 230171 5813
rect 498510 5810 498516 5812
rect 87781 5808 230171 5810
rect 87781 5752 87786 5808
rect 87842 5752 230110 5808
rect 230166 5752 230171 5808
rect 87781 5750 230171 5752
rect 87781 5747 87847 5750
rect 230105 5747 230171 5750
rect 498334 5750 498516 5810
rect 498334 5676 498394 5750
rect 498510 5748 498516 5750
rect 498580 5748 498586 5812
rect 583520 5796 584960 6036
rect 498326 5612 498332 5676
rect 498396 5612 498402 5676
rect 82629 5402 82695 5405
rect 92974 5402 92980 5404
rect 82629 5400 92980 5402
rect 82629 5344 82634 5400
rect 82690 5344 92980 5400
rect 82629 5342 92980 5344
rect 82629 5339 82695 5342
rect 92974 5340 92980 5342
rect 93044 5340 93050 5404
rect 89294 5204 89300 5268
rect 89364 5266 89370 5268
rect 266997 5266 267063 5269
rect 89364 5264 267063 5266
rect 89364 5208 267002 5264
rect 267058 5208 267063 5264
rect 89364 5206 267063 5208
rect 89364 5204 89370 5206
rect 266997 5203 267063 5206
rect 90398 5068 90404 5132
rect 90468 5130 90474 5132
rect 282453 5130 282519 5133
rect 90468 5128 282519 5130
rect 90468 5072 282458 5128
rect 282514 5072 282519 5128
rect 90468 5070 282519 5072
rect 90468 5068 90474 5070
rect 282453 5067 282519 5070
rect 16021 4994 16087 4997
rect 502190 4994 502196 4996
rect 16021 4992 502196 4994
rect 16021 4936 16026 4992
rect 16082 4936 502196 4992
rect 16021 4934 502196 4936
rect 16021 4931 16087 4934
rect 502190 4932 502196 4934
rect 502260 4932 502266 4996
rect 5257 4858 5323 4861
rect 503294 4858 503300 4860
rect 5257 4856 503300 4858
rect 5257 4800 5262 4856
rect 5318 4800 503300 4856
rect 5257 4798 503300 4800
rect 5257 4795 5323 4798
rect 503294 4796 503300 4798
rect 503364 4796 503370 4860
rect 86125 4724 86191 4725
rect 86125 4722 86172 4724
rect 86080 4720 86172 4722
rect 86080 4664 86130 4720
rect 86080 4662 86172 4664
rect 86125 4660 86172 4662
rect 86236 4660 86242 4724
rect 86125 4659 86191 4660
rect 164366 4388 164372 4452
rect 164436 4450 164442 4452
rect 169150 4450 169156 4452
rect 164436 4390 169156 4450
rect 164436 4388 164442 4390
rect 169150 4388 169156 4390
rect 169220 4388 169226 4452
rect 172462 4388 172468 4452
rect 172532 4450 172538 4452
rect 182030 4450 182036 4452
rect 172532 4390 182036 4450
rect 172532 4388 172538 4390
rect 182030 4388 182036 4390
rect 182100 4388 182106 4452
rect 329230 4388 329236 4452
rect 329300 4450 329306 4452
rect 337878 4450 337884 4452
rect 329300 4390 337884 4450
rect 329300 4388 329306 4390
rect 337878 4388 337884 4390
rect 337948 4388 337954 4452
rect 396022 4388 396028 4452
rect 396092 4450 396098 4452
rect 405590 4450 405596 4452
rect 396092 4390 405596 4450
rect 396092 4388 396098 4390
rect 405590 4388 405596 4390
rect 405660 4388 405666 4452
rect 415710 4388 415716 4452
rect 415780 4450 415786 4452
rect 424910 4450 424916 4452
rect 415780 4390 424916 4450
rect 415780 4388 415786 4390
rect 424910 4388 424916 4390
rect 424980 4388 424986 4452
rect 434662 4388 434668 4452
rect 434732 4450 434738 4452
rect 443310 4450 443316 4452
rect 434732 4390 443316 4450
rect 434732 4388 434738 4390
rect 443310 4388 443316 4390
rect 443380 4388 443386 4452
rect 444414 4252 444420 4316
rect 444484 4314 444490 4316
rect 457478 4314 457484 4316
rect 444484 4254 457484 4314
rect 444484 4252 444490 4254
rect 457478 4252 457484 4254
rect 457548 4252 457554 4316
rect 84377 4180 84443 4181
rect 86401 4180 86467 4181
rect 84326 4178 84332 4180
rect 84286 4118 84332 4178
rect 84396 4176 84443 4180
rect 86350 4178 86356 4180
rect 84438 4120 84443 4176
rect 84326 4116 84332 4118
rect 84396 4116 84443 4120
rect 86310 4118 86356 4178
rect 86420 4176 86467 4180
rect 86462 4120 86467 4176
rect 86350 4116 86356 4118
rect 86420 4116 86467 4120
rect 84377 4115 84443 4116
rect 86401 4115 86467 4116
rect 318885 4178 318951 4181
rect 318885 4176 319178 4178
rect 318885 4120 318890 4176
rect 318946 4120 319178 4176
rect 318885 4118 319178 4120
rect 318885 4115 318951 4118
rect 70301 4042 70367 4045
rect 271505 4042 271571 4045
rect 70301 4040 271571 4042
rect 70301 3984 70306 4040
rect 70362 3984 271510 4040
rect 271566 3984 271571 4040
rect 70301 3982 271571 3984
rect 70301 3979 70367 3982
rect 271505 3979 271571 3982
rect 271689 4042 271755 4045
rect 275277 4042 275343 4045
rect 275870 4042 275876 4044
rect 271689 4040 275202 4042
rect 271689 3984 271694 4040
rect 271750 3984 275202 4040
rect 271689 3982 275202 3984
rect 271689 3979 271755 3982
rect 81433 3906 81499 3909
rect 84326 3906 84332 3908
rect 81433 3904 84332 3906
rect 81433 3848 81438 3904
rect 81494 3848 84332 3904
rect 81433 3846 84332 3848
rect 81433 3843 81499 3846
rect 84326 3844 84332 3846
rect 84396 3844 84402 3908
rect 88517 3906 88583 3909
rect 89110 3906 89116 3908
rect 88517 3904 89116 3906
rect 88517 3848 88522 3904
rect 88578 3848 89116 3904
rect 88517 3846 89116 3848
rect 88517 3843 88583 3846
rect 89110 3844 89116 3846
rect 89180 3844 89186 3908
rect 90725 3906 90791 3909
rect 89302 3904 90791 3906
rect 89302 3848 90730 3904
rect 90786 3848 90791 3904
rect 89302 3846 90791 3848
rect 79041 3770 79107 3773
rect 86350 3770 86356 3772
rect 79041 3768 86356 3770
rect 79041 3712 79046 3768
rect 79102 3712 86356 3768
rect 79041 3710 86356 3712
rect 79041 3707 79107 3710
rect 86350 3708 86356 3710
rect 86420 3708 86426 3772
rect 87086 3708 87092 3772
rect 87156 3770 87162 3772
rect 89302 3770 89362 3846
rect 90725 3843 90791 3846
rect 90909 3906 90975 3909
rect 92422 3906 92428 3908
rect 90909 3904 92428 3906
rect 90909 3848 90914 3904
rect 90970 3848 92428 3904
rect 90909 3846 92428 3848
rect 90909 3843 90975 3846
rect 92422 3844 92428 3846
rect 92492 3844 92498 3908
rect 93526 3844 93532 3908
rect 93596 3906 93602 3908
rect 263409 3906 263475 3909
rect 275142 3906 275202 3982
rect 275277 4040 275876 4042
rect 275277 3984 275282 4040
rect 275338 3984 275876 4040
rect 275277 3982 275876 3984
rect 275277 3979 275343 3982
rect 275870 3980 275876 3982
rect 275940 3980 275946 4044
rect 278865 4042 278931 4045
rect 318793 4042 318859 4045
rect 278865 4040 318859 4042
rect 278865 3984 278870 4040
rect 278926 3984 318798 4040
rect 318854 3984 318859 4040
rect 278865 3982 318859 3984
rect 319118 4042 319178 4118
rect 384982 4116 384988 4180
rect 385052 4178 385058 4180
rect 394601 4178 394667 4181
rect 385052 4176 394667 4178
rect 385052 4120 394606 4176
rect 394662 4120 394667 4176
rect 385052 4118 394667 4120
rect 385052 4116 385058 4118
rect 394601 4115 394667 4118
rect 479374 4116 479380 4180
rect 479444 4178 479450 4180
rect 485630 4178 485636 4180
rect 479444 4118 485636 4178
rect 479444 4116 479450 4118
rect 485630 4116 485636 4118
rect 485700 4116 485706 4180
rect 356789 4042 356855 4045
rect 319118 4040 356855 4042
rect 319118 3984 356794 4040
rect 356850 3984 356855 4040
rect 319118 3982 356855 3984
rect 278865 3979 278931 3982
rect 318793 3979 318859 3982
rect 356789 3979 356855 3982
rect 357249 4042 357315 4045
rect 494697 4042 494763 4045
rect 357249 4040 494763 4042
rect 357249 3984 357254 4040
rect 357310 3984 494702 4040
rect 494758 3984 494763 4040
rect 357249 3982 494763 3984
rect 357249 3979 357315 3982
rect 494697 3979 494763 3982
rect 495617 4042 495683 4045
rect 500166 4042 500172 4044
rect 495617 4040 500172 4042
rect 495617 3984 495622 4040
rect 495678 3984 500172 4040
rect 495617 3982 500172 3984
rect 495617 3979 495683 3982
rect 500166 3980 500172 3982
rect 500236 3980 500242 4044
rect 318742 3906 318748 3908
rect 93596 3904 263475 3906
rect 93596 3848 263414 3904
rect 263470 3848 263475 3904
rect 93596 3846 263475 3848
rect 93596 3844 93602 3846
rect 263409 3843 263475 3846
rect 270358 3846 275018 3906
rect 275142 3846 318748 3906
rect 115749 3770 115815 3773
rect 87156 3710 89362 3770
rect 93166 3768 115815 3770
rect 93166 3712 115754 3768
rect 115810 3712 115815 3768
rect 93166 3710 115815 3712
rect 87156 3708 87162 3710
rect 88190 3572 88196 3636
rect 88260 3634 88266 3636
rect 93166 3634 93226 3710
rect 115749 3707 115815 3710
rect 115933 3770 115999 3773
rect 116710 3770 116716 3772
rect 115933 3768 116716 3770
rect 115933 3712 115938 3768
rect 115994 3712 116716 3768
rect 115933 3710 116716 3712
rect 115933 3707 115999 3710
rect 116710 3708 116716 3710
rect 116780 3708 116786 3772
rect 116853 3770 116919 3773
rect 162117 3770 162183 3773
rect 163497 3770 163563 3773
rect 163998 3770 164004 3772
rect 116853 3768 162183 3770
rect 116853 3712 116858 3768
rect 116914 3712 162122 3768
rect 162178 3712 162183 3768
rect 116853 3710 162183 3712
rect 116853 3707 116919 3710
rect 162117 3707 162183 3710
rect 162902 3710 163146 3770
rect 88260 3574 93226 3634
rect 95141 3634 95207 3637
rect 143441 3634 143507 3637
rect 153101 3634 153167 3637
rect 162761 3634 162827 3637
rect 162902 3634 162962 3710
rect 95141 3632 125610 3634
rect 95141 3576 95146 3632
rect 95202 3576 125610 3632
rect 95141 3574 125610 3576
rect 88260 3572 88266 3574
rect 95141 3571 95207 3574
rect 82537 3498 82603 3501
rect 85573 3498 85639 3501
rect 82537 3496 85639 3498
rect 82537 3440 82542 3496
rect 82598 3440 85578 3496
rect 85634 3440 85639 3496
rect 82537 3438 85639 3440
rect 82537 3435 82603 3438
rect 85573 3435 85639 3438
rect 90725 3498 90791 3501
rect 122005 3498 122071 3501
rect 90725 3496 122071 3498
rect 90725 3440 90730 3496
rect 90786 3440 122010 3496
rect 122066 3440 122071 3496
rect 90725 3438 122071 3440
rect 90725 3435 90791 3438
rect 122005 3435 122071 3438
rect 122782 3436 122788 3500
rect 122852 3498 122858 3500
rect 123017 3498 123083 3501
rect 125550 3500 125610 3574
rect 143441 3632 143642 3634
rect 143441 3576 143446 3632
rect 143502 3576 143642 3632
rect 143441 3574 143642 3576
rect 153020 3632 153210 3634
rect 153020 3576 153106 3632
rect 153162 3576 153210 3632
rect 153020 3574 153210 3576
rect 143441 3571 143507 3574
rect 143582 3500 143642 3574
rect 153101 3571 153210 3574
rect 162761 3632 162962 3634
rect 162761 3576 162766 3632
rect 162822 3576 162962 3632
rect 162761 3574 162962 3576
rect 163086 3634 163146 3710
rect 163497 3768 164004 3770
rect 163497 3712 163502 3768
rect 163558 3712 164004 3768
rect 163497 3710 164004 3712
rect 163497 3707 163563 3710
rect 163998 3708 164004 3710
rect 164068 3708 164074 3772
rect 164693 3770 164759 3773
rect 206921 3770 206987 3773
rect 164693 3768 206987 3770
rect 164693 3712 164698 3768
rect 164754 3712 206926 3768
rect 206982 3712 206987 3768
rect 164693 3710 206987 3712
rect 164693 3707 164759 3710
rect 206921 3707 206987 3710
rect 207054 3708 207060 3772
rect 207124 3770 207130 3772
rect 207473 3770 207539 3773
rect 207124 3768 207539 3770
rect 207124 3712 207478 3768
rect 207534 3712 207539 3768
rect 207124 3710 207539 3712
rect 207124 3708 207130 3710
rect 207473 3707 207539 3710
rect 218094 3708 218100 3772
rect 218164 3770 218170 3772
rect 219341 3770 219407 3773
rect 218164 3768 219407 3770
rect 218164 3712 219346 3768
rect 219402 3712 219407 3768
rect 218164 3710 219407 3712
rect 218164 3708 218170 3710
rect 219341 3707 219407 3710
rect 220077 3770 220143 3773
rect 257429 3770 257495 3773
rect 220077 3768 257495 3770
rect 220077 3712 220082 3768
rect 220138 3712 257434 3768
rect 257490 3712 257495 3768
rect 220077 3710 257495 3712
rect 220077 3707 220143 3710
rect 257429 3707 257495 3710
rect 259821 3770 259887 3773
rect 270358 3770 270418 3846
rect 259821 3768 270418 3770
rect 259821 3712 259826 3768
rect 259882 3712 270418 3768
rect 259821 3710 270418 3712
rect 270493 3770 270559 3773
rect 271638 3770 271644 3772
rect 270493 3768 271644 3770
rect 270493 3712 270498 3768
rect 270554 3712 271644 3768
rect 270493 3710 271644 3712
rect 259821 3707 259887 3710
rect 270493 3707 270559 3710
rect 271638 3708 271644 3710
rect 271708 3708 271714 3772
rect 274958 3770 275018 3846
rect 318742 3844 318748 3846
rect 318812 3844 318818 3908
rect 319110 3844 319116 3908
rect 319180 3906 319186 3908
rect 356973 3906 357039 3909
rect 319180 3904 357039 3906
rect 319180 3848 356978 3904
rect 357034 3848 357039 3904
rect 319180 3846 357039 3848
rect 319180 3844 319186 3846
rect 356973 3843 357039 3846
rect 357249 3906 357315 3909
rect 495382 3906 495388 3908
rect 357249 3904 495388 3906
rect 357249 3848 357254 3904
rect 357310 3848 495388 3904
rect 357249 3846 495388 3848
rect 357249 3843 357315 3846
rect 495382 3844 495388 3846
rect 495452 3844 495458 3908
rect 495525 3906 495591 3909
rect 502006 3906 502012 3908
rect 495525 3904 502012 3906
rect 495525 3848 495530 3904
rect 495586 3848 502012 3904
rect 495525 3846 502012 3848
rect 495525 3843 495591 3846
rect 502006 3844 502012 3846
rect 502076 3844 502082 3908
rect 318742 3770 318748 3772
rect 274958 3710 318748 3770
rect 318742 3708 318748 3710
rect 318812 3708 318818 3772
rect 319253 3770 319319 3773
rect 320030 3770 320036 3772
rect 319253 3768 320036 3770
rect 319253 3712 319258 3768
rect 319314 3712 320036 3768
rect 319253 3710 320036 3712
rect 319253 3707 319319 3710
rect 320030 3708 320036 3710
rect 320100 3708 320106 3772
rect 342294 3708 342300 3772
rect 342364 3770 342370 3772
rect 343081 3770 343147 3773
rect 342364 3768 343147 3770
rect 342364 3712 343086 3768
rect 343142 3712 343147 3768
rect 342364 3710 343147 3712
rect 342364 3708 342370 3710
rect 343081 3707 343147 3710
rect 351821 3770 351887 3773
rect 357382 3770 357388 3772
rect 351821 3768 357388 3770
rect 351821 3712 351826 3768
rect 351882 3712 357388 3768
rect 351821 3710 357388 3712
rect 351821 3707 351887 3710
rect 357382 3708 357388 3710
rect 357452 3708 357458 3772
rect 365662 3708 365668 3772
rect 365732 3770 365738 3772
rect 394601 3770 394667 3773
rect 396022 3770 396028 3772
rect 365732 3710 375298 3770
rect 365732 3708 365738 3710
rect 182081 3634 182147 3637
rect 241513 3634 241579 3637
rect 163086 3574 172530 3634
rect 162761 3571 162827 3574
rect 122852 3496 123083 3498
rect 122852 3440 123022 3496
rect 123078 3440 123083 3496
rect 122852 3438 123083 3440
rect 122852 3436 122858 3438
rect 123017 3435 123083 3438
rect 125542 3436 125548 3500
rect 125612 3436 125618 3500
rect 125726 3436 125732 3500
rect 125796 3498 125802 3500
rect 133822 3498 133828 3500
rect 125796 3438 133828 3498
rect 125796 3436 125802 3438
rect 133822 3436 133828 3438
rect 133892 3436 133898 3500
rect 143574 3436 143580 3500
rect 143644 3436 143650 3500
rect 148041 3498 148107 3501
rect 153150 3500 153210 3571
rect 148174 3498 148180 3500
rect 148041 3496 148180 3498
rect 148041 3440 148046 3496
rect 148102 3440 148180 3496
rect 148041 3438 148180 3440
rect 148041 3435 148107 3438
rect 148174 3436 148180 3438
rect 148244 3436 148250 3500
rect 153142 3436 153148 3500
rect 153212 3436 153218 3500
rect 162117 3498 162183 3501
rect 162853 3498 162919 3501
rect 172470 3500 172530 3574
rect 182081 3632 241579 3634
rect 182081 3576 182086 3632
rect 182142 3576 241518 3632
rect 241574 3576 241579 3632
rect 182081 3574 241579 3576
rect 182081 3571 182147 3574
rect 241513 3571 241579 3574
rect 259361 3634 259427 3637
rect 288382 3634 288388 3636
rect 259361 3632 288388 3634
rect 259361 3576 259366 3632
rect 259422 3576 288388 3632
rect 259361 3574 288388 3576
rect 259361 3571 259427 3574
rect 288382 3572 288388 3574
rect 288452 3572 288458 3636
rect 298001 3634 298067 3637
rect 307702 3634 307708 3636
rect 298001 3632 307708 3634
rect 298001 3576 298006 3632
rect 298062 3576 307708 3632
rect 298001 3574 307708 3576
rect 298001 3571 298067 3574
rect 307702 3572 307708 3574
rect 307772 3572 307778 3636
rect 317270 3572 317276 3636
rect 317340 3634 317346 3636
rect 327022 3634 327028 3636
rect 317340 3574 327028 3634
rect 317340 3572 317346 3574
rect 327022 3572 327028 3574
rect 327092 3572 327098 3636
rect 332593 3634 332659 3637
rect 335353 3634 335419 3637
rect 332593 3632 335419 3634
rect 332593 3576 332598 3632
rect 332654 3576 335358 3632
rect 335414 3576 335419 3632
rect 332593 3574 335419 3576
rect 375238 3634 375298 3710
rect 394601 3768 396028 3770
rect 394601 3712 394606 3768
rect 394662 3712 396028 3768
rect 394601 3710 396028 3712
rect 394601 3707 394667 3710
rect 396022 3708 396028 3710
rect 396092 3708 396098 3772
rect 400857 3770 400923 3773
rect 405641 3770 405707 3773
rect 400857 3768 405707 3770
rect 400857 3712 400862 3768
rect 400918 3712 405646 3768
rect 405702 3712 405707 3768
rect 400857 3710 405707 3712
rect 400857 3707 400923 3710
rect 405641 3707 405707 3710
rect 442257 3770 442323 3773
rect 451457 3770 451523 3773
rect 442257 3768 451523 3770
rect 442257 3712 442262 3768
rect 442318 3712 451462 3768
rect 451518 3712 451523 3768
rect 442257 3710 451523 3712
rect 442257 3707 442323 3710
rect 451457 3707 451523 3710
rect 460974 3708 460980 3772
rect 461044 3770 461050 3772
rect 462446 3770 462452 3772
rect 461044 3710 462452 3770
rect 461044 3708 461050 3710
rect 462446 3708 462452 3710
rect 462516 3708 462522 3772
rect 463233 3770 463299 3773
rect 463550 3770 463556 3772
rect 463233 3768 463556 3770
rect 463233 3712 463238 3768
rect 463294 3712 463556 3768
rect 463233 3710 463556 3712
rect 463233 3707 463299 3710
rect 463550 3708 463556 3710
rect 463620 3708 463626 3772
rect 463693 3770 463759 3773
rect 470593 3770 470659 3773
rect 478689 3772 478755 3773
rect 478638 3770 478644 3772
rect 463693 3768 470659 3770
rect 463693 3712 463698 3768
rect 463754 3712 470598 3768
rect 470654 3712 470659 3768
rect 463693 3710 470659 3712
rect 478598 3710 478644 3770
rect 478708 3768 478755 3772
rect 478750 3712 478755 3768
rect 463693 3707 463759 3710
rect 470593 3707 470659 3710
rect 478638 3708 478644 3710
rect 478708 3708 478755 3712
rect 478689 3707 478755 3708
rect 482369 3770 482435 3773
rect 495065 3770 495131 3773
rect 482369 3768 495131 3770
rect 482369 3712 482374 3768
rect 482430 3712 495070 3768
rect 495126 3712 495131 3768
rect 482369 3710 495131 3712
rect 482369 3707 482435 3710
rect 495065 3707 495131 3710
rect 495198 3708 495204 3772
rect 495268 3770 495274 3772
rect 507710 3770 507716 3772
rect 495268 3710 507716 3770
rect 495268 3708 495274 3710
rect 507710 3708 507716 3710
rect 507780 3708 507786 3772
rect 521694 3708 521700 3772
rect 521764 3770 521770 3772
rect 531078 3770 531084 3772
rect 521764 3710 531084 3770
rect 521764 3708 521770 3710
rect 531078 3708 531084 3710
rect 531148 3708 531154 3772
rect 557942 3708 557948 3772
rect 558012 3770 558018 3772
rect 558361 3770 558427 3773
rect 558012 3768 558427 3770
rect 558012 3712 558366 3768
rect 558422 3712 558427 3768
rect 558012 3710 558427 3712
rect 558012 3708 558018 3710
rect 558361 3707 558427 3710
rect 384982 3634 384988 3636
rect 375238 3574 384988 3634
rect 332593 3571 332659 3574
rect 335353 3571 335419 3574
rect 384982 3572 384988 3574
rect 385052 3572 385058 3636
rect 425145 3634 425211 3637
rect 425462 3634 425468 3636
rect 425145 3632 425468 3634
rect 425145 3576 425150 3632
rect 425206 3576 425468 3632
rect 425145 3574 425468 3576
rect 425145 3571 425211 3574
rect 425462 3572 425468 3574
rect 425532 3572 425538 3636
rect 435817 3634 435883 3637
rect 495382 3634 495388 3636
rect 435817 3632 495388 3634
rect 435817 3576 435822 3632
rect 435878 3576 495388 3632
rect 435817 3574 495388 3576
rect 435817 3571 435883 3574
rect 495382 3572 495388 3574
rect 495452 3572 495458 3636
rect 495566 3572 495572 3636
rect 495636 3634 495642 3636
rect 500033 3634 500099 3637
rect 495636 3632 500099 3634
rect 495636 3576 500038 3632
rect 500094 3576 500099 3632
rect 495636 3574 500099 3576
rect 495636 3572 495642 3574
rect 500033 3571 500099 3574
rect 162117 3496 162919 3498
rect 162117 3440 162122 3496
rect 162178 3440 162858 3496
rect 162914 3440 162919 3496
rect 162117 3438 162919 3440
rect 162117 3435 162183 3438
rect 162853 3435 162919 3438
rect 172462 3436 172468 3500
rect 172532 3436 172538 3500
rect 175365 3498 175431 3501
rect 176510 3498 176516 3500
rect 175365 3496 176516 3498
rect 175365 3440 175370 3496
rect 175426 3440 176516 3496
rect 175365 3438 176516 3440
rect 175365 3435 175431 3438
rect 176510 3436 176516 3438
rect 176580 3436 176586 3500
rect 206921 3498 206987 3501
rect 220077 3498 220143 3501
rect 206921 3496 220143 3498
rect 206921 3440 206926 3496
rect 206982 3440 220082 3496
rect 220138 3440 220143 3496
rect 206921 3438 220143 3440
rect 206921 3435 206987 3438
rect 220077 3435 220143 3438
rect 220261 3498 220327 3501
rect 499798 3498 499804 3500
rect 220261 3496 499804 3498
rect 220261 3440 220266 3496
rect 220322 3440 499804 3496
rect 220261 3438 499804 3440
rect 220261 3435 220327 3438
rect 499798 3436 499804 3438
rect 499868 3436 499874 3500
rect 80830 3300 80836 3364
rect 80900 3362 80906 3364
rect 162853 3362 162919 3365
rect 80900 3360 162919 3362
rect 80900 3304 162858 3360
rect 162914 3304 162919 3360
rect 80900 3302 162919 3304
rect 80900 3300 80906 3302
rect 162853 3299 162919 3302
rect 163313 3362 163379 3365
rect 460841 3362 460907 3365
rect 163313 3360 460907 3362
rect 163313 3304 163318 3360
rect 163374 3304 460846 3360
rect 460902 3304 460907 3360
rect 163313 3302 460907 3304
rect 163313 3299 163379 3302
rect 460841 3299 460907 3302
rect 464429 3362 464495 3365
rect 498326 3362 498332 3364
rect 464429 3360 498332 3362
rect 464429 3304 464434 3360
rect 464490 3304 498332 3360
rect 464429 3302 498332 3304
rect 464429 3299 464495 3302
rect 498326 3300 498332 3302
rect 498396 3300 498402 3364
rect 86217 3226 86283 3229
rect 299105 3226 299171 3229
rect 86217 3224 299171 3226
rect 86217 3168 86222 3224
rect 86278 3168 299110 3224
rect 299166 3168 299171 3224
rect 86217 3166 299171 3168
rect 86217 3163 86283 3166
rect 299105 3163 299171 3166
rect 301405 3226 301471 3229
rect 495750 3226 495756 3228
rect 301405 3224 495756 3226
rect 301405 3168 301410 3224
rect 301466 3168 495756 3224
rect 301405 3166 495756 3168
rect 301405 3163 301471 3166
rect 495750 3164 495756 3166
rect 495820 3164 495826 3228
rect 499062 3226 499068 3228
rect 495942 3166 499068 3226
rect 84694 3028 84700 3092
rect 84764 3090 84770 3092
rect 107561 3090 107627 3093
rect 84764 3088 107627 3090
rect 84764 3032 107566 3088
rect 107622 3032 107627 3088
rect 84764 3030 107627 3032
rect 84764 3028 84770 3030
rect 107561 3027 107627 3030
rect 107694 3028 107700 3092
rect 107764 3090 107770 3092
rect 108757 3090 108823 3093
rect 107764 3088 108823 3090
rect 107764 3032 108762 3088
rect 108818 3032 108823 3088
rect 107764 3030 108823 3032
rect 107764 3028 107770 3030
rect 108757 3027 108823 3030
rect 108941 3090 109007 3093
rect 238385 3090 238451 3093
rect 108941 3088 238451 3090
rect 108941 3032 108946 3088
rect 109002 3032 238390 3088
rect 238446 3032 238451 3088
rect 108941 3030 238451 3032
rect 108941 3027 109007 3030
rect 238385 3027 238451 3030
rect 243486 3028 243492 3092
rect 243556 3090 243562 3092
rect 243556 3030 244474 3090
rect 243556 3028 243562 3030
rect 94497 2954 94563 2957
rect 101254 2954 101260 2956
rect 94497 2952 101260 2954
rect 94497 2896 94502 2952
rect 94558 2896 101260 2952
rect 94497 2894 101260 2896
rect 94497 2891 94563 2894
rect 101254 2892 101260 2894
rect 101324 2892 101330 2956
rect 114737 2954 114803 2957
rect 114870 2954 114876 2956
rect 114737 2952 114876 2954
rect 114737 2896 114742 2952
rect 114798 2896 114876 2952
rect 114737 2894 114876 2896
rect 114737 2891 114803 2894
rect 114870 2892 114876 2894
rect 114940 2892 114946 2956
rect 122005 2954 122071 2957
rect 125409 2954 125475 2957
rect 122005 2952 125475 2954
rect 122005 2896 122010 2952
rect 122066 2896 125414 2952
rect 125470 2896 125475 2952
rect 122005 2894 125475 2896
rect 122005 2891 122071 2894
rect 125409 2891 125475 2894
rect 133822 2892 133828 2956
rect 133892 2954 133898 2956
rect 143441 2954 143507 2957
rect 153101 2956 153167 2957
rect 133892 2952 143507 2954
rect 133892 2896 143446 2952
rect 143502 2896 143507 2952
rect 133892 2894 143507 2896
rect 133892 2892 133898 2894
rect 143441 2891 143507 2894
rect 143574 2892 143580 2956
rect 143644 2954 143650 2956
rect 153101 2954 153148 2956
rect 143644 2952 153148 2954
rect 153212 2954 153218 2956
rect 162761 2954 162827 2957
rect 153212 2952 162827 2954
rect 143644 2896 153106 2952
rect 153212 2896 162766 2952
rect 162822 2896 162827 2952
rect 143644 2894 153148 2896
rect 143644 2892 143650 2894
rect 153101 2892 153148 2894
rect 153212 2894 162827 2896
rect 153212 2892 153218 2894
rect 153101 2891 153167 2892
rect 162761 2891 162827 2894
rect 172462 2892 172468 2956
rect 172532 2954 172538 2956
rect 182081 2954 182147 2957
rect 172532 2952 182147 2954
rect 172532 2896 182086 2952
rect 182142 2896 182147 2952
rect 172532 2894 182147 2896
rect 172532 2892 172538 2894
rect 182081 2891 182147 2894
rect 218145 2954 218211 2957
rect 220261 2954 220327 2957
rect 218145 2952 220327 2954
rect 218145 2896 218150 2952
rect 218206 2896 220266 2952
rect 220322 2896 220327 2952
rect 218145 2894 220327 2896
rect 244414 2954 244474 3030
rect 252502 3028 252508 3092
rect 252572 3090 252578 3092
rect 253841 3090 253907 3093
rect 267590 3090 267596 3092
rect 252572 3088 253907 3090
rect 252572 3032 253846 3088
rect 253902 3032 253907 3088
rect 252572 3030 253907 3032
rect 252572 3028 252578 3030
rect 253841 3027 253907 3030
rect 253982 3030 267596 3090
rect 253982 2954 254042 3030
rect 267590 3028 267596 3030
rect 267660 3028 267666 3092
rect 271505 3090 271571 3093
rect 280061 3090 280127 3093
rect 271505 3088 280127 3090
rect 271505 3032 271510 3088
rect 271566 3032 280066 3088
rect 280122 3032 280127 3088
rect 271505 3030 280127 3032
rect 271505 3027 271571 3030
rect 280061 3027 280127 3030
rect 288382 3028 288388 3092
rect 288452 3090 288458 3092
rect 298001 3090 298067 3093
rect 288452 3088 298067 3090
rect 288452 3032 298006 3088
rect 298062 3032 298067 3088
rect 288452 3030 298067 3032
rect 288452 3028 288458 3030
rect 298001 3027 298067 3030
rect 301998 3028 302004 3092
rect 302068 3090 302074 3092
rect 306230 3090 306236 3092
rect 302068 3030 306236 3090
rect 302068 3028 302074 3030
rect 306230 3028 306236 3030
rect 306300 3028 306306 3092
rect 315982 3028 315988 3092
rect 316052 3090 316058 3092
rect 325550 3090 325556 3092
rect 316052 3030 325556 3090
rect 316052 3028 316058 3030
rect 325550 3028 325556 3030
rect 325620 3028 325626 3092
rect 332593 3090 332659 3093
rect 325696 3088 332659 3090
rect 325696 3032 332598 3088
rect 332654 3032 332659 3088
rect 325696 3030 332659 3032
rect 244414 2894 254042 2954
rect 218145 2891 218211 2894
rect 220261 2891 220327 2894
rect 264462 2892 264468 2956
rect 264532 2954 264538 2956
rect 268878 2954 268884 2956
rect 264532 2894 268884 2954
rect 264532 2892 264538 2894
rect 268878 2892 268884 2894
rect 268948 2892 268954 2956
rect 307702 2892 307708 2956
rect 307772 2954 307778 2956
rect 317270 2954 317276 2956
rect 307772 2894 317276 2954
rect 307772 2892 307778 2894
rect 317270 2892 317276 2894
rect 317340 2892 317346 2956
rect 318742 2892 318748 2956
rect 318812 2954 318818 2956
rect 325696 2954 325756 3030
rect 332593 3027 332659 3030
rect 335353 3090 335419 3093
rect 351821 3090 351887 3093
rect 335353 3088 351887 3090
rect 335353 3032 335358 3088
rect 335414 3032 351826 3088
rect 351882 3032 351887 3088
rect 335353 3030 351887 3032
rect 335353 3027 335419 3030
rect 351821 3027 351887 3030
rect 357382 3028 357388 3092
rect 357452 3090 357458 3092
rect 365662 3090 365668 3092
rect 357452 3030 365668 3090
rect 357452 3028 357458 3030
rect 365662 3028 365668 3030
rect 365732 3028 365738 3092
rect 378542 3028 378548 3092
rect 378612 3090 378618 3092
rect 379646 3090 379652 3092
rect 378612 3030 379652 3090
rect 378612 3028 378618 3030
rect 379646 3028 379652 3030
rect 379716 3028 379722 3092
rect 396022 3028 396028 3092
rect 396092 3090 396098 3092
rect 400857 3090 400923 3093
rect 396092 3088 400923 3090
rect 396092 3032 400862 3088
rect 400918 3032 400923 3088
rect 396092 3030 400923 3032
rect 396092 3028 396098 3030
rect 400857 3027 400923 3030
rect 417550 3028 417556 3092
rect 417620 3090 417626 3092
rect 419206 3090 419212 3092
rect 417620 3030 419212 3090
rect 417620 3028 417626 3030
rect 419206 3028 419212 3030
rect 419276 3028 419282 3092
rect 436134 3028 436140 3092
rect 436204 3090 436210 3092
rect 437422 3090 437428 3092
rect 436204 3030 437428 3090
rect 436204 3028 436210 3030
rect 437422 3028 437428 3030
rect 437492 3028 437498 3092
rect 442993 3090 443059 3093
rect 495942 3090 496002 3166
rect 499062 3164 499068 3166
rect 499132 3164 499138 3228
rect 442993 3088 496002 3090
rect 442993 3032 442998 3088
rect 443054 3032 496002 3088
rect 442993 3030 496002 3032
rect 442993 3027 443059 3030
rect 496118 3028 496124 3092
rect 496188 3090 496194 3092
rect 501638 3090 501644 3092
rect 496188 3030 501644 3090
rect 496188 3028 496194 3030
rect 501638 3028 501644 3030
rect 501708 3028 501714 3092
rect 513966 3028 513972 3092
rect 514036 3090 514042 3092
rect 520038 3090 520044 3092
rect 514036 3030 520044 3090
rect 514036 3028 514042 3030
rect 520038 3028 520044 3030
rect 520108 3028 520114 3092
rect 318812 2894 325756 2954
rect 318812 2892 318818 2894
rect 327022 2892 327028 2956
rect 327092 2954 327098 2956
rect 332409 2954 332475 2957
rect 327092 2952 332475 2954
rect 327092 2896 332414 2952
rect 332470 2896 332475 2952
rect 327092 2894 332475 2896
rect 327092 2892 327098 2894
rect 332409 2891 332475 2894
rect 335302 2892 335308 2956
rect 335372 2954 335378 2956
rect 340822 2954 340828 2956
rect 335372 2894 340828 2954
rect 335372 2892 335378 2894
rect 340822 2892 340828 2894
rect 340892 2892 340898 2956
rect 425053 2954 425119 2957
rect 442257 2954 442323 2957
rect 425053 2952 442323 2954
rect 425053 2896 425058 2952
rect 425114 2896 442262 2952
rect 442318 2896 442323 2952
rect 425053 2894 442323 2896
rect 425053 2891 425119 2894
rect 442257 2891 442323 2894
rect 459645 2954 459711 2957
rect 506422 2954 506428 2956
rect 459645 2952 506428 2954
rect 459645 2896 459650 2952
rect 459706 2896 506428 2952
rect 459645 2894 506428 2896
rect 459645 2891 459711 2894
rect 506422 2892 506428 2894
rect 506492 2892 506498 2956
rect 99373 2818 99439 2821
rect 108941 2818 109007 2821
rect 99373 2816 109007 2818
rect 99373 2760 99378 2816
rect 99434 2760 108946 2816
rect 109002 2760 109007 2816
rect 99373 2758 109007 2760
rect 99373 2755 99439 2758
rect 108941 2755 109007 2758
rect 118693 2818 118759 2821
rect 122925 2818 122991 2821
rect 118693 2816 122991 2818
rect 118693 2760 118698 2816
rect 118754 2760 122930 2816
rect 122986 2760 122991 2816
rect 118693 2758 122991 2760
rect 118693 2755 118759 2758
rect 122925 2755 122991 2758
rect 241513 2818 241579 2821
rect 259361 2818 259427 2821
rect 241513 2816 259427 2818
rect 241513 2760 241518 2816
rect 241574 2760 259366 2816
rect 259422 2760 259427 2816
rect 241513 2758 259427 2760
rect 241513 2755 241579 2758
rect 259361 2755 259427 2758
rect 451457 2818 451523 2821
rect 463693 2818 463759 2821
rect 451457 2816 463759 2818
rect 451457 2760 451462 2816
rect 451518 2760 463698 2816
rect 463754 2760 463759 2816
rect 451457 2758 463759 2760
rect 451457 2755 451523 2758
rect 463693 2755 463759 2758
rect 470593 2818 470659 2821
rect 482369 2818 482435 2821
rect 470593 2816 478522 2818
rect 470593 2760 470598 2816
rect 470654 2760 478522 2816
rect 470593 2758 478522 2760
rect 470593 2755 470659 2758
rect 451590 2620 451596 2684
rect 451660 2682 451666 2684
rect 461342 2682 461348 2684
rect 451660 2622 461348 2682
rect 451660 2620 451666 2622
rect 461342 2620 461348 2622
rect 461412 2620 461418 2684
rect 478462 2682 478522 2758
rect 479014 2816 482435 2818
rect 479014 2760 482374 2816
rect 482430 2760 482435 2816
rect 479014 2758 482435 2760
rect 479014 2682 479074 2758
rect 482369 2755 482435 2758
rect 486550 2756 486556 2820
rect 486620 2818 486626 2820
rect 486969 2818 487035 2821
rect 486620 2816 487035 2818
rect 486620 2760 486974 2816
rect 487030 2760 487035 2816
rect 486620 2758 487035 2760
rect 486620 2756 486626 2758
rect 486969 2755 487035 2758
rect 490557 2818 490623 2821
rect 507853 2818 507919 2821
rect 490557 2816 507919 2818
rect 490557 2760 490562 2816
rect 490618 2760 507858 2816
rect 507914 2760 507919 2816
rect 490557 2758 507919 2760
rect 490557 2755 490623 2758
rect 507853 2755 507919 2758
rect 478462 2622 479074 2682
rect 470542 2484 470548 2548
rect 470612 2546 470618 2548
rect 479374 2546 479380 2548
rect 470612 2486 479380 2546
rect 470612 2484 470618 2486
rect 479374 2484 479380 2486
rect 479444 2484 479450 2548
<< via3 >>
rect 92244 700708 92308 700772
rect 89484 700572 89548 700636
rect 93348 700436 93412 700500
rect 91876 700300 91940 700364
rect 90220 699756 90284 699820
rect 505692 696900 505756 696964
rect 89484 695464 89548 695468
rect 89484 695408 89534 695464
rect 89534 695408 89548 695464
rect 89484 695404 89548 695408
rect 89852 689284 89916 689348
rect 89484 674792 89548 674796
rect 89484 674736 89534 674792
rect 89534 674736 89548 674792
rect 89484 674732 89548 674736
rect 89484 665272 89548 665276
rect 89484 665216 89534 665272
rect 89534 665216 89548 665272
rect 89484 665212 89548 665216
rect 89484 655480 89548 655484
rect 89484 655424 89534 655480
rect 89534 655424 89548 655480
rect 89484 655420 89548 655424
rect 89484 645960 89548 645964
rect 89484 645904 89534 645960
rect 89534 645904 89548 645960
rect 89484 645900 89548 645904
rect 89484 636168 89548 636172
rect 89484 636112 89534 636168
rect 89534 636112 89548 636168
rect 89484 636108 89548 636112
rect 89484 626648 89548 626652
rect 89484 626592 89534 626648
rect 89534 626592 89548 626648
rect 89484 626588 89548 626592
rect 89300 626452 89364 626516
rect 89484 626452 89548 626516
rect 89484 596184 89548 596188
rect 89484 596128 89498 596184
rect 89498 596128 89548 596184
rect 89484 596124 89548 596128
rect 87644 585652 87708 585716
rect 89668 584972 89732 585036
rect 88196 584836 88260 584900
rect 172468 584836 172532 584900
rect 91692 584700 91756 584764
rect 172652 584700 172716 584764
rect 501644 584836 501708 584900
rect 506244 584700 506308 584764
rect 88380 584564 88444 584628
rect 97764 584428 97828 584492
rect 233924 584428 233988 584492
rect 87276 584292 87340 584356
rect 88564 584156 88628 584220
rect 92612 584020 92676 584084
rect 84516 583884 84580 583948
rect 92060 583808 92124 583812
rect 92060 583752 92110 583808
rect 92110 583752 92124 583808
rect 92060 583748 92124 583752
rect 93532 583748 93596 583812
rect 233188 583748 233252 583812
rect 298140 583748 298204 583812
rect 499068 583748 499132 583812
rect 499436 583884 499500 583948
rect 509372 583748 509436 583812
rect 84700 582932 84764 582996
rect 500356 582932 500420 582996
rect 89484 582796 89548 582860
rect 106044 582796 106108 582860
rect 501276 582660 501340 582724
rect 506060 582524 506124 582588
rect 86724 582388 86788 582452
rect 89116 582116 89180 582180
rect 113772 582252 113836 582316
rect 505876 582388 505940 582452
rect 162348 582252 162412 582316
rect 181668 582252 181732 582316
rect 190684 582252 190748 582316
rect 200988 582252 201052 582316
rect 316540 582252 316604 582316
rect 326476 582252 326540 582316
rect 412772 582252 412836 582316
rect 423076 582252 423140 582316
rect 431908 582252 431972 582316
rect 442212 582252 442276 582316
rect 451964 582252 452028 582316
rect 461348 582252 461412 582316
rect 470548 582252 470612 582316
rect 480852 582252 480916 582316
rect 489868 582252 489932 582316
rect 510660 582252 510724 582316
rect 210372 582116 210436 582180
rect 260788 582116 260852 582180
rect 277532 582116 277596 582180
rect 287836 582116 287900 582180
rect 297220 582116 297284 582180
rect 306604 582116 306668 582180
rect 316724 582116 316788 582180
rect 326292 582116 326356 582180
rect 393452 582116 393516 582180
rect 403756 582116 403820 582180
rect 412588 582116 412652 582180
rect 422892 582116 422956 582180
rect 491708 582116 491772 582180
rect 85252 581980 85316 582044
rect 89852 581980 89916 582044
rect 151676 581980 151740 582044
rect 156460 581980 156524 582044
rect 221228 581980 221292 582044
rect 229324 581980 229388 582044
rect 249748 581980 249812 582044
rect 268516 581980 268580 582044
rect 277716 581980 277780 582044
rect 287652 581980 287716 582044
rect 297404 581980 297468 582044
rect 306052 581980 306116 582044
rect 497412 581980 497476 582044
rect 84884 581844 84948 581908
rect 91324 581844 91388 581908
rect 91692 581844 91756 581908
rect 249012 581844 249076 581908
rect 258948 581844 259012 581908
rect 268332 581844 268396 581908
rect 498148 581844 498212 581908
rect 85620 581708 85684 581772
rect 88012 581708 88076 581772
rect 335860 581708 335924 581772
rect 350396 581708 350460 581772
rect 355364 581708 355428 581772
rect 364748 581708 364812 581772
rect 374132 581708 374196 581772
rect 384436 581708 384500 581772
rect 393268 581708 393332 581772
rect 403572 581708 403636 581772
rect 498332 581708 498396 581772
rect 86356 581572 86420 581636
rect 108988 581572 109052 581636
rect 128124 581572 128188 581636
rect 128308 581572 128372 581636
rect 137876 581572 137940 581636
rect 157196 581572 157260 581636
rect 84332 581436 84396 581500
rect 85436 581496 85500 581500
rect 85436 581440 85486 581496
rect 85486 581440 85500 581496
rect 85436 581436 85500 581440
rect 113588 581436 113652 581500
rect 123340 581436 123404 581500
rect 87460 581300 87524 581364
rect 89300 581360 89364 581364
rect 89300 581304 89314 581360
rect 89314 581304 89364 581360
rect 89300 581300 89364 581304
rect 90036 581300 90100 581364
rect 90588 581300 90652 581364
rect 91692 581360 91756 581364
rect 91692 581304 91742 581360
rect 91742 581304 91756 581360
rect 91692 581300 91756 581304
rect 92428 581300 92492 581364
rect 93164 581360 93228 581364
rect 93164 581304 93214 581360
rect 93214 581304 93228 581360
rect 93164 581300 93228 581304
rect 109356 581300 109420 581364
rect 186268 581572 186332 581636
rect 195836 581572 195900 581636
rect 191052 581436 191116 581500
rect 205588 581572 205652 581636
rect 224908 581572 224972 581636
rect 244228 581572 244292 581636
rect 260604 581572 260668 581636
rect 321876 581572 321940 581636
rect 336044 581572 336108 581636
rect 345612 581572 345676 581636
rect 346900 581632 346964 581636
rect 346900 581576 346914 581632
rect 346914 581576 346964 581632
rect 346900 581572 346964 581576
rect 351684 581632 351748 581636
rect 351684 581576 351698 581632
rect 351698 581576 351748 581632
rect 351684 581572 351748 581576
rect 355180 581572 355244 581636
rect 360148 581572 360212 581636
rect 365116 581572 365180 581636
rect 373948 581572 374012 581636
rect 384252 581572 384316 581636
rect 384804 581632 384868 581636
rect 384804 581576 384854 581632
rect 384854 581576 384868 581632
rect 384804 581572 384868 581576
rect 389772 581632 389836 581636
rect 389772 581576 389786 581632
rect 389786 581576 389836 581632
rect 389772 581572 389836 581576
rect 391796 581632 391860 581636
rect 391796 581576 391810 581632
rect 391810 581576 391860 581632
rect 391796 581572 391860 581576
rect 498700 581572 498764 581636
rect 499988 581572 500052 581636
rect 83780 581164 83844 581228
rect 94268 581164 94332 581228
rect 85804 581028 85868 581092
rect 104388 581164 104452 581228
rect 108804 581164 108868 581228
rect 118556 581164 118620 581228
rect 109356 581028 109420 581092
rect 113588 581028 113652 581092
rect 113772 581028 113836 581092
rect 137324 581164 137388 581228
rect 82308 580892 82372 580956
rect 86356 580892 86420 580956
rect 94268 580892 94332 580956
rect 104388 580892 104452 580956
rect 118556 580756 118620 580820
rect 123340 581028 123404 581092
rect 128124 581028 128188 581092
rect 128308 581028 128372 581092
rect 137508 581028 137572 581092
rect 138060 581028 138124 581092
rect 137324 580892 137388 580956
rect 151676 581164 151740 581228
rect 156092 581300 156156 581364
rect 138428 581028 138492 581092
rect 156092 581028 156156 581092
rect 156460 581164 156524 581228
rect 161428 581164 161492 581228
rect 162348 581164 162412 581228
rect 181668 581164 181732 581228
rect 186268 581164 186332 581228
rect 190500 581164 190564 581228
rect 190684 581164 190748 581228
rect 200988 581164 201052 581228
rect 205588 581164 205652 581228
rect 224908 581164 224972 581228
rect 506428 581436 506492 581500
rect 231900 581360 231964 581364
rect 231900 581304 231950 581360
rect 231950 581304 231964 581360
rect 231900 581300 231964 581304
rect 157196 581028 157260 581092
rect 210372 581028 210436 581092
rect 221228 581028 221292 581092
rect 229324 581028 229388 581092
rect 244228 581164 244292 581228
rect 249748 581164 249812 581228
rect 358676 581360 358740 581364
rect 358676 581304 358726 581360
rect 358726 581304 358740 581360
rect 260604 581164 260668 581228
rect 260788 581164 260852 581228
rect 268516 581164 268580 581228
rect 277532 581164 277596 581228
rect 287836 581164 287900 581228
rect 297220 581164 297284 581228
rect 306604 581164 306668 581228
rect 316724 581164 316788 581228
rect 326292 581164 326356 581228
rect 335860 581164 335924 581228
rect 350396 581164 350460 581228
rect 355180 581164 355244 581228
rect 358676 581300 358740 581304
rect 360148 581164 360212 581228
rect 374132 581164 374196 581228
rect 384436 581164 384500 581228
rect 393452 581164 393516 581228
rect 403756 581164 403820 581228
rect 412772 581164 412836 581228
rect 423076 581164 423140 581228
rect 432092 581164 432156 581228
rect 437428 581164 437492 581228
rect 456564 581164 456628 581228
rect 456748 581164 456812 581228
rect 470732 581164 470796 581228
rect 476068 581164 476132 581228
rect 489868 581164 489932 581228
rect 495388 581164 495452 581228
rect 499988 581164 500052 581228
rect 509188 581164 509252 581228
rect 550588 581300 550652 581364
rect 249012 581028 249076 581092
rect 258948 581028 259012 581092
rect 268332 581028 268396 581092
rect 277716 581028 277780 581092
rect 287652 581028 287716 581092
rect 297404 581028 297468 581092
rect 306052 581028 306116 581092
rect 316540 581028 316604 581092
rect 326476 581028 326540 581092
rect 336044 581028 336108 581092
rect 345612 581028 345676 581092
rect 355364 581028 355428 581092
rect 364748 581028 364812 581092
rect 373948 581028 374012 581092
rect 384252 581028 384316 581092
rect 393268 581028 393332 581092
rect 403572 581028 403636 581092
rect 412588 581028 412652 581092
rect 422892 581028 422956 581092
rect 431908 581028 431972 581092
rect 442212 581028 442276 581092
rect 451964 581028 452028 581092
rect 461348 581028 461412 581092
rect 470548 581028 470612 581092
rect 480852 581028 480916 581092
rect 489868 581028 489932 581092
rect 550588 581028 550652 581092
rect 179276 580892 179340 580956
rect 195836 580892 195900 580956
rect 389772 580892 389836 580956
rect 384804 580756 384868 580820
rect 501092 580756 501156 580820
rect 161428 580620 161492 580684
rect 169708 580620 169772 580684
rect 391796 580620 391860 580684
rect 99972 580484 100036 580548
rect 113772 580484 113836 580548
rect 114508 580484 114572 580548
rect 123708 580484 123772 580548
rect 124260 580484 124324 580548
rect 137140 580484 137204 580548
rect 142108 580484 142172 580548
rect 151492 580484 151556 580548
rect 151860 580484 151924 580548
rect 161244 580484 161308 580548
rect 166212 580484 166276 580548
rect 167684 580484 167748 580548
rect 197308 580484 197372 580548
rect 206876 580484 206940 580548
rect 216628 580484 216692 580548
rect 226196 580484 226260 580548
rect 358676 580484 358740 580548
rect 502012 580484 502076 580548
rect 86908 580348 86972 580412
rect 231900 580348 231964 580412
rect 245700 580348 245764 580412
rect 254900 580348 254964 580412
rect 260972 580348 261036 580412
rect 270356 580348 270420 580412
rect 272564 580348 272628 580412
rect 273852 580348 273916 580412
rect 282316 580348 282380 580412
rect 283420 580348 283484 580412
rect 291884 580348 291948 580412
rect 293172 580348 293236 580412
rect 330708 580348 330772 580412
rect 331812 580348 331876 580412
rect 338068 580348 338132 580412
rect 341380 580348 341444 580412
rect 346900 580348 346964 580412
rect 91140 580212 91204 580276
rect 321876 580212 321940 580276
rect 351684 580212 351748 580276
rect 91508 580076 91572 580140
rect 93716 580076 93780 580140
rect 169708 580076 169772 580140
rect 179276 580076 179340 580140
rect 318748 580076 318812 580140
rect 328316 580076 328380 580140
rect 432092 580076 432156 580140
rect 437428 580076 437492 580140
rect 456564 580076 456628 580140
rect 456748 580076 456812 580140
rect 470732 580076 470796 580140
rect 476068 580076 476132 580140
rect 491708 580076 491772 580140
rect 86724 579940 86788 580004
rect 87644 579940 87708 580004
rect 88932 579940 88996 580004
rect 94084 579940 94148 580004
rect 489868 579940 489932 580004
rect 495388 579940 495452 580004
rect 90404 579804 90468 579868
rect 92612 579804 92676 579868
rect 97764 579804 97828 579868
rect 508084 577628 508148 577692
rect 506980 575452 507044 575516
rect 501276 573684 501340 573748
rect 501276 573548 501340 573612
rect 501828 573548 501892 573612
rect 501460 572188 501524 572252
rect 501460 571916 501524 571980
rect 501828 571916 501892 571980
rect 79732 570012 79796 570076
rect 505508 570012 505572 570076
rect 510108 559948 510172 560012
rect 501460 557092 501524 557156
rect 79548 555868 79612 555932
rect 82492 551788 82556 551852
rect 79364 548796 79428 548860
rect 501460 547844 501524 547908
rect 507900 545804 507964 545868
rect 507164 545396 507228 545460
rect 81388 545260 81452 545324
rect 506796 543900 506860 543964
rect 506796 543628 506860 543692
rect 502564 542268 502628 542332
rect 82124 539548 82188 539612
rect 82630 539548 82694 539612
rect 506612 538732 506676 538796
rect 81572 538188 81636 538252
rect 502932 531388 502996 531452
rect 81204 531116 81268 531180
rect 81756 527580 81820 527644
rect 82492 523772 82556 523836
rect 501644 520100 501708 520164
rect 501644 519556 501708 519620
rect 82492 519284 82556 519348
rect 82492 519012 82556 519076
rect 82492 518740 82556 518804
rect 501276 517244 501340 517308
rect 502012 517244 502076 517308
rect 502196 517244 502260 517308
rect 501276 513708 501340 513772
rect 501276 511940 501340 512004
rect 502012 511940 502076 512004
rect 77156 510172 77220 510236
rect 82308 509552 82372 509556
rect 82308 509496 82358 509552
rect 82358 509496 82372 509552
rect 82308 509492 82372 509496
rect 504220 507180 504284 507244
rect 501276 506908 501340 506972
rect 501828 506772 501892 506836
rect 502196 506772 502260 506836
rect 82492 505744 82556 505748
rect 82492 505688 82542 505744
rect 82542 505688 82556 505744
rect 82492 505684 82556 505688
rect 502380 503644 502444 503708
rect 82308 500848 82372 500852
rect 82308 500792 82358 500848
rect 82358 500792 82372 500848
rect 82308 500788 82372 500792
rect 501828 500788 501892 500852
rect 82308 498068 82372 498132
rect 82308 497176 82372 497180
rect 82308 497120 82358 497176
rect 82358 497120 82372 497176
rect 82308 497116 82372 497120
rect 82124 495756 82188 495820
rect 501828 493308 501892 493372
rect 506796 492628 506860 492692
rect 506980 492628 507044 492692
rect 81940 491948 82004 492012
rect 82492 486160 82556 486164
rect 82492 486104 82542 486160
rect 82542 486104 82556 486160
rect 82492 486100 82556 486104
rect 508268 485964 508332 486028
rect 82492 484876 82556 484940
rect 82492 481204 82556 481268
rect 82492 481128 82556 481132
rect 82492 481072 82542 481128
rect 82542 481072 82556 481128
rect 82492 481068 82556 481072
rect 501828 478620 501892 478684
rect 502012 478620 502076 478684
rect 82492 475824 82556 475828
rect 82492 475768 82542 475824
rect 82542 475768 82556 475824
rect 82492 475764 82556 475768
rect 503668 475356 503732 475420
rect 501276 474812 501340 474876
rect 82492 474192 82556 474196
rect 82492 474136 82506 474192
rect 82506 474136 82556 474192
rect 82492 474132 82556 474136
rect 82492 473588 82556 473652
rect 82492 473512 82556 473516
rect 82492 473456 82542 473512
rect 82542 473456 82556 473512
rect 82492 473452 82556 473456
rect 82492 471064 82556 471068
rect 82492 471008 82542 471064
rect 82542 471008 82556 471064
rect 82492 471004 82556 471008
rect 509740 467876 509804 467940
rect 82492 466168 82556 466172
rect 82492 466112 82506 466168
rect 82506 466112 82556 466168
rect 82492 466108 82556 466112
rect 506796 464748 506860 464812
rect 501460 464476 501524 464540
rect 502196 464476 502260 464540
rect 501644 464340 501708 464404
rect 501460 464204 501524 464268
rect 502748 461212 502812 461276
rect 82492 458008 82556 458012
rect 82492 457952 82542 458008
rect 82542 457952 82556 458008
rect 82492 457948 82556 457952
rect 82308 456860 82372 456924
rect 101628 456512 101692 456516
rect 101628 456456 101642 456512
rect 101642 456456 101692 456512
rect 101628 456452 101692 456456
rect 501644 454820 501708 454884
rect 502012 454744 502076 454748
rect 502012 454688 502062 454744
rect 502062 454688 502076 454744
rect 502012 454684 502076 454688
rect 3924 452372 3988 452436
rect 101444 451888 101508 451892
rect 101444 451832 101494 451888
rect 101494 451832 101508 451888
rect 101444 451828 101508 451832
rect 503668 450604 503732 450668
rect 502196 448972 502260 449036
rect 504588 447068 504652 447132
rect 507164 444484 507228 444548
rect 507164 444348 507228 444412
rect 501460 443260 501524 443324
rect 501276 442444 501340 442508
rect 501460 442444 501524 442508
rect 501460 442172 501524 442236
rect 501276 439724 501340 439788
rect 82492 438968 82556 438972
rect 82492 438912 82542 438968
rect 82542 438912 82556 438968
rect 82492 438908 82556 438912
rect 501460 438092 501524 438156
rect 502012 438092 502076 438156
rect 82492 435432 82556 435436
rect 82492 435376 82542 435432
rect 82542 435376 82556 435432
rect 82492 435372 82556 435376
rect 506980 434616 507044 434620
rect 506980 434560 507030 434616
rect 507030 434560 507044 434616
rect 506980 434556 507044 434560
rect 79180 432652 79244 432716
rect 82492 431216 82556 431220
rect 82492 431160 82542 431216
rect 82542 431160 82556 431216
rect 82492 431156 82556 431160
rect 504220 427892 504284 427956
rect 501276 427756 501340 427820
rect 504220 427620 504284 427684
rect 506796 425444 506860 425508
rect 506980 425232 507044 425236
rect 506980 425176 507030 425232
rect 507030 425176 507044 425232
rect 506980 425172 507044 425176
rect 507164 425172 507228 425236
rect 504404 425036 504468 425100
rect 506796 425036 506860 425100
rect 507164 425036 507228 425100
rect 502012 423812 502076 423876
rect 501828 423676 501892 423740
rect 501828 423404 501892 423468
rect 507716 422588 507780 422652
rect 78996 422044 79060 422108
rect 501276 418236 501340 418300
rect 502012 414080 502076 414084
rect 502012 414024 502062 414080
rect 502062 414024 502076 414080
rect 502012 414020 502076 414024
rect 502196 413748 502260 413812
rect 501276 411436 501340 411500
rect 501276 409940 501340 410004
rect 504036 408580 504100 408644
rect 504404 408580 504468 408644
rect 503852 408444 503916 408508
rect 82492 406464 82556 406468
rect 82492 406408 82542 406464
rect 82542 406408 82556 406464
rect 82492 406404 82556 406408
rect 501828 405724 501892 405788
rect 501828 405588 501892 405652
rect 506980 405648 507044 405652
rect 506980 405592 507030 405648
rect 507030 405592 507044 405648
rect 506980 405588 507044 405592
rect 501460 403684 501524 403748
rect 82492 401568 82556 401572
rect 82492 401512 82542 401568
rect 82542 401512 82556 401568
rect 82492 401508 82556 401512
rect 501828 400828 501892 400892
rect 502196 400828 502260 400892
rect 501828 400692 501892 400756
rect 82492 400148 82556 400212
rect 504036 398788 504100 398852
rect 502012 398712 502076 398716
rect 502012 398656 502062 398712
rect 502062 398656 502076 398712
rect 502012 398652 502076 398656
rect 504404 398652 504468 398716
rect 82492 396128 82556 396132
rect 82492 396072 82506 396128
rect 82506 396072 82556 396128
rect 82492 396068 82556 396072
rect 506980 396128 507044 396132
rect 506980 396072 507030 396128
rect 507030 396072 507044 396128
rect 506980 396068 507044 396072
rect 502196 394632 502260 394636
rect 502196 394576 502246 394632
rect 502246 394576 502260 394632
rect 502196 394572 502260 394576
rect 506980 394632 507044 394636
rect 506980 394576 507030 394632
rect 507030 394576 507044 394632
rect 506980 394572 507044 394576
rect 503300 394300 503364 394364
rect 80836 394028 80900 394092
rect 82308 394028 82372 394092
rect 80836 393076 80900 393140
rect 501644 391852 501708 391916
rect 501828 391716 501892 391780
rect 82492 391172 82556 391236
rect 503300 388316 503364 388380
rect 504036 387228 504100 387292
rect 502196 387152 502260 387156
rect 502196 387096 502246 387152
rect 502246 387096 502260 387152
rect 502196 387092 502260 387096
rect 506980 387152 507044 387156
rect 506980 387096 507030 387152
rect 507030 387096 507044 387152
rect 506980 387092 507044 387096
rect 80836 386956 80900 387020
rect 82492 385792 82556 385796
rect 82492 385736 82542 385792
rect 82542 385736 82556 385792
rect 82492 385732 82556 385736
rect 80836 385596 80900 385660
rect 82308 385656 82372 385660
rect 82308 385600 82358 385656
rect 82358 385600 82372 385656
rect 82308 385596 82372 385600
rect 501460 385052 501524 385116
rect 502012 385052 502076 385116
rect 78812 383420 78876 383484
rect 503300 382468 503364 382532
rect 507532 382468 507596 382532
rect 78628 376348 78692 376412
rect 82492 371920 82556 371924
rect 82492 371864 82506 371920
rect 82506 371864 82556 371920
rect 82492 371860 82556 371864
rect 82308 369064 82372 369068
rect 82308 369008 82358 369064
rect 82358 369008 82372 369064
rect 82308 369004 82372 369008
rect 82308 368868 82372 368932
rect 82492 368732 82556 368796
rect 82492 368112 82556 368116
rect 82492 368056 82506 368112
rect 82506 368056 82556 368112
rect 82492 368052 82556 368056
rect 82492 364848 82556 364852
rect 82492 364792 82506 364848
rect 82506 364792 82556 364848
rect 82492 364788 82556 364792
rect 82492 364652 82556 364716
rect 82492 362884 82556 362948
rect 82492 362748 82556 362812
rect 82308 360224 82372 360228
rect 82308 360168 82358 360224
rect 82358 360168 82372 360224
rect 82308 360164 82372 360168
rect 82630 360088 82694 360092
rect 82630 360032 82634 360088
rect 82634 360032 82690 360088
rect 82690 360032 82694 360088
rect 82630 360028 82694 360032
rect 82630 359348 82694 359412
rect 501460 358532 501524 358596
rect 502012 358532 502076 358596
rect 82630 358048 82694 358052
rect 82630 357992 82634 358048
rect 82634 357992 82690 358048
rect 82690 357992 82694 358048
rect 82630 357988 82694 357992
rect 503116 355676 503180 355740
rect 501276 351596 501340 351660
rect 501460 350508 501524 350572
rect 501460 349828 501524 349892
rect 504588 349828 504652 349892
rect 504036 349556 504100 349620
rect 504588 349556 504652 349620
rect 504404 347652 504468 347716
rect 82492 347032 82556 347036
rect 82492 346976 82542 347032
rect 82542 346976 82556 347032
rect 82492 346972 82556 346976
rect 501460 346428 501524 346492
rect 501460 346292 501524 346356
rect 506980 345068 507044 345132
rect 507348 345068 507412 345132
rect 502196 344992 502260 344996
rect 502196 344936 502210 344992
rect 502210 344936 502260 344992
rect 502196 344932 502260 344936
rect 501276 344796 501340 344860
rect 501460 344252 501524 344316
rect 82630 341728 82694 341732
rect 82630 341672 82634 341728
rect 82634 341672 82690 341728
rect 82690 341672 82694 341728
rect 82630 341668 82694 341672
rect 82492 339628 82556 339692
rect 82308 339008 82372 339012
rect 82308 338952 82358 339008
rect 82358 338952 82372 339008
rect 82308 338948 82372 338952
rect 501460 338948 501524 339012
rect 502012 338948 502076 339012
rect 504036 338948 504100 339012
rect 504588 338948 504652 339012
rect 502012 338812 502076 338876
rect 504588 338872 504652 338876
rect 504588 338816 504602 338872
rect 504602 338816 504652 338872
rect 504588 338812 504652 338816
rect 80836 337996 80900 338060
rect 82492 336772 82556 336836
rect 82492 335064 82556 335068
rect 82492 335008 82542 335064
rect 82542 335008 82556 335064
rect 82492 335004 82556 335008
rect 82492 332148 82556 332212
rect 82308 331256 82372 331260
rect 82308 331200 82358 331256
rect 82358 331200 82372 331256
rect 82308 331196 82372 331200
rect 82492 331196 82556 331260
rect 82492 331120 82556 331124
rect 82492 331064 82542 331120
rect 82542 331064 82556 331120
rect 82492 331060 82556 331064
rect 506796 328400 506860 328404
rect 506796 328344 506846 328400
rect 506846 328344 506860 328400
rect 506796 328340 506860 328344
rect 80836 328068 80900 328132
rect 78260 327796 78324 327860
rect 80836 327796 80900 327860
rect 504588 326436 504652 326500
rect 504036 326300 504100 326364
rect 504588 326300 504652 326364
rect 504036 326164 504100 326228
rect 501644 325620 501708 325684
rect 506796 323640 506860 323644
rect 506796 323584 506846 323640
rect 506846 323584 506860 323640
rect 506796 323580 506860 323584
rect 507532 319500 507596 319564
rect 507532 318820 507596 318884
rect 82492 317384 82556 317388
rect 82492 317328 82506 317384
rect 82506 317328 82556 317384
rect 82492 317324 82556 317328
rect 504588 316780 504652 316844
rect 504036 316644 504100 316708
rect 504588 316644 504652 316708
rect 504036 316508 504100 316572
rect 82492 316296 82556 316300
rect 82492 316240 82506 316296
rect 82506 316240 82556 316296
rect 82492 316236 82556 316240
rect 507348 315964 507412 316028
rect 501828 315828 501892 315892
rect 503300 313244 503364 313308
rect 82492 312352 82556 312356
rect 82492 312296 82506 312352
rect 82506 312296 82556 312352
rect 82492 312292 82556 312296
rect 501644 308484 501708 308548
rect 82492 307456 82556 307460
rect 82492 307400 82506 307456
rect 82506 307400 82556 307456
rect 82492 307396 82556 307400
rect 504588 307124 504652 307188
rect 504036 306988 504100 307052
rect 504588 306988 504652 307052
rect 501460 306852 501524 306916
rect 501644 306852 501708 306916
rect 81020 298828 81084 298892
rect 82492 297800 82556 297804
rect 82492 297744 82542 297800
rect 82542 297744 82556 297800
rect 82492 297740 82556 297744
rect 82492 297468 82556 297532
rect 504036 297468 504100 297532
rect 504588 297468 504652 297532
rect 504404 297332 504468 297396
rect 506980 297392 507044 297396
rect 506980 297336 507030 297392
rect 507030 297336 507044 297392
rect 506980 297332 507044 297336
rect 82492 296788 82556 296852
rect 78260 295428 78324 295492
rect 80836 293388 80900 293452
rect 82492 293388 82556 293452
rect 82492 292028 82556 292092
rect 82308 291076 82372 291140
rect 502012 290456 502076 290460
rect 502012 290400 502026 290456
rect 502026 290400 502076 290456
rect 502012 290396 502076 290400
rect 506980 290396 507044 290460
rect 507348 290396 507412 290460
rect 501460 290260 501524 290324
rect 504220 290124 504284 290188
rect 501460 289988 501524 290052
rect 82492 289096 82556 289100
rect 82492 289040 82542 289096
rect 82542 289040 82556 289096
rect 82492 289036 82556 289040
rect 501276 289036 501340 289100
rect 501644 289036 501708 289100
rect 504036 286996 504100 287060
rect 504220 286996 504284 287060
rect 501460 286316 501524 286380
rect 501828 286316 501892 286380
rect 501276 284684 501340 284748
rect 501460 282372 501524 282436
rect 502012 282296 502076 282300
rect 502012 282240 502026 282296
rect 502026 282240 502076 282296
rect 502012 282236 502076 282240
rect 501276 281420 501340 281484
rect 78260 280876 78324 280940
rect 82308 280876 82372 280940
rect 507348 280740 507412 280804
rect 501644 276524 501708 276588
rect 501460 276252 501524 276316
rect 501828 275844 501892 275908
rect 501460 275164 501524 275228
rect 501460 275028 501524 275092
rect 501460 274892 501524 274956
rect 502012 274892 502076 274956
rect 501276 274076 501340 274140
rect 502196 274076 502260 274140
rect 78260 273940 78324 274004
rect 78260 273396 78324 273460
rect 501644 273260 501708 273324
rect 501460 273124 501524 273188
rect 501460 272852 501524 272916
rect 501644 272580 501708 272644
rect 501460 272444 501524 272508
rect 501276 272308 501340 272372
rect 504588 271764 504652 271828
rect 501276 270812 501340 270876
rect 80836 270540 80900 270604
rect 502012 270540 502076 270604
rect 506980 270540 507044 270604
rect 501276 270404 501340 270468
rect 504588 270268 504652 270332
rect 78260 269588 78324 269652
rect 501276 268228 501340 268292
rect 502012 267140 502076 267204
rect 501276 267004 501340 267068
rect 504588 267004 504652 267068
rect 82630 266188 82694 266252
rect 501276 263468 501340 263532
rect 507532 263604 507596 263668
rect 502012 263332 502076 263396
rect 77892 262788 77956 262852
rect 82630 262788 82694 262852
rect 501644 262380 501708 262444
rect 506980 261428 507044 261492
rect 507348 261428 507412 261492
rect 78260 260748 78324 260812
rect 82630 260748 82694 260812
rect 82630 260204 82694 260268
rect 501276 260204 501340 260268
rect 501828 259796 501892 259860
rect 501276 258708 501340 258772
rect 501276 256668 501340 256732
rect 501460 256260 501524 256324
rect 501828 256260 501892 256324
rect 501460 256124 501524 256188
rect 77708 255444 77772 255508
rect 77892 255444 77956 255508
rect 502196 255580 502260 255644
rect 501644 255444 501708 255508
rect 502196 255444 502260 255508
rect 501644 255308 501708 255372
rect 501828 255036 501892 255100
rect 82492 254824 82556 254828
rect 82492 254768 82542 254824
rect 82542 254768 82556 254824
rect 82492 254764 82556 254768
rect 501828 254492 501892 254556
rect 501644 254084 501708 254148
rect 77892 253948 77956 254012
rect 82492 253948 82556 254012
rect 501276 253132 501340 253196
rect 501460 253132 501524 253196
rect 82492 252784 82556 252788
rect 82492 252728 82542 252784
rect 82542 252728 82556 252784
rect 82492 252724 82556 252728
rect 77708 252316 77772 252380
rect 78260 252316 78324 252380
rect 501644 251908 501708 251972
rect 504036 251908 504100 251972
rect 501644 251772 501708 251836
rect 502196 251772 502260 251836
rect 503484 249732 503548 249796
rect 504220 249732 504284 249796
rect 501276 249596 501340 249660
rect 504404 249596 504468 249660
rect 501460 249324 501524 249388
rect 501460 249052 501524 249116
rect 88748 248024 88812 248028
rect 88748 247968 88762 248024
rect 88762 247968 88812 248024
rect 88748 247964 88812 247968
rect 77524 247828 77588 247892
rect 88380 247752 88444 247756
rect 88380 247696 88430 247752
rect 88430 247696 88444 247752
rect 88380 247692 88444 247696
rect 501460 246604 501524 246668
rect 504220 246468 504284 246532
rect 501460 246060 501524 246124
rect 504036 246060 504100 246124
rect 502196 244836 502260 244900
rect 502196 244700 502260 244764
rect 501460 244564 501524 244628
rect 501828 244564 501892 244628
rect 501460 244428 501524 244492
rect 502012 244428 502076 244492
rect 501460 244292 501524 244356
rect 502012 244156 502076 244220
rect 501644 242660 501708 242724
rect 78260 242524 78324 242588
rect 501276 242524 501340 242588
rect 81020 241436 81084 241500
rect 501460 242388 501524 242452
rect 501460 242116 501524 242180
rect 501828 242252 501892 242316
rect 503484 242116 503548 242180
rect 504036 242116 504100 242180
rect 507348 242116 507412 242180
rect 501644 241980 501708 242044
rect 503484 241980 503548 242044
rect 501460 241708 501524 241772
rect 507532 241708 507596 241772
rect 501460 241436 501524 241500
rect 501644 241436 501708 241500
rect 80836 241300 80900 241364
rect 81204 241300 81268 241364
rect 81388 241300 81452 241364
rect 80836 240756 80900 240820
rect 81204 240756 81268 240820
rect 81388 240756 81452 240820
rect 81020 239396 81084 239460
rect 82538 239456 82602 239460
rect 82538 239400 82542 239456
rect 82542 239400 82598 239456
rect 82598 239400 82602 239456
rect 82538 239396 82602 239400
rect 82492 238368 82556 238372
rect 82492 238312 82506 238368
rect 82506 238312 82556 238368
rect 82492 238308 82556 238312
rect 504404 238988 504468 239052
rect 501276 238036 501340 238100
rect 501828 238036 501892 238100
rect 501460 237764 501524 237828
rect 501644 237764 501708 237828
rect 78076 237628 78140 237692
rect 501828 237628 501892 237692
rect 501460 237492 501524 237556
rect 501644 237492 501708 237556
rect 501276 237220 501340 237284
rect 501828 237220 501892 237284
rect 80284 237008 80348 237012
rect 80284 236952 80334 237008
rect 80334 236952 80348 237008
rect 80284 236948 80348 236952
rect 82492 236948 82556 237012
rect 82492 236132 82556 236196
rect 501276 235724 501340 235788
rect 501276 235588 501340 235652
rect 503484 235588 503548 235652
rect 82492 235104 82556 235108
rect 82492 235048 82506 235104
rect 82506 235048 82556 235104
rect 82492 235044 82556 235048
rect 504588 235452 504652 235516
rect 504036 235316 504100 235380
rect 504588 235316 504652 235380
rect 506980 235376 507044 235380
rect 506980 235320 507030 235376
rect 507030 235320 507044 235376
rect 506980 235316 507044 235320
rect 82492 234772 82556 234836
rect 82492 233684 82556 233748
rect 82492 233412 82556 233476
rect 502012 233140 502076 233204
rect 88748 233064 88812 233068
rect 88748 233008 88762 233064
rect 88762 233008 88812 233064
rect 88748 233004 88812 233008
rect 87828 232792 87892 232796
rect 87828 232736 87878 232792
rect 87878 232736 87892 232792
rect 87828 232732 87892 232736
rect 82308 232596 82372 232660
rect 82492 232596 82556 232660
rect 502380 231780 502444 231844
rect 502380 231236 502444 231300
rect 82492 230964 82556 231028
rect 78260 230828 78324 230892
rect 82492 230828 82556 230892
rect 82308 230556 82372 230620
rect 82492 229468 82556 229532
rect 82492 229196 82556 229260
rect 503484 229060 503548 229124
rect 82492 227836 82556 227900
rect 84516 226808 84580 226812
rect 84516 226752 84566 226808
rect 84566 226752 84580 226808
rect 84516 226748 84580 226752
rect 86172 226808 86236 226812
rect 86172 226752 86186 226808
rect 86186 226752 86236 226808
rect 86172 226748 86236 226752
rect 501828 226612 501892 226676
rect 502196 226612 502260 226676
rect 502196 226476 502260 226540
rect 82308 225660 82372 225724
rect 501276 225116 501340 225180
rect 501276 224844 501340 224908
rect 82492 223348 82556 223412
rect 501460 223620 501524 223684
rect 501460 222532 501524 222596
rect 501276 222124 501340 222188
rect 501276 221580 501340 221644
rect 504036 221988 504100 222052
rect 504404 221988 504468 222052
rect 504588 221852 504652 221916
rect 501276 221444 501340 221508
rect 501828 221444 501892 221508
rect 502012 221444 502076 221508
rect 82492 220084 82556 220148
rect 78260 219948 78324 220012
rect 82492 219948 82556 220012
rect 82492 219812 82556 219876
rect 501460 220220 501524 220284
rect 501828 219948 501892 220012
rect 502196 219948 502260 220012
rect 502196 219812 502260 219876
rect 501460 219676 501524 219740
rect 502012 216276 502076 216340
rect 501460 215868 501524 215932
rect 502196 215732 502260 215796
rect 504036 214508 504100 214572
rect 504404 214508 504468 214572
rect 502196 211788 502260 211852
rect 501276 211516 501340 211580
rect 504588 211516 504652 211580
rect 504036 210700 504100 210764
rect 82630 210428 82694 210492
rect 82308 209340 82372 209404
rect 502012 209204 502076 209268
rect 82492 209068 82556 209132
rect 82308 207980 82372 208044
rect 82630 207708 82694 207772
rect 77708 206212 77772 206276
rect 78260 206212 78324 206276
rect 77524 206076 77588 206140
rect 78260 206076 78324 206140
rect 501460 204852 501524 204916
rect 502150 204036 502214 204100
rect 501276 203628 501340 203692
rect 501460 203356 501524 203420
rect 504588 203356 504652 203420
rect 501460 203220 501524 203284
rect 502012 203220 502076 203284
rect 77892 203084 77956 203148
rect 82492 203084 82556 203148
rect 82492 202948 82556 203012
rect 78076 202676 78140 202740
rect 82492 201996 82556 202060
rect 77156 201860 77220 201924
rect 82492 201860 82556 201924
rect 82492 201724 82556 201788
rect 501276 203084 501340 203148
rect 501644 202132 501708 202196
rect 502196 202132 502260 202196
rect 82630 201588 82694 201652
rect 82308 201452 82372 201516
rect 82308 201180 82372 201244
rect 82492 201044 82556 201108
rect 76052 200908 76116 200972
rect 77524 200908 77588 200972
rect 82308 200772 82372 200836
rect 501460 201180 501524 201244
rect 501276 200364 501340 200428
rect 502012 200364 502076 200428
rect 78260 200228 78324 200292
rect 82492 199548 82556 199612
rect 501644 199412 501708 199476
rect 504036 199412 504100 199476
rect 504036 199276 504100 199340
rect 77156 198052 77220 198116
rect 501828 198052 501892 198116
rect 502012 197372 502076 197436
rect 502012 196828 502076 196892
rect 501460 196692 501524 196756
rect 502012 196692 502076 196756
rect 501460 196284 501524 196348
rect 504588 196284 504652 196348
rect 501276 196148 501340 196212
rect 501460 195740 501524 195804
rect 501460 195468 501524 195532
rect 82630 195332 82694 195396
rect 82492 195196 82556 195260
rect 82630 194984 82694 194988
rect 82630 194928 82634 194984
rect 82634 194928 82690 194984
rect 82690 194928 82694 194984
rect 82630 194924 82694 194928
rect 82630 194848 82694 194852
rect 82630 194792 82634 194848
rect 82634 194792 82690 194848
rect 82690 194792 82694 194848
rect 82630 194788 82694 194792
rect 77708 194652 77772 194716
rect 501460 194380 501524 194444
rect 506980 193836 507044 193900
rect 507348 193836 507412 193900
rect 501460 193156 501524 193220
rect 504588 193156 504652 193220
rect 503484 193020 503548 193084
rect 503484 192884 503548 192948
rect 504036 192884 504100 192948
rect 82492 192340 82556 192404
rect 82630 192340 82694 192404
rect 82492 191932 82556 191996
rect 82630 191388 82694 191452
rect 501276 191388 501340 191452
rect 504588 191388 504652 191452
rect 501276 191252 501340 191316
rect 501644 191252 501708 191316
rect 82492 191116 82556 191180
rect 82492 190844 82556 190908
rect 501460 191116 501524 191180
rect 501644 191116 501708 191180
rect 502196 191116 502260 191180
rect 501460 190980 501524 191044
rect 502012 190980 502076 191044
rect 502012 190844 502076 190908
rect 503484 190844 503548 190908
rect 502196 190708 502260 190772
rect 82308 190436 82372 190500
rect 82630 190300 82694 190364
rect 501276 189756 501340 189820
rect 82492 188668 82556 188732
rect 78260 188396 78324 188460
rect 82492 187308 82556 187372
rect 82630 187096 82694 187100
rect 82630 187040 82634 187096
rect 82634 187040 82690 187096
rect 82690 187040 82694 187096
rect 82630 187036 82694 187040
rect 82492 186900 82556 186964
rect 502012 186900 502076 186964
rect 503484 186900 503548 186964
rect 504220 186764 504284 186828
rect 502196 186356 502260 186420
rect 501276 186220 501340 186284
rect 77524 184588 77588 184652
rect 504404 185812 504468 185876
rect 501460 184724 501524 184788
rect 501644 184724 501708 184788
rect 501828 184724 501892 184788
rect 502012 184724 502076 184788
rect 501828 184452 501892 184516
rect 502012 184452 502076 184516
rect 501276 184316 501340 184380
rect 501460 184316 501524 184380
rect 501644 184316 501708 184380
rect 502196 183772 502260 183836
rect 504220 183772 504284 183836
rect 502196 183636 502260 183700
rect 503484 183636 503548 183700
rect 502012 183500 502076 183564
rect 501460 182276 501524 182340
rect 502012 182276 502076 182340
rect 502196 182004 502260 182068
rect 501460 181868 501524 181932
rect 502196 181868 502260 181932
rect 501460 181732 501524 181796
rect 82492 181324 82556 181388
rect 82308 181052 82372 181116
rect 507532 181052 507596 181116
rect 502196 180100 502260 180164
rect 77892 179964 77956 180028
rect 501460 179964 501524 180028
rect 503484 180100 503548 180164
rect 82492 179828 82556 179892
rect 87322 179888 87386 179892
rect 87322 179832 87326 179888
rect 87326 179832 87382 179888
rect 87382 179832 87386 179888
rect 87322 179828 87386 179832
rect 88748 179888 88812 179892
rect 88748 179832 88762 179888
rect 88762 179832 88812 179888
rect 88748 179828 88812 179832
rect 501276 179148 501340 179212
rect 502196 178876 502260 178940
rect 82492 178604 82556 178668
rect 501276 178468 501340 178532
rect 504588 178468 504652 178532
rect 82492 178332 82556 178396
rect 501460 178332 501524 178396
rect 501460 178196 501524 178260
rect 501460 178060 501524 178124
rect 502012 177244 502076 177308
rect 501460 177108 501524 177172
rect 502012 177108 502076 177172
rect 501460 176972 501524 177036
rect 501276 175748 501340 175812
rect 504220 175748 504284 175812
rect 501276 175612 501340 175676
rect 502012 175612 502076 175676
rect 502012 175476 502076 175540
rect 502196 175476 502260 175540
rect 502196 175340 502260 175404
rect 82308 174524 82372 174588
rect 82630 175068 82694 175132
rect 82492 173844 82556 173908
rect 82630 173708 82694 173772
rect 502196 173980 502260 174044
rect 501644 173300 501708 173364
rect 501644 173164 501708 173228
rect 502196 173028 502260 173092
rect 504220 173164 504284 173228
rect 506980 173164 507044 173228
rect 507348 173164 507412 173228
rect 77892 172348 77956 172412
rect 82630 172348 82694 172412
rect 501276 172348 501340 172412
rect 504588 172348 504652 172412
rect 82492 171804 82556 171868
rect 82492 171532 82556 171596
rect 87322 171592 87386 171596
rect 87322 171536 87326 171592
rect 87326 171536 87382 171592
rect 87382 171536 87386 171592
rect 87322 171532 87386 171536
rect 87644 171592 87708 171596
rect 87644 171536 87658 171592
rect 87658 171536 87708 171592
rect 87644 171532 87708 171536
rect 82630 171396 82694 171460
rect 501828 171124 501892 171188
rect 82630 170988 82694 171052
rect 82124 170580 82188 170644
rect 82492 170444 82556 170508
rect 82630 170444 82694 170508
rect 501644 170444 501708 170508
rect 502012 170444 502076 170508
rect 502196 170172 502260 170236
rect 82492 170036 82556 170100
rect 82124 169764 82188 169828
rect 501828 166364 501892 166428
rect 501828 165956 501892 166020
rect 502012 165956 502076 166020
rect 502012 165820 502076 165884
rect 78260 165548 78324 165612
rect 504588 165412 504652 165476
rect 503484 165004 503548 165068
rect 503484 164868 503548 164932
rect 504220 164868 504284 164932
rect 506980 164868 507044 164932
rect 507348 164868 507412 164932
rect 501460 163780 501524 163844
rect 501460 163644 501524 163708
rect 501460 162828 501524 162892
rect 501460 162420 501524 162484
rect 501644 162284 501708 162348
rect 82492 162148 82556 162212
rect 501276 161740 501340 161804
rect 501276 161332 501340 161396
rect 504036 161332 504100 161396
rect 82492 160788 82556 160852
rect 501644 160788 501708 160852
rect 502012 160788 502076 160852
rect 77892 159020 77956 159084
rect 82308 159020 82372 159084
rect 501828 158884 501892 158948
rect 502012 158748 502076 158812
rect 504588 158068 504652 158132
rect 501276 157932 501340 157996
rect 504036 157932 504100 157996
rect 501644 157448 501708 157452
rect 501644 157392 501658 157448
rect 501658 157392 501708 157448
rect 501644 157388 501708 157392
rect 504588 157388 504652 157452
rect 82492 157252 82556 157316
rect 82308 156708 82372 156772
rect 82630 156708 82694 156772
rect 501460 156572 501524 156636
rect 503484 155756 503548 155820
rect 504220 155756 504284 155820
rect 502196 155620 502260 155684
rect 503484 155620 503548 155684
rect 502196 155212 502260 155276
rect 506980 155212 507044 155276
rect 507348 155212 507412 155276
rect 501460 152084 501524 152148
rect 501460 150860 501524 150924
rect 82492 149636 82556 149700
rect 501460 148820 501524 148884
rect 501460 148548 501524 148612
rect 507348 148548 507412 148612
rect 501276 147460 501340 147524
rect 507532 147324 507596 147388
rect 501460 147188 501524 147252
rect 503484 146916 503548 146980
rect 82308 146780 82372 146844
rect 501460 145964 501524 146028
rect 501460 145828 501524 145892
rect 507348 145828 507412 145892
rect 506980 145556 507044 145620
rect 507348 145556 507412 145620
rect 82308 144468 82372 144532
rect 503484 143924 503548 143988
rect 82492 143108 82556 143172
rect 82492 141884 82556 141948
rect 501276 140524 501340 140588
rect 501276 140388 501340 140452
rect 501276 140252 501340 140316
rect 501460 140116 501524 140180
rect 501828 140040 501892 140044
rect 501828 139984 501878 140040
rect 501878 139984 501892 140040
rect 501828 139980 501892 139984
rect 501828 139844 501892 139908
rect 506244 139300 506308 139364
rect 506980 139300 507044 139364
rect 503484 138756 503548 138820
rect 501460 138620 501524 138684
rect 501828 138620 501892 138684
rect 503484 138620 503548 138684
rect 504036 138620 504100 138684
rect 501460 138484 501524 138548
rect 501460 138348 501524 138412
rect 502012 137940 502076 138004
rect 501644 137804 501708 137868
rect 502012 137668 502076 137732
rect 80836 137396 80900 137460
rect 80836 137260 80900 137324
rect 82492 137396 82556 137460
rect 82308 137260 82372 137324
rect 501276 136988 501340 137052
rect 501276 136716 501340 136780
rect 501828 136580 501892 136644
rect 504036 137260 504100 137324
rect 501460 136308 501524 136372
rect 82308 136036 82372 136100
rect 82492 136036 82556 136100
rect 82308 135900 82372 135964
rect 501460 135084 501524 135148
rect 504036 135084 504100 135148
rect 504036 134948 504100 135012
rect 501460 134812 501524 134876
rect 501644 134812 501708 134876
rect 501276 133452 501340 133516
rect 507348 133860 507412 133924
rect 506244 131956 506308 132020
rect 501276 130868 501340 130932
rect 77524 130460 77588 130524
rect 504036 130596 504100 130660
rect 504036 130460 504100 130524
rect 82492 128964 82556 129028
rect 501276 126108 501340 126172
rect 504036 125972 504100 126036
rect 503484 125156 503548 125220
rect 504036 125156 504100 125220
rect 502196 125020 502260 125084
rect 502196 124884 502260 124948
rect 503484 124884 503548 124948
rect 77892 123932 77956 123996
rect 83780 123932 83844 123996
rect 84332 123932 84396 123996
rect 86724 123932 86788 123996
rect 88380 123932 88444 123996
rect 90772 123932 90836 123996
rect 90956 123932 91020 123996
rect 107700 123932 107764 123996
rect 463556 123932 463620 123996
rect 491892 123932 491956 123996
rect 493548 123932 493612 123996
rect 497964 123932 498028 123996
rect 498332 123932 498396 123996
rect 499068 123932 499132 123996
rect 499620 123932 499684 123996
rect 500724 123932 500788 123996
rect 122788 123796 122852 123860
rect 425468 123796 425532 123860
rect 493180 123796 493244 123860
rect 497228 123796 497292 123860
rect 499436 123796 499500 123860
rect 90956 123660 91020 123724
rect 91140 123660 91204 123724
rect 207060 123660 207124 123724
rect 320036 123660 320100 123724
rect 82676 123524 82740 123588
rect 87460 123524 87524 123588
rect 218100 123524 218164 123588
rect 234108 123524 234172 123588
rect 235212 123524 235276 123588
rect 240180 123524 240244 123588
rect 253060 123524 253124 123588
rect 275876 123524 275940 123588
rect 498516 123524 498580 123588
rect 499436 123660 499500 123724
rect 501276 123796 501340 123860
rect 500908 123660 500972 123724
rect 499804 123524 499868 123588
rect 86172 123388 86236 123452
rect 92612 123388 92676 123452
rect 252508 123388 252572 123452
rect 258028 123388 258092 123452
rect 260052 123388 260116 123452
rect 88564 123252 88628 123316
rect 93716 123252 93780 123316
rect 209820 123252 209884 123316
rect 219204 123252 219268 123316
rect 84700 123116 84764 123180
rect 271644 123116 271708 123180
rect 277348 123388 277412 123452
rect 295196 123388 295260 123452
rect 296668 123388 296732 123452
rect 314516 123388 314580 123452
rect 315988 123388 316052 123452
rect 333836 123388 333900 123452
rect 335308 123388 335372 123452
rect 353156 123388 353220 123452
rect 354628 123388 354692 123452
rect 372476 123388 372540 123452
rect 373948 123388 374012 123452
rect 391796 123388 391860 123452
rect 393268 123388 393332 123452
rect 411116 123388 411180 123452
rect 412588 123388 412652 123452
rect 277532 123252 277596 123316
rect 285628 123252 285692 123316
rect 296852 123252 296916 123316
rect 304948 123252 305012 123316
rect 316172 123252 316236 123316
rect 324268 123252 324332 123316
rect 335492 123252 335556 123316
rect 343588 123252 343652 123316
rect 354812 123252 354876 123316
rect 362908 123252 362972 123316
rect 374132 123252 374196 123316
rect 382228 123252 382292 123316
rect 393452 123252 393516 123316
rect 401548 123252 401612 123316
rect 412772 123252 412836 123316
rect 469260 123388 469324 123452
rect 478644 123388 478708 123452
rect 493364 123388 493428 123452
rect 466316 123252 466380 123316
rect 474044 123252 474108 123316
rect 478276 123252 478340 123316
rect 500540 123388 500604 123452
rect 500724 123252 500788 123316
rect 493180 123116 493244 123180
rect 499436 123116 499500 123180
rect 499804 123116 499868 123180
rect 77524 122980 77588 123044
rect 86908 122980 86972 123044
rect 88932 122980 88996 123044
rect 92612 122980 92676 123044
rect 285628 122980 285692 123044
rect 295196 122980 295260 123044
rect 304948 122980 305012 123044
rect 314516 122980 314580 123044
rect 324268 122980 324332 123044
rect 333836 122980 333900 123044
rect 343588 122980 343652 123044
rect 353156 122980 353220 123044
rect 362908 122980 362972 123044
rect 372476 122980 372540 123044
rect 382228 122980 382292 123044
rect 391796 122980 391860 123044
rect 401548 122980 401612 123044
rect 411116 122980 411180 123044
rect 493364 122980 493428 123044
rect 500724 122980 500788 123044
rect 99236 122844 99300 122908
rect 369900 122844 369964 122908
rect 379284 122844 379348 122908
rect 417556 122844 417620 122908
rect 420132 122844 420196 122908
rect 425100 122844 425164 122908
rect 434484 122844 434548 122908
rect 469444 122844 469508 122908
rect 478644 122844 478708 122908
rect 486556 122844 486620 122908
rect 88932 122708 88996 122772
rect 87828 122572 87892 122636
rect 78628 122300 78692 122364
rect 89300 122708 89364 122772
rect 91324 122708 91388 122772
rect 237236 122708 237300 122772
rect 89484 122572 89548 122636
rect 90588 122632 90652 122636
rect 90588 122576 90638 122632
rect 90638 122576 90652 122632
rect 90588 122572 90652 122576
rect 91876 122572 91940 122636
rect 114324 122572 114388 122636
rect 114692 122572 114756 122636
rect 172468 122572 172532 122636
rect 191972 122572 192036 122636
rect 500356 122632 500420 122636
rect 500356 122576 500370 122632
rect 500370 122576 500420 122632
rect 500356 122572 500420 122576
rect 507716 122572 507780 122636
rect 90036 122436 90100 122500
rect 506612 122436 506676 122500
rect 89300 122300 89364 122364
rect 92796 122300 92860 122364
rect 191788 122300 191852 122364
rect 508084 122300 508148 122364
rect 83780 122224 83844 122228
rect 83780 122168 83830 122224
rect 83830 122168 83844 122224
rect 83780 122164 83844 122168
rect 84884 122164 84948 122228
rect 114692 122164 114756 122228
rect 230428 122164 230492 122228
rect 269068 122164 269132 122228
rect 288388 122164 288452 122228
rect 299428 122164 299492 122228
rect 299612 122164 299676 122228
rect 327028 122164 327092 122228
rect 346348 122164 346412 122228
rect 365668 122164 365732 122228
rect 434668 122164 434732 122228
rect 444236 122164 444300 122228
rect 478276 122164 478340 122228
rect 478644 122164 478708 122228
rect 491892 122164 491956 122228
rect 495388 122164 495452 122228
rect 497412 122164 497476 122228
rect 84516 122028 84580 122092
rect 87276 122028 87340 122092
rect 91508 122028 91572 122092
rect 90588 121892 90652 121956
rect 172468 121756 172532 121820
rect 318748 122028 318812 122092
rect 319116 122028 319180 122092
rect 338068 122028 338132 122092
rect 338436 122028 338500 122092
rect 504588 122028 504652 122092
rect 215156 121892 215220 121956
rect 215524 121892 215588 121956
rect 237236 121892 237300 121956
rect 243492 121756 243556 121820
rect 259316 121756 259380 121820
rect 269068 121756 269132 121820
rect 281212 121756 281276 121820
rect 293172 121756 293236 121820
rect 318748 121892 318812 121956
rect 319116 121892 319180 121956
rect 338068 121892 338132 121956
rect 338620 121892 338684 121956
rect 506796 121892 506860 121956
rect 301452 121756 301516 121820
rect 322612 121756 322676 121820
rect 93716 121620 93780 121684
rect 230612 121620 230676 121684
rect 288388 121620 288452 121684
rect 327028 121620 327092 121684
rect 331076 121620 331140 121684
rect 344876 121620 344940 121684
rect 347084 121620 347148 121684
rect 365668 121620 365732 121684
rect 502932 121620 502996 121684
rect 89668 121484 89732 121548
rect 85068 121348 85132 121412
rect 116716 121348 116780 121412
rect 499436 121408 499500 121412
rect 499436 121352 499450 121408
rect 499450 121352 499500 121408
rect 499436 121348 499500 121352
rect 90220 121212 90284 121276
rect 505692 121212 505756 121276
rect 114324 121076 114388 121140
rect 495388 121076 495452 121140
rect 496492 121076 496556 121140
rect 501460 121076 501524 121140
rect 495940 120940 496004 121004
rect 498332 121000 498396 121004
rect 498332 120944 498382 121000
rect 498382 120944 498396 121000
rect 498332 120940 498396 120944
rect 498516 121000 498580 121004
rect 498516 120944 498566 121000
rect 498566 120944 498580 121000
rect 498516 120940 498580 120944
rect 501092 120940 501156 121004
rect 501644 120804 501708 120868
rect 82860 120668 82924 120732
rect 88196 120668 88260 120732
rect 501092 120668 501156 120732
rect 498516 120532 498580 120596
rect 507164 120396 507228 120460
rect 498700 120260 498764 120324
rect 499620 120260 499684 120324
rect 499988 120320 500052 120324
rect 499988 120264 500038 120320
rect 500038 120264 500052 120320
rect 499988 120260 500052 120264
rect 193260 120124 193324 120188
rect 196572 120124 196636 120188
rect 408540 120124 408604 120188
rect 422892 120124 422956 120188
rect 446628 120124 446692 120188
rect 453620 120124 453684 120188
rect 331260 119988 331324 120052
rect 340644 119988 340708 120052
rect 376708 119988 376772 120052
rect 85252 119852 85316 119916
rect 93348 119716 93412 119780
rect 92244 119580 92308 119644
rect 509740 119580 509804 119644
rect 87828 119172 87892 119236
rect 509372 119172 509436 119236
rect 89852 119036 89916 119100
rect 85620 118900 85684 118964
rect 394740 118900 394804 118964
rect 399524 118900 399588 118964
rect 453988 118900 454052 118964
rect 457300 118900 457364 118964
rect 497412 118900 497476 118964
rect 92612 118764 92676 118828
rect 174492 118628 174556 118692
rect 183324 118628 183388 118692
rect 186268 118628 186332 118692
rect 190500 118628 190564 118692
rect 251220 118628 251284 118692
rect 265572 118628 265636 118692
rect 269804 118628 269868 118692
rect 273668 118628 273732 118692
rect 315988 118628 316052 118692
rect 326844 118628 326908 118692
rect 394556 118628 394620 118692
rect 425100 118628 425164 118692
rect 434300 118628 434364 118692
rect 495940 118220 496004 118284
rect 504036 118220 504100 118284
rect 83228 118008 83292 118012
rect 83228 117952 83242 118008
rect 83242 117952 83292 118008
rect 83228 117948 83292 117952
rect 499804 117948 499868 118012
rect 493548 117192 493612 117196
rect 493548 117136 493562 117192
rect 493562 117136 493612 117192
rect 493548 117132 493612 117136
rect 85988 116920 86052 116924
rect 85988 116864 86038 116920
rect 86038 116864 86052 116920
rect 85988 116860 86052 116864
rect 86908 116724 86972 116788
rect 498332 116724 498396 116788
rect 505692 116724 505756 116788
rect 506244 116724 506308 116788
rect 78996 116588 79060 116652
rect 82308 116452 82372 116516
rect 500724 116180 500788 116244
rect 503484 116180 503548 116244
rect 499068 116044 499132 116108
rect 88012 115364 88076 115428
rect 88380 115364 88444 115428
rect 501276 115364 501340 115428
rect 504404 115228 504468 115292
rect 78812 115092 78876 115156
rect 500356 114608 500420 114612
rect 500356 114552 500406 114608
rect 500406 114552 500420 114608
rect 500356 114548 500420 114552
rect 500172 113188 500236 113252
rect 338068 111420 338132 111484
rect 473308 111420 473372 111484
rect 501092 111284 501156 111348
rect 87276 111148 87340 111212
rect 338068 111148 338132 111212
rect 473308 111148 473372 111212
rect 81204 111012 81268 111076
rect 396028 110876 396092 110940
rect 453988 110876 454052 110940
rect 396028 110604 396092 110668
rect 453988 110604 454052 110668
rect 500172 109712 500236 109716
rect 500172 109656 500186 109712
rect 500186 109656 500236 109712
rect 500172 109652 500236 109656
rect 82860 106932 82924 106996
rect 83412 106932 83476 106996
rect 84332 106992 84396 106996
rect 84332 106936 84346 106992
rect 84346 106936 84396 106992
rect 84332 106932 84396 106936
rect 86724 106932 86788 106996
rect 498516 106932 498580 106996
rect 499436 106932 499500 106996
rect 85988 106448 86052 106452
rect 85988 106392 86038 106448
rect 86038 106392 86052 106448
rect 85988 106388 86052 106392
rect 83228 106312 83292 106316
rect 83228 106256 83242 106312
rect 83242 106256 83292 106312
rect 83228 106252 83292 106256
rect 504404 105980 504468 106044
rect 85988 105844 86052 105908
rect 87092 105904 87156 105908
rect 87092 105848 87142 105904
rect 87142 105848 87156 105904
rect 87092 105844 87156 105848
rect 85988 105708 86052 105772
rect 83228 104816 83292 104820
rect 83228 104760 83278 104816
rect 83278 104760 83292 104816
rect 83228 104756 83292 104760
rect 500356 104756 500420 104820
rect 498884 104484 498948 104548
rect 499252 104484 499316 104548
rect 496860 102172 496924 102236
rect 497044 102172 497108 102236
rect 88196 101552 88260 101556
rect 88196 101496 88246 101552
rect 88246 101496 88260 101552
rect 88196 101492 88260 101496
rect 505692 101356 505756 101420
rect 84332 98696 84396 98700
rect 84332 98640 84346 98696
rect 84346 98640 84396 98696
rect 84332 98636 84396 98640
rect 504036 98636 504100 98700
rect 504404 98636 504468 98700
rect 82860 97956 82924 98020
rect 83412 97956 83476 98020
rect 289676 97064 289740 97068
rect 289676 97008 289726 97064
rect 289726 97008 289740 97064
rect 289676 97004 289740 97008
rect 500172 96792 500236 96796
rect 500172 96736 500186 96792
rect 500186 96736 500236 96792
rect 500172 96732 500236 96736
rect 504220 96732 504284 96796
rect 289676 96656 289740 96660
rect 289676 96600 289726 96656
rect 289726 96600 289740 96656
rect 289676 96596 289740 96600
rect 88196 96520 88260 96524
rect 88196 96464 88210 96520
rect 88210 96464 88260 96520
rect 88196 96460 88260 96464
rect 504220 96460 504284 96524
rect 88012 96384 88076 96388
rect 88012 96328 88026 96384
rect 88026 96328 88076 96384
rect 88012 96324 88076 96328
rect 83228 95296 83292 95300
rect 83228 95240 83278 95296
rect 83278 95240 83292 95296
rect 83228 95236 83292 95240
rect 499988 95160 500052 95164
rect 499988 95104 500002 95160
rect 500002 95104 500052 95160
rect 499988 95100 500052 95104
rect 88196 94616 88260 94620
rect 88196 94560 88210 94616
rect 88210 94560 88260 94616
rect 88196 94556 88260 94560
rect 500540 92848 500604 92852
rect 500540 92792 500590 92848
rect 500590 92792 500604 92848
rect 500540 92788 500604 92792
rect 88012 92712 88076 92716
rect 88012 92656 88026 92712
rect 88026 92656 88076 92712
rect 88012 92652 88076 92656
rect 500724 92712 500788 92716
rect 500724 92656 500738 92712
rect 500738 92656 500788 92712
rect 500724 92652 500788 92656
rect 88012 92380 88076 92444
rect 499436 92380 499500 92444
rect 499252 92244 499316 92308
rect 88012 91972 88076 92036
rect 500540 91760 500604 91764
rect 500540 91704 500590 91760
rect 500590 91704 500604 91760
rect 500540 91700 500604 91704
rect 87644 88300 87708 88364
rect 88196 88300 88260 88364
rect 504036 87680 504100 87684
rect 504036 87624 504050 87680
rect 504050 87624 504100 87680
rect 504036 87620 504100 87624
rect 501092 86940 501156 87004
rect 506060 86940 506124 87004
rect 83228 86864 83292 86868
rect 83228 86808 83278 86864
rect 83278 86808 83292 86864
rect 83228 86804 83292 86808
rect 84332 86320 84396 86324
rect 84332 86264 84382 86320
rect 84382 86264 84396 86320
rect 84332 86260 84396 86264
rect 87092 86320 87156 86324
rect 87092 86264 87142 86320
rect 87142 86264 87156 86320
rect 87092 86260 87156 86264
rect 82860 84900 82924 84964
rect 83412 84900 83476 84964
rect 502564 84764 502628 84828
rect 87460 84220 87524 84284
rect 87644 84220 87708 84284
rect 88012 84084 88076 84148
rect 88012 83812 88076 83876
rect 501092 82996 501156 83060
rect 500356 82860 500420 82924
rect 504220 80200 504284 80204
rect 504220 80144 504270 80200
rect 504270 80144 504284 80200
rect 504220 80140 504284 80144
rect 508268 80004 508332 80068
rect 82860 78644 82924 78708
rect 83412 78644 83476 78708
rect 84332 78024 84396 78028
rect 84332 77968 84382 78024
rect 84382 77968 84396 78024
rect 84332 77964 84396 77968
rect 87092 78024 87156 78028
rect 87092 77968 87142 78024
rect 87142 77968 87156 78024
rect 87092 77964 87156 77968
rect 87644 78024 87708 78028
rect 87644 77968 87658 78024
rect 87658 77968 87708 78024
rect 87644 77964 87708 77968
rect 88196 78024 88260 78028
rect 88196 77968 88246 78024
rect 88246 77968 88260 78024
rect 88196 77964 88260 77968
rect 83228 77344 83292 77348
rect 83228 77288 83278 77344
rect 83278 77288 83292 77344
rect 83228 77284 83292 77288
rect 504036 77344 504100 77348
rect 504036 77288 504050 77344
rect 504050 77288 504100 77344
rect 504036 77284 504100 77288
rect 504220 77344 504284 77348
rect 504220 77288 504270 77344
rect 504270 77288 504284 77344
rect 504220 77284 504284 77288
rect 500356 77208 500420 77212
rect 500356 77152 500406 77208
rect 500406 77152 500420 77208
rect 500356 77148 500420 77152
rect 83274 77072 83338 77076
rect 83274 77016 83278 77072
rect 83278 77016 83334 77072
rect 83334 77016 83338 77072
rect 83274 77012 83338 77016
rect 499252 72932 499316 72996
rect 152780 70348 152844 70412
rect 88196 69184 88260 69188
rect 88196 69128 88246 69184
rect 88246 69128 88260 69184
rect 88196 69124 88260 69128
rect 500356 68368 500420 68372
rect 500356 68312 500406 68368
rect 500406 68312 500420 68368
rect 500356 68308 500420 68312
rect 83228 67688 83292 67692
rect 83228 67632 83278 67688
rect 83278 67632 83292 67688
rect 83228 67628 83292 67632
rect 87644 67688 87708 67692
rect 87644 67632 87658 67688
rect 87658 67632 87708 67688
rect 87644 67628 87708 67632
rect 152780 67688 152844 67692
rect 152780 67632 152830 67688
rect 152830 67632 152844 67688
rect 152780 67628 152844 67632
rect 498516 67492 498580 67556
rect 85988 67220 86052 67284
rect 85988 67084 86052 67148
rect 82860 65452 82924 65516
rect 83412 65452 83476 65516
rect 85804 62792 85868 62796
rect 85804 62736 85818 62792
rect 85818 62736 85868 62792
rect 85804 62732 85868 62736
rect 498332 62792 498396 62796
rect 498332 62736 498382 62792
rect 498382 62736 498396 62792
rect 498332 62732 498396 62736
rect 87644 62188 87708 62252
rect 87460 61916 87524 61980
rect 152964 61432 153028 61436
rect 152964 61376 152978 61432
rect 152978 61376 153028 61432
rect 152964 61372 153028 61376
rect 501644 60692 501708 60756
rect 501828 60692 501892 60756
rect 83228 57896 83292 57900
rect 83228 57840 83278 57896
rect 83278 57840 83292 57896
rect 83228 57836 83292 57840
rect 87460 57896 87524 57900
rect 87460 57840 87510 57896
rect 87510 57840 87524 57896
rect 87460 57836 87524 57840
rect 498332 57836 498396 57900
rect 504036 57564 504100 57628
rect 504588 57564 504652 57628
rect 499988 56612 500052 56676
rect 500540 56536 500604 56540
rect 500540 56480 500554 56536
rect 500554 56480 500604 56536
rect 500540 56476 500604 56480
rect 82860 55796 82924 55860
rect 83412 55796 83476 55860
rect 499436 55252 499500 55316
rect 152964 50960 153028 50964
rect 152964 50904 153014 50960
rect 153014 50904 153028 50960
rect 152964 50900 153028 50904
rect 499988 49056 500052 49060
rect 499988 49000 500002 49056
rect 500002 49000 500052 49056
rect 499988 48996 500052 49000
rect 500356 49056 500420 49060
rect 500356 49000 500406 49056
rect 500406 49000 500420 49056
rect 500356 48996 500420 49000
rect 504220 48996 504284 49060
rect 504588 48996 504652 49060
rect 500540 48920 500604 48924
rect 500540 48864 500554 48920
rect 500554 48864 500604 48920
rect 500540 48860 500604 48864
rect 83228 48376 83292 48380
rect 83228 48320 83278 48376
rect 83278 48320 83292 48376
rect 83228 48316 83292 48320
rect 85804 48316 85868 48380
rect 87460 48376 87524 48380
rect 87460 48320 87510 48376
rect 87510 48320 87524 48376
rect 87460 48316 87524 48320
rect 498516 48316 498580 48380
rect 85988 48044 86052 48108
rect 85988 47772 86052 47836
rect 498516 44372 498580 44436
rect 498332 44236 498396 44300
rect 85804 43480 85868 43484
rect 85804 43424 85854 43480
rect 85854 43424 85868 43480
rect 85804 43420 85868 43424
rect 86724 40156 86788 40220
rect 87460 40156 87524 40220
rect 84332 39884 84396 39948
rect 84516 39884 84580 39948
rect 86540 39884 86604 39948
rect 87276 39884 87340 39948
rect 499988 38660 500052 38724
rect 504220 38660 504284 38724
rect 504404 38720 504468 38724
rect 504404 38664 504454 38720
rect 504454 38664 504468 38720
rect 504404 38660 504468 38664
rect 83228 38584 83292 38588
rect 83228 38528 83278 38584
rect 83278 38528 83292 38584
rect 83228 38524 83292 38528
rect 85804 37300 85868 37364
rect 499436 37300 499500 37364
rect 500540 37224 500604 37228
rect 500540 37168 500590 37224
rect 500590 37168 500604 37224
rect 500540 37164 500604 37168
rect 499620 37028 499684 37092
rect 87276 35260 87340 35324
rect 83412 35124 83476 35188
rect 498332 34368 498396 34372
rect 498332 34312 498346 34368
rect 498346 34312 498396 34368
rect 498332 34308 498396 34312
rect 499988 29684 500052 29748
rect 500356 29684 500420 29748
rect 500540 29744 500604 29748
rect 500540 29688 500590 29744
rect 500590 29688 500604 29744
rect 500540 29684 500604 29688
rect 83228 29004 83292 29068
rect 505876 29004 505940 29068
rect 85804 27568 85868 27572
rect 85804 27512 85854 27568
rect 85854 27512 85868 27568
rect 85804 27508 85868 27512
rect 497044 26284 497108 26348
rect 496860 26012 496924 26076
rect 498332 24924 498396 24988
rect 84332 23428 84396 23492
rect 84516 23428 84580 23492
rect 87460 23488 87524 23492
rect 87460 23432 87510 23488
rect 87510 23432 87524 23488
rect 87460 23428 87524 23432
rect 84332 23352 84396 23356
rect 84332 23296 84382 23352
rect 84382 23296 84396 23352
rect 84332 23292 84396 23296
rect 86540 22748 86604 22812
rect 507900 21932 507964 21996
rect 83228 19212 83292 19276
rect 85988 19272 86052 19276
rect 85988 19216 86002 19272
rect 86002 19216 86052 19272
rect 85988 19212 86052 19216
rect 498884 18940 498948 19004
rect 87460 18668 87524 18732
rect 499620 18668 499684 18732
rect 505508 18532 505572 18596
rect 85620 17988 85684 18052
rect 503668 17444 503732 17508
rect 503852 17308 503916 17372
rect 79180 17172 79244 17236
rect 503116 16356 503180 16420
rect 502380 16220 502444 16284
rect 504220 16084 504284 16148
rect 500540 15948 500604 16012
rect 498332 15268 498396 15332
rect 502748 14588 502812 14652
rect 81020 14452 81084 14516
rect 84332 13832 84396 13836
rect 84332 13776 84382 13832
rect 84382 13776 84396 13832
rect 84332 13772 84396 13776
rect 84332 13696 84396 13700
rect 84332 13640 84382 13696
rect 84382 13640 84396 13696
rect 84332 13636 84396 13640
rect 83044 12956 83108 13020
rect 82124 11732 82188 11796
rect 81756 11596 81820 11660
rect 79732 10508 79796 10572
rect 81572 10372 81636 10436
rect 504404 10236 504468 10300
rect 85620 9828 85684 9892
rect 85804 9692 85868 9756
rect 85988 9692 86052 9756
rect 498516 9752 498580 9756
rect 498516 9696 498530 9752
rect 498530 9696 498580 9752
rect 498516 9692 498580 9696
rect 85988 9420 86052 9484
rect 91692 8876 91756 8940
rect 500356 8876 500420 8940
rect 85804 8196 85868 8260
rect 93164 6836 93228 6900
rect 510660 6836 510724 6900
rect 85436 6700 85500 6764
rect 496860 6700 496924 6764
rect 79364 6564 79428 6628
rect 507532 6564 507596 6628
rect 81388 6428 81452 6492
rect 497412 6428 497476 6492
rect 79548 6292 79612 6356
rect 81940 6156 82004 6220
rect 88012 6020 88076 6084
rect 509188 6020 509252 6084
rect 92060 5884 92124 5948
rect 498516 5748 498580 5812
rect 498332 5612 498396 5676
rect 92980 5340 93044 5404
rect 89300 5204 89364 5268
rect 90404 5068 90468 5132
rect 502196 4932 502260 4996
rect 503300 4796 503364 4860
rect 86172 4720 86236 4724
rect 86172 4664 86186 4720
rect 86186 4664 86236 4720
rect 86172 4660 86236 4664
rect 164372 4388 164436 4452
rect 169156 4388 169220 4452
rect 172468 4388 172532 4452
rect 182036 4388 182100 4452
rect 329236 4388 329300 4452
rect 337884 4388 337948 4452
rect 396028 4388 396092 4452
rect 405596 4388 405660 4452
rect 415716 4388 415780 4452
rect 424916 4388 424980 4452
rect 434668 4388 434732 4452
rect 443316 4388 443380 4452
rect 444420 4252 444484 4316
rect 457484 4252 457548 4316
rect 84332 4176 84396 4180
rect 84332 4120 84382 4176
rect 84382 4120 84396 4176
rect 84332 4116 84396 4120
rect 86356 4176 86420 4180
rect 86356 4120 86406 4176
rect 86406 4120 86420 4176
rect 86356 4116 86420 4120
rect 84332 3844 84396 3908
rect 89116 3844 89180 3908
rect 86356 3708 86420 3772
rect 87092 3708 87156 3772
rect 92428 3844 92492 3908
rect 93532 3844 93596 3908
rect 275876 3980 275940 4044
rect 384988 4116 385052 4180
rect 479380 4116 479444 4180
rect 485636 4116 485700 4180
rect 500172 3980 500236 4044
rect 88196 3572 88260 3636
rect 116716 3708 116780 3772
rect 122788 3436 122852 3500
rect 164004 3708 164068 3772
rect 207060 3708 207124 3772
rect 218100 3708 218164 3772
rect 271644 3708 271708 3772
rect 318748 3844 318812 3908
rect 319116 3844 319180 3908
rect 495388 3844 495452 3908
rect 502012 3844 502076 3908
rect 318748 3708 318812 3772
rect 320036 3708 320100 3772
rect 342300 3708 342364 3772
rect 357388 3708 357452 3772
rect 365668 3708 365732 3772
rect 125548 3436 125612 3500
rect 125732 3436 125796 3500
rect 133828 3436 133892 3500
rect 143580 3436 143644 3500
rect 148180 3436 148244 3500
rect 153148 3436 153212 3500
rect 288388 3572 288452 3636
rect 307708 3572 307772 3636
rect 317276 3572 317340 3636
rect 327028 3572 327092 3636
rect 396028 3708 396092 3772
rect 460980 3708 461044 3772
rect 462452 3708 462516 3772
rect 463556 3708 463620 3772
rect 478644 3768 478708 3772
rect 478644 3712 478694 3768
rect 478694 3712 478708 3768
rect 478644 3708 478708 3712
rect 495204 3708 495268 3772
rect 507716 3708 507780 3772
rect 521700 3708 521764 3772
rect 531084 3708 531148 3772
rect 557948 3708 558012 3772
rect 384988 3572 385052 3636
rect 425468 3572 425532 3636
rect 495388 3572 495452 3636
rect 495572 3572 495636 3636
rect 172468 3436 172532 3500
rect 176516 3436 176580 3500
rect 499804 3436 499868 3500
rect 80836 3300 80900 3364
rect 498332 3300 498396 3364
rect 495756 3164 495820 3228
rect 84700 3028 84764 3092
rect 107700 3028 107764 3092
rect 243492 3028 243556 3092
rect 101260 2892 101324 2956
rect 114876 2892 114940 2956
rect 133828 2892 133892 2956
rect 143580 2892 143644 2956
rect 153148 2952 153212 2956
rect 153148 2896 153162 2952
rect 153162 2896 153212 2952
rect 153148 2892 153212 2896
rect 172468 2892 172532 2956
rect 252508 3028 252572 3092
rect 267596 3028 267660 3092
rect 288388 3028 288452 3092
rect 302004 3028 302068 3092
rect 306236 3028 306300 3092
rect 315988 3028 316052 3092
rect 325556 3028 325620 3092
rect 264468 2892 264532 2956
rect 268884 2892 268948 2956
rect 307708 2892 307772 2956
rect 317276 2892 317340 2956
rect 318748 2892 318812 2956
rect 357388 3028 357452 3092
rect 365668 3028 365732 3092
rect 378548 3028 378612 3092
rect 379652 3028 379716 3092
rect 396028 3028 396092 3092
rect 417556 3028 417620 3092
rect 419212 3028 419276 3092
rect 436140 3028 436204 3092
rect 437428 3028 437492 3092
rect 499068 3164 499132 3228
rect 496124 3028 496188 3092
rect 501644 3028 501708 3092
rect 513972 3028 514036 3092
rect 520044 3028 520108 3092
rect 327028 2892 327092 2956
rect 335308 2892 335372 2956
rect 340828 2892 340892 2956
rect 506428 2892 506492 2956
rect 451596 2620 451660 2684
rect 461348 2620 461412 2684
rect 486556 2756 486620 2820
rect 470548 2484 470612 2548
rect 479380 2484 479444 2548
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 3926 452437 3986 453102
rect 3923 452436 3989 452437
rect 3923 452372 3924 452436
rect 3988 452372 3989 452436
rect 3923 452371 3989 452372
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 79731 570076 79797 570077
rect 79731 570012 79732 570076
rect 79796 570012 79797 570076
rect 79731 570011 79797 570012
rect 79547 555932 79613 555933
rect 79547 555868 79548 555932
rect 79612 555868 79613 555932
rect 79547 555867 79613 555868
rect 79363 548860 79429 548861
rect 79363 548796 79364 548860
rect 79428 548796 79429 548860
rect 79363 548795 79429 548796
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 77155 510236 77221 510237
rect 77155 510172 77156 510236
rect 77220 510172 77221 510236
rect 77155 510171 77221 510172
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76054 200973 76114 216462
rect 76051 200972 76117 200973
rect 76051 200908 76052 200972
rect 76116 200908 76117 200972
rect 76051 200907 76117 200908
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 186054 77004 221498
rect 77158 201925 77218 510171
rect 79179 432716 79245 432717
rect 79179 432652 79180 432716
rect 79244 432652 79245 432716
rect 79179 432651 79245 432652
rect 78995 422108 79061 422109
rect 78995 422044 78996 422108
rect 79060 422044 79061 422108
rect 78995 422043 79061 422044
rect 78630 396218 78690 403462
rect 78811 383484 78877 383485
rect 78811 383420 78812 383484
rect 78876 383420 78877 383484
rect 78811 383419 78877 383420
rect 78262 375818 78322 382382
rect 78627 376412 78693 376413
rect 78627 376348 78628 376412
rect 78692 376348 78693 376412
rect 78627 376347 78693 376348
rect 78262 327861 78322 330702
rect 78259 327860 78325 327861
rect 78259 327796 78260 327860
rect 78324 327796 78325 327860
rect 78259 327795 78325 327796
rect 78262 298978 78322 302822
rect 77894 292858 77954 294662
rect 77526 273138 77586 283782
rect 78259 280940 78325 280941
rect 78259 280876 78260 280940
rect 78324 280876 78325 280940
rect 78259 280875 78325 280876
rect 78262 277898 78322 280875
rect 78262 274005 78322 274262
rect 78259 274004 78325 274005
rect 78259 273940 78260 274004
rect 78324 273940 78325 274004
rect 78259 273939 78325 273940
rect 78259 273460 78325 273461
rect 78259 273396 78260 273460
rect 78324 273396 78325 273460
rect 78259 273395 78325 273396
rect 78262 271098 78322 273395
rect 77894 264298 77954 266102
rect 77891 262852 77957 262853
rect 77891 262788 77892 262852
rect 77956 262788 77957 262852
rect 77891 262787 77957 262788
rect 77894 260218 77954 262787
rect 78259 260812 78325 260813
rect 78259 260748 78260 260812
rect 78324 260748 78325 260812
rect 78259 260747 78325 260748
rect 77894 255509 77954 258622
rect 77707 255508 77773 255509
rect 77707 255444 77708 255508
rect 77772 255444 77773 255508
rect 77707 255443 77773 255444
rect 77891 255508 77957 255509
rect 77891 255444 77892 255508
rect 77956 255444 77957 255508
rect 77891 255443 77957 255444
rect 77710 252381 77770 255443
rect 77891 254012 77957 254013
rect 77891 253948 77892 254012
rect 77956 253948 77957 254012
rect 77891 253947 77957 253948
rect 77707 252380 77773 252381
rect 77707 252316 77708 252380
rect 77772 252316 77773 252380
rect 77707 252315 77773 252316
rect 77894 242538 77954 253947
rect 78262 252738 78322 260747
rect 78259 252380 78325 252381
rect 78259 252316 78260 252380
rect 78324 252316 78325 252380
rect 78259 252315 78325 252316
rect 78262 245258 78322 252315
rect 78259 242588 78325 242589
rect 78259 242524 78260 242588
rect 78324 242524 78325 242588
rect 78259 242523 78325 242524
rect 78262 241178 78322 242523
rect 78262 230893 78322 233462
rect 78259 230892 78325 230893
rect 78259 230828 78260 230892
rect 78324 230828 78325 230892
rect 78259 230827 78325 230828
rect 77894 222818 77954 230742
rect 78259 220012 78325 220013
rect 78259 219948 78260 220012
rect 78324 219948 78325 220012
rect 78259 219947 78325 219948
rect 77894 216018 77954 219862
rect 77526 206141 77586 208302
rect 77707 206276 77773 206277
rect 77707 206212 77708 206276
rect 77772 206212 77773 206276
rect 77707 206211 77773 206212
rect 77523 206140 77589 206141
rect 77523 206076 77524 206140
rect 77588 206076 77589 206140
rect 77523 206075 77589 206076
rect 77155 201924 77221 201925
rect 77155 201860 77156 201924
rect 77220 201860 77221 201924
rect 77155 201859 77221 201860
rect 77523 200972 77589 200973
rect 77523 200908 77524 200972
rect 77588 200908 77589 200972
rect 77523 200907 77589 200908
rect 77155 198116 77221 198117
rect 77155 198052 77156 198116
rect 77220 198052 77221 198116
rect 77155 198051 77221 198052
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 77158 3858 77218 198051
rect 77526 194258 77586 200907
rect 77710 194717 77770 206211
rect 77894 203149 77954 212382
rect 78262 206277 78322 219947
rect 78259 206276 78325 206277
rect 78259 206212 78260 206276
rect 78324 206212 78325 206276
rect 78259 206211 78325 206212
rect 78259 206140 78325 206141
rect 78259 206076 78260 206140
rect 78324 206076 78325 206140
rect 78259 206075 78325 206076
rect 78262 205818 78322 206075
rect 77891 203148 77957 203149
rect 77891 203084 77892 203148
rect 77956 203084 77957 203148
rect 77891 203083 77957 203084
rect 78075 202740 78141 202741
rect 78075 202676 78076 202740
rect 78140 202676 78141 202740
rect 78075 202675 78141 202676
rect 78078 195618 78138 202675
rect 78262 200293 78322 202862
rect 78259 200292 78325 200293
rect 78259 200228 78260 200292
rect 78324 200228 78325 200292
rect 78259 200227 78325 200228
rect 77707 194716 77773 194717
rect 77707 194652 77708 194716
rect 77772 194652 77773 194716
rect 77707 194651 77773 194652
rect 77894 184058 77954 191302
rect 78259 188460 78325 188461
rect 78259 188396 78260 188460
rect 78324 188396 78325 188460
rect 78259 188395 78325 188396
rect 77891 180028 77957 180029
rect 77891 179964 77892 180028
rect 77956 179964 77957 180028
rect 77891 179963 77957 179964
rect 77894 177258 77954 179963
rect 78262 176578 78322 188395
rect 77891 172412 77957 172413
rect 77891 172348 77892 172412
rect 77956 172348 77957 172412
rect 77891 172347 77957 172348
rect 77894 162978 77954 172347
rect 78262 167058 78322 168862
rect 77891 159084 77957 159085
rect 77891 159020 77892 159084
rect 77956 159020 77957 159084
rect 77891 159019 77957 159020
rect 77894 155498 77954 159019
rect 78262 152098 78322 158662
rect 77526 130525 77586 130782
rect 77523 130524 77589 130525
rect 77523 130460 77524 130524
rect 77588 130460 77589 130524
rect 77523 130459 77589 130460
rect 77526 123045 77586 130102
rect 77894 123997 77954 150502
rect 78262 129658 78322 141662
rect 77891 123996 77957 123997
rect 77891 123932 77892 123996
rect 77956 123932 77957 123996
rect 77891 123931 77957 123932
rect 77523 123044 77589 123045
rect 77523 122980 77524 123044
rect 77588 122980 77589 123044
rect 77523 122979 77589 122980
rect 78630 122365 78690 376347
rect 78627 122364 78693 122365
rect 78627 122300 78628 122364
rect 78692 122300 78693 122364
rect 78627 122299 78693 122300
rect 78814 115157 78874 383419
rect 78998 116653 79058 422043
rect 78995 116652 79061 116653
rect 78995 116588 78996 116652
rect 79060 116588 79061 116652
rect 78995 116587 79061 116588
rect 78811 115156 78877 115157
rect 78811 115092 78812 115156
rect 78876 115092 78877 115156
rect 78811 115091 78877 115092
rect 79182 17237 79242 432651
rect 79179 17236 79245 17237
rect 79179 17172 79180 17236
rect 79244 17172 79245 17236
rect 79179 17171 79245 17172
rect 79366 6629 79426 548795
rect 79363 6628 79429 6629
rect 79363 6564 79364 6628
rect 79428 6564 79429 6628
rect 79363 6563 79429 6564
rect 79550 6357 79610 555867
rect 79734 10573 79794 570011
rect 80004 549654 80604 585098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 89483 700636 89549 700637
rect 89483 700572 89484 700636
rect 89548 700572 89549 700636
rect 89483 700571 89549 700572
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 89486 695469 89546 700571
rect 90219 699820 90285 699821
rect 90219 699756 90220 699820
rect 90284 699756 90285 699820
rect 90219 699755 90285 699756
rect 89483 695468 89549 695469
rect 89483 695404 89484 695468
rect 89548 695404 89549 695468
rect 89483 695403 89549 695404
rect 89851 689348 89917 689349
rect 89851 689284 89852 689348
rect 89916 689284 89917 689348
rect 89851 689283 89917 689284
rect 89854 684450 89914 689283
rect 89486 684390 89914 684450
rect 89486 674797 89546 684390
rect 89483 674796 89549 674797
rect 89483 674732 89484 674796
rect 89548 674732 89549 674796
rect 89483 674731 89549 674732
rect 89483 665276 89549 665277
rect 89483 665212 89484 665276
rect 89548 665212 89549 665276
rect 89483 665211 89549 665212
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 89486 655485 89546 665211
rect 89483 655484 89549 655485
rect 89483 655420 89484 655484
rect 89548 655420 89549 655484
rect 89483 655419 89549 655420
rect 89483 645964 89549 645965
rect 89483 645900 89484 645964
rect 89548 645900 89549 645964
rect 89483 645899 89549 645900
rect 89486 636173 89546 645899
rect 89483 636172 89549 636173
rect 89483 636108 89484 636172
rect 89548 636108 89549 636172
rect 89483 636107 89549 636108
rect 89483 626652 89549 626653
rect 89483 626588 89484 626652
rect 89548 626588 89549 626652
rect 89483 626587 89549 626588
rect 89486 626517 89546 626587
rect 89299 626516 89365 626517
rect 89299 626452 89300 626516
rect 89364 626452 89365 626516
rect 89299 626451 89365 626452
rect 89483 626516 89549 626517
rect 89483 626452 89484 626516
rect 89548 626452 89549 626516
rect 89483 626451 89549 626452
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 89302 617130 89362 626451
rect 89302 617070 89546 617130
rect 89486 596189 89546 617070
rect 89483 596188 89549 596189
rect 89483 596124 89484 596188
rect 89548 596124 89549 596188
rect 89483 596123 89549 596124
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 582000 84204 588698
rect 87643 585716 87709 585717
rect 87643 585652 87644 585716
rect 87708 585652 87709 585716
rect 87643 585651 87709 585652
rect 87275 584356 87341 584357
rect 87275 584292 87276 584356
rect 87340 584292 87341 584356
rect 87275 584291 87341 584292
rect 84515 583948 84581 583949
rect 84515 583884 84516 583948
rect 84580 583884 84581 583948
rect 84515 583883 84581 583884
rect 84331 581500 84397 581501
rect 84331 581436 84332 581500
rect 84396 581436 84397 581500
rect 84331 581435 84397 581436
rect 83779 581228 83845 581229
rect 83779 581164 83780 581228
rect 83844 581164 83845 581228
rect 83779 581163 83845 581164
rect 82307 580956 82373 580957
rect 82307 580892 82308 580956
rect 82372 580892 82373 580956
rect 82307 580891 82373 580892
rect 82310 570298 82370 580891
rect 83782 579050 83842 581163
rect 83046 578990 83842 579050
rect 82678 569618 82738 574822
rect 83046 570074 83106 578990
rect 84334 577690 84394 581435
rect 83782 577630 84394 577690
rect 83782 575058 83842 577630
rect 84518 575650 84578 583883
rect 84699 582996 84765 582997
rect 84699 582932 84700 582996
rect 84764 582932 84765 582996
rect 84699 582931 84765 582932
rect 84334 575590 84578 575650
rect 84334 574290 84394 575590
rect 84702 574970 84762 582931
rect 86723 582452 86789 582453
rect 86723 582388 86724 582452
rect 86788 582388 86789 582452
rect 86723 582387 86789 582388
rect 85251 582044 85317 582045
rect 85251 581980 85252 582044
rect 85316 581980 85317 582044
rect 85251 581979 85317 581980
rect 84883 581908 84949 581909
rect 84883 581844 84884 581908
rect 84948 581844 84949 581908
rect 84883 581843 84949 581844
rect 83782 574230 84394 574290
rect 84518 574910 84762 574970
rect 83782 571570 83842 574230
rect 84150 572250 84210 573462
rect 84518 572930 84578 574910
rect 84886 573698 84946 581843
rect 84518 572870 85130 572930
rect 84150 572190 84946 572250
rect 83782 571510 84210 571570
rect 84150 570074 84210 571510
rect 83046 570014 83842 570074
rect 84150 570014 84762 570074
rect 83414 563410 83474 565302
rect 83782 564770 83842 570014
rect 83782 564710 84026 564770
rect 83414 563350 83658 563410
rect 83598 559418 83658 563350
rect 83966 558650 84026 564710
rect 84334 561370 84394 569382
rect 83414 558590 84026 558650
rect 84150 561310 84394 561370
rect 82491 551852 82557 551853
rect 82491 551788 82492 551852
rect 82556 551850 82557 551852
rect 82556 551790 82922 551850
rect 82556 551788 82557 551790
rect 82491 551787 82557 551788
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 81387 545324 81453 545325
rect 81387 545260 81388 545324
rect 81452 545260 81453 545324
rect 82862 545322 82922 551790
rect 81387 545259 81453 545260
rect 82494 545262 82922 545322
rect 81203 531180 81269 531181
rect 81203 531116 81204 531180
rect 81268 531116 81269 531180
rect 81203 531115 81269 531116
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80838 487338 80898 504782
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80838 418658 80898 420462
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80838 393141 80898 393262
rect 80835 393140 80901 393141
rect 80835 393076 80836 393140
rect 80900 393076 80901 393140
rect 80835 393075 80901 393076
rect 80835 387020 80901 387021
rect 80835 386956 80836 387020
rect 80900 386956 80901 387020
rect 80835 386955 80901 386956
rect 80838 386018 80898 386955
rect 80835 385660 80901 385661
rect 80835 385596 80836 385660
rect 80900 385596 80901 385660
rect 80835 385595 80901 385596
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80838 356778 80898 385595
rect 80838 349978 80898 353822
rect 80838 346578 80898 349062
rect 80835 338060 80901 338061
rect 80835 337996 80836 338060
rect 80900 337996 80901 338060
rect 80835 337995 80901 337996
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80838 328898 80898 337995
rect 80835 327860 80901 327861
rect 80835 327796 80836 327860
rect 80900 327796 80901 327860
rect 80835 327795 80901 327796
rect 80838 313258 80898 327795
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80838 293453 80898 299422
rect 81019 298892 81085 298893
rect 81019 298828 81020 298892
rect 81084 298828 81085 298892
rect 81019 298827 81085 298828
rect 80835 293452 80901 293453
rect 80835 293388 80836 293452
rect 80900 293388 80901 293452
rect 80835 293387 80901 293388
rect 80835 270604 80901 270605
rect 80835 270540 80836 270604
rect 80900 270540 80901 270604
rect 80835 270539 80901 270540
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 237098 80604 261098
rect 80838 241365 80898 270539
rect 81022 241501 81082 298827
rect 81019 241500 81085 241501
rect 81019 241436 81020 241500
rect 81084 241436 81085 241500
rect 81019 241435 81085 241436
rect 81206 241365 81266 531115
rect 81390 241365 81450 545259
rect 81571 538252 81637 538253
rect 81571 538188 81572 538252
rect 81636 538188 81637 538252
rect 81571 538187 81637 538188
rect 80835 241364 80901 241365
rect 80835 241300 80836 241364
rect 80900 241300 80901 241364
rect 80835 241299 80901 241300
rect 81203 241364 81269 241365
rect 81203 241300 81204 241364
rect 81268 241300 81269 241364
rect 81203 241299 81269 241300
rect 81387 241364 81453 241365
rect 81387 241300 81388 241364
rect 81452 241300 81453 241364
rect 81387 241299 81453 241300
rect 80835 240820 80901 240821
rect 80835 240756 80836 240820
rect 80900 240756 80901 240820
rect 80835 240755 80901 240756
rect 81203 240820 81269 240821
rect 81203 240756 81204 240820
rect 81268 240756 81269 240820
rect 81203 240755 81269 240756
rect 81387 240820 81453 240821
rect 81387 240756 81388 240820
rect 81452 240756 81453 240820
rect 81387 240755 81453 240756
rect 80004 236862 80198 237098
rect 80434 236862 80604 237098
rect 80004 225654 80604 236862
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80838 137461 80898 240755
rect 81019 239460 81085 239461
rect 81019 239396 81020 239460
rect 81084 239396 81085 239460
rect 81019 239395 81085 239396
rect 80835 137460 80901 137461
rect 80835 137396 80836 137460
rect 80900 137396 80901 137460
rect 80835 137395 80901 137396
rect 80835 137324 80901 137325
rect 80835 137260 80836 137324
rect 80900 137260 80901 137324
rect 80835 137259 80901 137260
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 79731 10572 79797 10573
rect 79731 10508 79732 10572
rect 79796 10508 79797 10572
rect 79731 10507 79797 10508
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 79547 6356 79613 6357
rect 79547 6292 79548 6356
rect 79612 6292 79613 6356
rect 79547 6291 79613 6292
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 -4026 80604 9098
rect 80838 3365 80898 137259
rect 81022 14517 81082 239395
rect 81206 111077 81266 240755
rect 81203 111076 81269 111077
rect 81203 111012 81204 111076
rect 81268 111012 81269 111076
rect 81203 111011 81269 111012
rect 81019 14516 81085 14517
rect 81019 14452 81020 14516
rect 81084 14452 81085 14516
rect 81019 14451 81085 14452
rect 81390 6493 81450 240755
rect 81574 10437 81634 538187
rect 81755 527644 81821 527645
rect 81755 527580 81756 527644
rect 81820 527580 81821 527644
rect 81755 527579 81821 527580
rect 81758 11661 81818 527579
rect 82494 525330 82554 545262
rect 83414 545050 83474 558590
rect 84150 557970 84210 561310
rect 84702 560690 84762 570014
rect 83598 557910 84210 557970
rect 84334 560630 84762 560690
rect 83598 549810 83658 557910
rect 84334 549810 84394 560630
rect 83598 549750 84210 549810
rect 84334 549750 84762 549810
rect 84150 547090 84210 549750
rect 84702 549130 84762 549750
rect 82678 544990 83474 545050
rect 83598 547030 84210 547090
rect 84334 549070 84762 549130
rect 82678 539613 82738 544990
rect 83598 543778 83658 547030
rect 84334 544370 84394 549070
rect 84886 546410 84946 572190
rect 83966 544310 84394 544370
rect 84702 546350 84946 546410
rect 84702 544370 84762 546350
rect 84702 544310 84946 544370
rect 83966 543010 84026 544310
rect 82629 539612 82738 539613
rect 82629 539548 82630 539612
rect 82694 539550 82738 539612
rect 83046 542950 84026 543010
rect 82694 539548 82695 539550
rect 82629 539547 82695 539548
rect 83046 536890 83106 542950
rect 84150 537658 84210 539462
rect 83046 536830 83290 536890
rect 83230 536210 83290 536830
rect 82862 536150 83290 536210
rect 82862 534850 82922 536150
rect 83414 535530 83474 537422
rect 84518 536298 84578 543542
rect 83414 535470 83658 535530
rect 82862 534790 83290 534850
rect 82862 526690 82922 529942
rect 83230 527370 83290 534790
rect 83598 530090 83658 535470
rect 83782 530770 83842 536062
rect 84886 535530 84946 544310
rect 84150 535470 84946 535530
rect 84150 531450 84210 535470
rect 84150 531390 84946 531450
rect 83782 530710 84394 530770
rect 83598 530030 83842 530090
rect 83230 527310 83474 527370
rect 82862 526630 83290 526690
rect 82494 525270 82922 525330
rect 82491 523836 82557 523837
rect 82491 523772 82492 523836
rect 82556 523772 82557 523836
rect 82491 523771 82557 523772
rect 82494 519349 82554 523771
rect 82862 521250 82922 525270
rect 82678 521190 82922 521250
rect 82491 519348 82557 519349
rect 82491 519284 82492 519348
rect 82556 519284 82557 519348
rect 82491 519283 82557 519284
rect 82491 519076 82557 519077
rect 82491 519012 82492 519076
rect 82556 519012 82557 519076
rect 82491 519011 82557 519012
rect 82494 518805 82554 519011
rect 82491 518804 82557 518805
rect 82491 518740 82492 518804
rect 82556 518740 82557 518804
rect 82678 518802 82738 521190
rect 83230 519298 83290 526630
rect 83414 526010 83474 527310
rect 83782 526690 83842 530030
rect 84334 527370 84394 530710
rect 84334 527310 84762 527370
rect 83782 526630 84578 526690
rect 83414 525950 84394 526010
rect 84334 518802 84394 525950
rect 82678 518742 82922 518802
rect 82491 518739 82557 518740
rect 82307 509556 82373 509557
rect 82307 509492 82308 509556
rect 82372 509492 82373 509556
rect 82307 509491 82373 509492
rect 82310 501530 82370 509491
rect 82494 505749 82554 515662
rect 82862 513770 82922 518742
rect 84150 518742 84394 518802
rect 84150 515898 84210 518742
rect 84518 515130 84578 526630
rect 82678 513710 82922 513770
rect 84150 515070 84578 515130
rect 82491 505748 82557 505749
rect 82491 505684 82492 505748
rect 82556 505684 82557 505748
rect 82491 505683 82557 505684
rect 82678 504338 82738 513710
rect 84150 510234 84210 515070
rect 84702 514450 84762 527310
rect 84334 514390 84762 514450
rect 84334 511050 84394 514390
rect 84334 510990 84762 511050
rect 83782 510174 84210 510234
rect 83782 505018 83842 510174
rect 84702 509690 84762 510990
rect 84518 509630 84762 509690
rect 84518 508330 84578 509630
rect 84886 509554 84946 531390
rect 84150 508270 84578 508330
rect 84702 509494 84946 509554
rect 82310 501470 82738 501530
rect 82307 497180 82373 497181
rect 82307 497116 82308 497180
rect 82372 497116 82373 497180
rect 82307 497115 82373 497116
rect 82310 496858 82370 497115
rect 82123 495820 82189 495821
rect 82123 495756 82124 495820
rect 82188 495756 82189 495820
rect 82123 495755 82189 495756
rect 81939 492012 82005 492013
rect 81939 491948 81940 492012
rect 82004 491948 82005 492012
rect 81939 491947 82005 491948
rect 81755 11660 81821 11661
rect 81755 11596 81756 11660
rect 81820 11596 81821 11660
rect 81755 11595 81821 11596
rect 81571 10436 81637 10437
rect 81571 10372 81572 10436
rect 81636 10372 81637 10436
rect 81571 10371 81637 10372
rect 81387 6492 81453 6493
rect 81387 6428 81388 6492
rect 81452 6428 81453 6492
rect 81387 6427 81453 6428
rect 81942 6221 82002 491947
rect 82126 170645 82186 495755
rect 82678 487930 82738 501470
rect 83230 489290 83290 504102
rect 84150 502890 84210 508270
rect 84702 504930 84762 509494
rect 85070 504930 85130 572870
rect 83598 502830 84210 502890
rect 84518 504870 84762 504930
rect 84886 504870 85130 504930
rect 83598 501618 83658 502830
rect 82494 487870 82738 487930
rect 82862 489230 83290 489290
rect 82494 487250 82554 487870
rect 82310 487190 82554 487250
rect 82310 479770 82370 487190
rect 82491 486164 82557 486165
rect 82491 486100 82492 486164
rect 82556 486100 82557 486164
rect 82491 486099 82557 486100
rect 82494 485890 82554 486099
rect 82862 485890 82922 489230
rect 82494 485830 82922 485890
rect 83230 485890 83290 487102
rect 83230 485830 83658 485890
rect 82491 484940 82557 484941
rect 82491 484876 82492 484940
rect 82556 484876 82557 484940
rect 82491 484875 82557 484876
rect 82494 481269 82554 484875
rect 82491 481268 82557 481269
rect 82491 481204 82492 481268
rect 82556 481204 82557 481268
rect 82491 481203 82557 481204
rect 82491 481132 82557 481133
rect 82491 481068 82492 481132
rect 82556 481130 82557 481132
rect 82556 481070 82922 481130
rect 82556 481068 82557 481070
rect 82491 481067 82557 481068
rect 82310 479710 82554 479770
rect 82494 475829 82554 479710
rect 82491 475828 82557 475829
rect 82491 475764 82492 475828
rect 82556 475764 82557 475828
rect 82491 475763 82557 475764
rect 82862 474330 82922 481070
rect 82494 474270 82922 474330
rect 82494 474197 82554 474270
rect 82491 474196 82557 474197
rect 82491 474132 82492 474196
rect 82556 474132 82557 474196
rect 82491 474131 82557 474132
rect 82491 473652 82557 473653
rect 82491 473588 82492 473652
rect 82556 473650 82557 473652
rect 82556 473590 82738 473650
rect 82556 473588 82557 473590
rect 82491 473587 82557 473588
rect 82491 473516 82557 473517
rect 82491 473452 82492 473516
rect 82556 473452 82557 473516
rect 82491 473451 82557 473452
rect 82494 471069 82554 473451
rect 82678 472290 82738 473590
rect 83230 473058 83290 481662
rect 83598 472970 83658 485830
rect 83782 477050 83842 500702
rect 84518 498810 84578 504870
rect 84886 504250 84946 504870
rect 84886 504190 85130 504250
rect 84518 498750 84946 498810
rect 84334 493370 84394 497982
rect 83966 493310 84394 493370
rect 83966 492010 84026 493310
rect 84334 492010 84394 492542
rect 83966 491950 84210 492010
rect 84334 491950 84578 492010
rect 84150 485890 84210 491950
rect 84518 486658 84578 491950
rect 84150 485830 84578 485890
rect 84518 479858 84578 485830
rect 83782 476990 84394 477050
rect 83598 472910 84026 472970
rect 82678 472230 83474 472290
rect 82491 471068 82557 471069
rect 82491 471004 82492 471068
rect 82556 471004 82557 471068
rect 82491 471003 82557 471004
rect 83414 468978 83474 472230
rect 82491 466172 82557 466173
rect 82491 466108 82492 466172
rect 82556 466170 82557 466172
rect 82556 466110 83290 466170
rect 82556 466108 82557 466110
rect 82491 466107 82557 466108
rect 83230 462090 83290 466110
rect 83414 465490 83474 467382
rect 83414 465430 83658 465490
rect 83230 462030 83474 462090
rect 82491 458012 82557 458013
rect 82491 457948 82492 458012
rect 82556 458010 82557 458012
rect 82556 457950 82738 458010
rect 82556 457948 82557 457950
rect 82491 457947 82557 457948
rect 82307 456924 82373 456925
rect 82307 456860 82308 456924
rect 82372 456860 82373 456924
rect 82307 456859 82373 456860
rect 82310 407010 82370 456859
rect 82491 438972 82557 438973
rect 82491 438908 82492 438972
rect 82556 438970 82557 438972
rect 82678 438970 82738 457950
rect 83414 457330 83474 462030
rect 82556 438910 82738 438970
rect 82862 457270 83474 457330
rect 82556 438908 82557 438910
rect 82491 438907 82557 438908
rect 82491 435436 82557 435437
rect 82491 435372 82492 435436
rect 82556 435372 82557 435436
rect 82491 435371 82557 435372
rect 82494 431221 82554 435371
rect 82491 431220 82557 431221
rect 82491 431156 82492 431220
rect 82556 431156 82557 431220
rect 82491 431155 82557 431156
rect 82310 406950 82738 407010
rect 82491 406468 82557 406469
rect 82491 406404 82492 406468
rect 82556 406404 82557 406468
rect 82491 406403 82557 406404
rect 82494 401573 82554 406403
rect 82491 401572 82557 401573
rect 82491 401508 82492 401572
rect 82556 401508 82557 401572
rect 82491 401507 82557 401508
rect 82491 400212 82557 400213
rect 82491 400148 82492 400212
rect 82556 400210 82557 400212
rect 82678 400210 82738 406950
rect 82556 400150 82738 400210
rect 82556 400148 82557 400150
rect 82491 400147 82557 400148
rect 82862 399530 82922 457270
rect 83598 455970 83658 465430
rect 83598 455910 83842 455970
rect 83782 433530 83842 455910
rect 83598 433470 83842 433530
rect 83598 404290 83658 433470
rect 83966 420698 84026 472910
rect 84334 465490 84394 476990
rect 84150 465430 84394 465490
rect 84150 455970 84210 465430
rect 84518 458010 84578 478942
rect 84334 457950 84578 458010
rect 84334 456922 84394 457950
rect 84334 456862 84762 456922
rect 84150 455910 84394 455970
rect 84334 442370 84394 455910
rect 84334 442310 84578 442370
rect 84518 434210 84578 442310
rect 84150 434150 84578 434210
rect 84150 427410 84210 434150
rect 84150 427350 84578 427410
rect 84150 414490 84210 418422
rect 84518 417890 84578 427350
rect 83414 404230 83658 404290
rect 83966 414430 84210 414490
rect 84334 417830 84578 417890
rect 83414 403698 83474 404230
rect 83966 402930 84026 414430
rect 83230 402870 84026 402930
rect 83230 402250 83290 402870
rect 82678 399470 82922 399530
rect 83046 402190 83290 402250
rect 82678 396898 82738 399470
rect 82491 396132 82557 396133
rect 82491 396068 82492 396132
rect 82556 396130 82557 396132
rect 82556 396070 82738 396130
rect 82556 396068 82557 396070
rect 82491 396067 82557 396068
rect 82307 394092 82373 394093
rect 82307 394028 82308 394092
rect 82372 394028 82373 394092
rect 82307 394027 82373 394028
rect 82310 390010 82370 394027
rect 82678 393410 82738 396070
rect 83046 394178 83106 402190
rect 84334 401570 84394 417830
rect 83966 401510 84394 401570
rect 83414 395450 83474 396662
rect 83414 395390 83658 395450
rect 82494 393350 82738 393410
rect 82494 391237 82554 393350
rect 83598 392818 83658 395390
rect 82491 391236 82557 391237
rect 82491 391172 82492 391236
rect 82556 391172 82557 391236
rect 82491 391171 82557 391172
rect 82310 389950 82922 390010
rect 82491 385796 82557 385797
rect 82491 385732 82492 385796
rect 82556 385732 82557 385796
rect 82491 385731 82557 385732
rect 82307 385660 82373 385661
rect 82307 385596 82308 385660
rect 82372 385596 82373 385660
rect 82307 385595 82373 385596
rect 82310 369069 82370 385595
rect 82494 371925 82554 385731
rect 82862 377858 82922 389950
rect 83046 382530 83106 392582
rect 83966 392050 84026 401510
rect 83598 391990 84026 392050
rect 83046 382470 83290 382530
rect 83230 375730 83290 382470
rect 83598 378450 83658 391990
rect 84702 390010 84762 456862
rect 84334 389950 84762 390010
rect 84334 384570 84394 389950
rect 84150 384510 84394 384570
rect 84150 382618 84210 384510
rect 84886 383482 84946 498750
rect 84702 383422 84946 383482
rect 84702 380490 84762 383422
rect 85070 383210 85130 504190
rect 84886 383150 85130 383210
rect 84886 381850 84946 383150
rect 84886 381790 85130 381850
rect 84702 380430 84946 380490
rect 83598 378390 84210 378450
rect 83046 375670 83290 375730
rect 83046 374370 83106 375670
rect 82862 374310 83106 374370
rect 82491 371924 82557 371925
rect 82491 371860 82492 371924
rect 82556 371860 82557 371924
rect 82491 371859 82557 371860
rect 82307 369068 82373 369069
rect 82307 369004 82308 369068
rect 82372 369004 82373 369068
rect 82307 369003 82373 369004
rect 82307 368932 82373 368933
rect 82307 368868 82308 368932
rect 82372 368868 82373 368932
rect 82862 368930 82922 374310
rect 82307 368867 82373 368868
rect 82494 368870 82922 368930
rect 82310 368658 82370 368867
rect 82494 368797 82554 368870
rect 82491 368796 82557 368797
rect 82491 368732 82492 368796
rect 82556 368732 82557 368796
rect 82491 368731 82557 368732
rect 82310 368598 83290 368658
rect 82491 368116 82557 368117
rect 82491 368052 82492 368116
rect 82556 368052 82557 368116
rect 82491 368051 82557 368052
rect 82494 366210 82554 368051
rect 82310 366150 82554 366210
rect 82310 362130 82370 366150
rect 82491 364852 82557 364853
rect 82491 364788 82492 364852
rect 82556 364850 82557 364852
rect 82862 364850 82922 367422
rect 83230 366210 83290 368598
rect 83782 367658 83842 377622
rect 84150 377178 84210 378390
rect 84150 375730 84210 376262
rect 83966 375670 84210 375730
rect 83966 373010 84026 375670
rect 83966 372950 84210 373010
rect 82556 364790 82922 364850
rect 83046 366150 83290 366210
rect 82556 364788 82557 364790
rect 82491 364787 82557 364788
rect 82491 364716 82557 364717
rect 82491 364652 82492 364716
rect 82556 364652 82557 364716
rect 82491 364651 82557 364652
rect 82494 362949 82554 364651
rect 82491 362948 82557 362949
rect 82491 362884 82492 362948
rect 82556 362884 82557 362948
rect 82491 362883 82557 362884
rect 82491 362812 82557 362813
rect 82491 362748 82492 362812
rect 82556 362810 82557 362812
rect 82556 362750 82922 362810
rect 82556 362748 82557 362750
rect 82491 362747 82557 362748
rect 82310 362070 82738 362130
rect 82307 360228 82373 360229
rect 82307 360164 82308 360228
rect 82372 360164 82373 360228
rect 82678 360226 82738 362070
rect 82307 360163 82373 360164
rect 82494 360166 82738 360226
rect 82310 339013 82370 360163
rect 82494 347037 82554 360166
rect 82629 360092 82695 360093
rect 82629 360028 82630 360092
rect 82694 360090 82695 360092
rect 82862 360090 82922 362750
rect 82694 360030 82922 360090
rect 82694 360028 82695 360030
rect 82629 360027 82695 360028
rect 83046 359498 83106 366150
rect 84150 365530 84210 372950
rect 84518 367570 84578 375582
rect 84518 367510 84762 367570
rect 84702 366890 84762 367510
rect 83598 365470 84210 365530
rect 84334 366830 84762 366890
rect 82629 359412 82695 359413
rect 82629 359348 82630 359412
rect 82694 359410 82695 359412
rect 82694 359348 82738 359410
rect 82629 359347 82738 359348
rect 82678 358730 82738 359347
rect 83598 359410 83658 365470
rect 84334 364850 84394 366830
rect 83782 364790 84394 364850
rect 83782 360090 83842 364790
rect 84886 362130 84946 380430
rect 84702 362070 84946 362130
rect 83782 360030 84394 360090
rect 83598 359350 84210 359410
rect 82678 358670 84026 358730
rect 82629 358052 82695 358053
rect 82629 357988 82630 358052
rect 82694 358050 82695 358052
rect 82694 357990 83106 358050
rect 82694 357988 82695 357990
rect 82629 357987 82695 357988
rect 83046 357778 83106 357990
rect 83046 357718 83290 357778
rect 82632 357310 82774 357370
rect 82632 356418 82692 357310
rect 83230 356418 83290 357718
rect 82632 356358 82738 356418
rect 82678 353970 82738 356358
rect 82862 356358 83290 356418
rect 82862 354650 82922 356358
rect 82862 354590 83290 354650
rect 82678 353910 82922 353970
rect 82862 353378 82922 353910
rect 83230 350570 83290 354590
rect 83598 354058 83658 356270
rect 82862 350510 83290 350570
rect 82491 347036 82557 347037
rect 82491 346972 82492 347036
rect 82556 346972 82557 347036
rect 82491 346971 82557 346972
rect 82629 341732 82695 341733
rect 82629 341668 82630 341732
rect 82694 341730 82695 341732
rect 82862 341730 82922 350510
rect 82694 341670 82922 341730
rect 82694 341668 82695 341670
rect 82629 341667 82695 341668
rect 82491 339692 82557 339693
rect 82491 339628 82492 339692
rect 82556 339690 82557 339692
rect 82678 339690 82738 340902
rect 82556 339630 82738 339690
rect 82556 339628 82557 339630
rect 82491 339627 82557 339628
rect 82307 339012 82373 339013
rect 82307 338948 82308 339012
rect 82372 338948 82373 339012
rect 82307 338947 82373 338948
rect 82491 336836 82557 336837
rect 82491 336772 82492 336836
rect 82556 336772 82557 336836
rect 82491 336771 82557 336772
rect 82494 335069 82554 336771
rect 82491 335068 82557 335069
rect 82491 335004 82492 335068
rect 82556 335004 82557 335068
rect 82491 335003 82557 335004
rect 83230 331618 83290 349742
rect 83598 341138 83658 353142
rect 83966 334930 84026 358670
rect 83598 334870 84026 334930
rect 82307 331260 82373 331261
rect 82307 331196 82308 331260
rect 82372 331196 82373 331260
rect 82307 331195 82373 331196
rect 82491 331260 82557 331261
rect 82491 331196 82492 331260
rect 82556 331258 82557 331260
rect 82556 331198 82738 331258
rect 82556 331196 82557 331198
rect 82491 331195 82557 331196
rect 82310 316570 82370 331195
rect 82491 331124 82557 331125
rect 82491 331060 82492 331124
rect 82556 331060 82557 331124
rect 82491 331059 82557 331060
rect 82494 317389 82554 331059
rect 82678 320650 82738 331198
rect 83598 330850 83658 334870
rect 84150 332890 84210 359350
rect 84334 346490 84394 360030
rect 84702 349298 84762 362070
rect 84334 346430 84946 346490
rect 84518 343178 84578 345662
rect 84886 340370 84946 346430
rect 83966 332830 84210 332890
rect 84334 340310 84946 340370
rect 83966 332298 84026 332830
rect 83046 330790 83658 330850
rect 83046 321418 83106 330790
rect 83414 320650 83474 328662
rect 83782 322098 83842 327982
rect 84334 327858 84394 340310
rect 84850 339630 84946 339690
rect 84334 327798 84762 327858
rect 84334 322778 84394 327302
rect 84702 322010 84762 327798
rect 84150 321950 84762 322010
rect 82678 320590 82922 320650
rect 82491 317388 82557 317389
rect 82491 317324 82492 317388
rect 82556 317324 82557 317388
rect 82491 317323 82557 317324
rect 82310 316510 82738 316570
rect 82491 316300 82557 316301
rect 82491 316236 82492 316300
rect 82556 316236 82557 316300
rect 82491 316235 82557 316236
rect 82494 312357 82554 316235
rect 82491 312356 82557 312357
rect 82491 312292 82492 312356
rect 82556 312292 82557 312356
rect 82491 312291 82557 312292
rect 82491 307460 82557 307461
rect 82491 307396 82492 307460
rect 82556 307396 82557 307460
rect 82491 307395 82557 307396
rect 82494 297805 82554 307395
rect 82491 297804 82557 297805
rect 82491 297740 82492 297804
rect 82556 297740 82557 297804
rect 82491 297739 82557 297740
rect 82491 297532 82557 297533
rect 82491 297468 82492 297532
rect 82556 297530 82557 297532
rect 82678 297530 82738 316510
rect 82556 297470 82738 297530
rect 82556 297468 82557 297470
rect 82491 297467 82557 297468
rect 82491 296852 82557 296853
rect 82491 296788 82492 296852
rect 82556 296850 82557 296852
rect 82862 296850 82922 320590
rect 83230 320590 83474 320650
rect 83230 318610 83290 320590
rect 83782 319290 83842 321182
rect 83782 319230 84026 319290
rect 83230 318550 83658 318610
rect 83230 308410 83290 313022
rect 83230 308350 83474 308410
rect 83414 300250 83474 308350
rect 82556 296790 82922 296850
rect 83230 300190 83474 300250
rect 82556 296788 82557 296790
rect 82491 296787 82557 296788
rect 83230 295578 83290 300190
rect 83598 299658 83658 318550
rect 83598 294130 83658 298742
rect 83966 294898 84026 319230
rect 84150 299570 84210 321950
rect 84666 321270 84762 321330
rect 84702 307458 84762 321270
rect 84518 307398 84762 307458
rect 84518 303058 84578 307398
rect 84518 300250 84578 302142
rect 84518 300190 84762 300250
rect 84150 299510 84578 299570
rect 84518 298210 84578 299510
rect 84150 298150 84578 298210
rect 84150 295490 84210 298150
rect 84702 296170 84762 300190
rect 84666 296110 84762 296170
rect 84150 295430 84578 295490
rect 83598 294070 84210 294130
rect 82491 293452 82557 293453
rect 82491 293388 82492 293452
rect 82556 293450 82557 293452
rect 82556 293390 83842 293450
rect 82556 293388 82557 293390
rect 82491 293387 82557 293388
rect 82491 292092 82557 292093
rect 82491 292028 82492 292092
rect 82556 292090 82557 292092
rect 82556 292030 82738 292090
rect 82556 292028 82557 292030
rect 82491 292027 82557 292028
rect 82307 291140 82373 291141
rect 82307 291076 82308 291140
rect 82372 291076 82373 291140
rect 82307 291075 82373 291076
rect 82310 280941 82370 291075
rect 82491 289100 82557 289101
rect 82491 289036 82492 289100
rect 82556 289036 82557 289100
rect 82491 289035 82557 289036
rect 82307 280940 82373 280941
rect 82307 280876 82308 280940
rect 82372 280876 82373 280940
rect 82307 280875 82373 280876
rect 82494 254829 82554 289035
rect 82678 266253 82738 292030
rect 83046 283250 83106 292622
rect 83046 283190 83658 283250
rect 83598 279170 83658 283190
rect 83414 279110 83658 279170
rect 83782 279170 83842 293390
rect 84150 290050 84210 294070
rect 84518 293450 84578 295430
rect 83966 289990 84210 290050
rect 84334 293390 84578 293450
rect 83966 280938 84026 289990
rect 84334 284018 84394 293390
rect 84886 287070 84946 339630
rect 84702 287010 84946 287070
rect 84702 281890 84762 287010
rect 84334 281830 84762 281890
rect 84334 281298 84394 281830
rect 84702 281150 84946 281210
rect 84702 280938 84762 281150
rect 83966 280878 84762 280938
rect 84150 279170 84210 279702
rect 83782 279110 84210 279170
rect 83046 273730 83106 276982
rect 82629 266252 82738 266253
rect 82629 266188 82630 266252
rect 82694 266190 82738 266252
rect 82862 273670 83106 273730
rect 82694 266188 82695 266190
rect 82629 266187 82695 266188
rect 82862 265570 82922 273670
rect 83414 270330 83474 279110
rect 84518 277810 84578 280382
rect 84518 277750 84762 277810
rect 84298 277350 84578 277410
rect 84518 275770 84578 277350
rect 84150 275710 84578 275770
rect 84150 273730 84210 275710
rect 84702 275090 84762 277750
rect 83598 273670 84210 273730
rect 84334 275030 84762 275090
rect 83598 270602 83658 273670
rect 83966 271690 84026 272902
rect 84334 272370 84394 275030
rect 84886 274410 84946 281150
rect 84702 274350 84946 274410
rect 84702 273818 84762 274350
rect 84334 272310 84946 272370
rect 83966 271630 84210 271690
rect 84150 270602 84210 271630
rect 83598 270542 84026 270602
rect 84150 270542 84394 270602
rect 83966 270330 84026 270542
rect 83414 270270 83842 270330
rect 83966 270270 84210 270330
rect 83414 266338 83474 269502
rect 82678 265510 82922 265570
rect 82678 262853 82738 265510
rect 83782 264890 83842 270270
rect 82629 262852 82738 262853
rect 82629 262788 82630 262852
rect 82694 262790 82738 262852
rect 82862 264830 83842 264890
rect 82694 262788 82695 262790
rect 82629 262787 82695 262788
rect 82629 260812 82695 260813
rect 82629 260748 82630 260812
rect 82694 260810 82695 260812
rect 82862 260810 82922 264830
rect 82694 260750 82922 260810
rect 82694 260748 82695 260750
rect 82629 260747 82695 260748
rect 82629 260268 82695 260269
rect 82629 260204 82630 260268
rect 82694 260266 82695 260268
rect 82694 260204 82738 260266
rect 82629 260203 82738 260204
rect 82491 254828 82557 254829
rect 82491 254764 82492 254828
rect 82556 254764 82557 254828
rect 82491 254763 82557 254764
rect 82678 254690 82738 260203
rect 83046 255458 83106 259982
rect 83414 259450 83474 264062
rect 84150 260810 84210 270270
rect 83598 260750 84210 260810
rect 83598 260130 83658 260750
rect 83598 260070 84026 260130
rect 83966 259450 84026 260070
rect 84334 259450 84394 270542
rect 83230 259390 83474 259450
rect 83598 259390 84026 259450
rect 84150 259390 84394 259450
rect 83230 256730 83290 259390
rect 83598 256730 83658 259390
rect 84150 258858 84210 259390
rect 83230 256670 83474 256730
rect 83598 256670 84210 256730
rect 82310 254630 82738 254690
rect 82310 252922 82370 254630
rect 82491 254012 82557 254013
rect 82491 253948 82492 254012
rect 82556 254010 82557 254012
rect 83414 254010 83474 256670
rect 82556 253950 83474 254010
rect 82556 253948 82557 253950
rect 82491 253947 82557 253948
rect 83782 253330 83842 255222
rect 84150 254690 84210 256670
rect 84518 254690 84578 270862
rect 82862 253270 83842 253330
rect 83966 254630 84210 254690
rect 84334 254630 84578 254690
rect 82310 252862 82738 252922
rect 82491 252788 82557 252789
rect 82491 252724 82492 252788
rect 82556 252724 82557 252788
rect 82491 252723 82557 252724
rect 82494 239594 82554 252723
rect 82310 239534 82554 239594
rect 82310 232661 82370 239534
rect 82537 239460 82603 239461
rect 82537 239396 82538 239460
rect 82602 239458 82603 239460
rect 82678 239458 82738 252862
rect 82602 239398 82738 239458
rect 82602 239396 82603 239398
rect 82537 239395 82603 239396
rect 82491 238372 82557 238373
rect 82491 238308 82492 238372
rect 82556 238370 82557 238372
rect 82862 238370 82922 253270
rect 83230 252738 83658 252786
rect 83230 252726 83510 252738
rect 83230 246530 83290 252726
rect 83966 247978 84026 254630
rect 84334 252786 84394 254630
rect 84334 252726 84762 252786
rect 83230 246470 84578 246530
rect 82556 238310 82922 238370
rect 82556 238308 82557 238310
rect 82491 238307 82557 238308
rect 82491 237012 82557 237013
rect 82491 236948 82492 237012
rect 82556 237010 82557 237012
rect 82862 237010 82922 237542
rect 82556 236950 82922 237010
rect 82556 236948 82557 236950
rect 82491 236947 82557 236948
rect 83230 236330 83290 242302
rect 83598 238458 83658 241622
rect 83966 237690 84026 245022
rect 82862 236270 83290 236330
rect 83598 237630 84026 237690
rect 82491 236196 82557 236197
rect 82491 236132 82492 236196
rect 82556 236132 82557 236196
rect 82491 236131 82557 236132
rect 82494 235874 82554 236131
rect 82491 235108 82557 235109
rect 82491 235044 82492 235108
rect 82556 235044 82557 235108
rect 82491 235043 82557 235044
rect 82494 234970 82554 235043
rect 82862 234970 82922 236270
rect 82494 234910 82922 234970
rect 82491 234836 82557 234837
rect 82491 234772 82492 234836
rect 82556 234834 82557 234836
rect 83598 234834 83658 237630
rect 84114 236950 84210 237010
rect 84150 236010 84210 236950
rect 84518 236010 84578 246470
rect 83966 235950 84578 236010
rect 82556 234774 83106 234834
rect 83598 234774 83842 234834
rect 82556 234772 82557 234774
rect 82491 234771 82557 234772
rect 83046 234290 83106 234774
rect 83046 234230 83658 234290
rect 82491 233748 82557 233749
rect 82491 233684 82492 233748
rect 82556 233746 82557 233748
rect 82678 233746 82738 234142
rect 82556 233686 82738 233746
rect 82556 233684 82557 233686
rect 82491 233683 82557 233684
rect 82494 233550 82958 233610
rect 82494 233477 82554 233550
rect 82491 233476 82557 233477
rect 82491 233412 82492 233476
rect 82556 233412 82557 233476
rect 82491 233411 82557 233412
rect 82307 232660 82373 232661
rect 82307 232596 82308 232660
rect 82372 232596 82373 232660
rect 82307 232595 82373 232596
rect 82491 232660 82557 232661
rect 82491 232596 82492 232660
rect 82556 232658 82557 232660
rect 82556 232598 82922 232658
rect 82556 232596 82557 232598
rect 82491 232595 82557 232596
rect 82494 231029 82554 232102
rect 82862 231658 82922 232598
rect 82491 231028 82557 231029
rect 82491 230964 82492 231028
rect 82556 230964 82557 231028
rect 82491 230963 82557 230964
rect 82491 230892 82557 230893
rect 82491 230828 82492 230892
rect 82556 230828 82557 230892
rect 82491 230827 82557 230828
rect 82494 230754 82554 230827
rect 82494 230694 83290 230754
rect 82307 230620 82373 230621
rect 82307 230556 82308 230620
rect 82372 230556 82373 230620
rect 82307 230555 82373 230556
rect 82310 228170 82370 230555
rect 82491 229260 82557 229261
rect 82491 229196 82492 229260
rect 82556 229196 82557 229260
rect 82491 229195 82557 229196
rect 82494 228850 82554 229195
rect 82494 228790 83106 228850
rect 82310 228110 82406 228170
rect 82491 227900 82557 227901
rect 82491 227836 82492 227900
rect 82556 227836 82557 227900
rect 82491 227835 82557 227836
rect 82494 226350 82554 227835
rect 82494 226290 82738 226350
rect 82307 225724 82373 225725
rect 82307 225660 82308 225724
rect 82372 225660 82373 225724
rect 82307 225659 82373 225660
rect 82310 209405 82370 225659
rect 82678 224178 82738 226290
rect 82491 223412 82557 223413
rect 82491 223348 82492 223412
rect 82556 223410 82557 223412
rect 83046 223410 83106 228790
rect 82556 223350 83106 223410
rect 82556 223348 82557 223350
rect 82491 223347 82557 223348
rect 83230 220826 83290 230694
rect 83598 220826 83658 234230
rect 83782 233746 83842 234774
rect 83966 234290 84026 235950
rect 84150 234630 84210 235950
rect 84150 234570 84394 234630
rect 84334 234290 84394 234570
rect 83966 234230 84210 234290
rect 84334 234230 84624 234290
rect 83782 233686 84026 233746
rect 83966 227578 84026 233686
rect 84150 228170 84210 234230
rect 84564 233250 84624 234230
rect 84518 233190 84624 233250
rect 84150 228110 84394 228170
rect 84334 226810 84394 228110
rect 84518 226813 84578 233190
rect 83966 226750 84394 226810
rect 84515 226812 84581 226813
rect 83966 220826 84026 226750
rect 84515 226748 84516 226812
rect 84580 226748 84581 226812
rect 84515 226747 84581 226748
rect 84334 225450 84394 226390
rect 84334 225390 84578 225450
rect 82494 220766 83290 220826
rect 83414 220766 83658 220826
rect 83782 220766 84026 220826
rect 82494 220149 82554 220766
rect 83414 220690 83474 220766
rect 83782 220690 83842 220766
rect 84518 220690 84578 225390
rect 83230 220630 83474 220690
rect 83598 220630 83842 220690
rect 83966 220630 84578 220690
rect 82491 220148 82557 220149
rect 82491 220084 82492 220148
rect 82556 220084 82557 220148
rect 82491 220083 82557 220084
rect 82491 220012 82557 220013
rect 82491 219948 82492 220012
rect 82556 220010 82557 220012
rect 83230 220010 83290 220630
rect 83598 220010 83658 220630
rect 82556 219950 83290 220010
rect 83414 219950 83658 220010
rect 82556 219948 82557 219950
rect 82491 219947 82557 219948
rect 82491 219876 82557 219877
rect 82491 219812 82492 219876
rect 82556 219812 82557 219876
rect 82491 219811 82557 219812
rect 82494 215930 82554 219811
rect 83414 219418 83474 219950
rect 82494 215870 82922 215930
rect 82629 210492 82695 210493
rect 82629 210428 82630 210492
rect 82694 210490 82695 210492
rect 82862 210490 82922 215870
rect 82694 210430 82922 210490
rect 82694 210428 82695 210430
rect 82629 210427 82695 210428
rect 82307 209404 82373 209405
rect 82307 209340 82308 209404
rect 82372 209340 82373 209404
rect 82307 209339 82373 209340
rect 83046 209130 83106 219182
rect 83966 217970 84026 220630
rect 84702 219874 84762 252726
rect 84334 219814 84762 219874
rect 84334 219418 84394 219814
rect 83782 217910 84026 217970
rect 84150 218590 84430 218650
rect 83782 216698 83842 217910
rect 84150 217378 84210 218590
rect 84886 217290 84946 272310
rect 84518 217230 84946 217290
rect 83598 214570 83658 215102
rect 83598 214510 83842 214570
rect 83414 209130 83474 213742
rect 83782 209130 83842 214510
rect 82862 209070 83106 209130
rect 83230 209070 83474 209130
rect 83598 209070 83842 209130
rect 82862 208450 82922 209070
rect 82494 208390 82922 208450
rect 82307 208044 82373 208045
rect 82307 207980 82308 208044
rect 82372 207980 82373 208044
rect 82307 207979 82373 207980
rect 82310 201517 82370 207979
rect 82494 203149 82554 208390
rect 82629 207772 82695 207773
rect 82629 207708 82630 207772
rect 82694 207770 82695 207772
rect 83230 207770 83290 209070
rect 83598 208450 83658 209070
rect 83966 208450 84026 215782
rect 84518 214658 84578 217230
rect 85070 216610 85130 381790
rect 85034 216550 85130 216610
rect 84886 213210 84946 215782
rect 82694 207710 83290 207770
rect 83414 208390 83658 208450
rect 83782 208390 84026 208450
rect 84334 213150 84946 213210
rect 82694 207708 82695 207710
rect 82629 207707 82695 207708
rect 82491 203148 82557 203149
rect 82491 203084 82492 203148
rect 82556 203084 82557 203148
rect 83046 203146 83106 206262
rect 83414 203690 83474 208390
rect 83782 206498 83842 208390
rect 84334 205138 84394 213150
rect 84702 210578 84762 211702
rect 85254 209810 85314 581979
rect 85619 581772 85685 581773
rect 85619 581708 85620 581772
rect 85684 581708 85685 581772
rect 85619 581707 85685 581708
rect 85435 581500 85501 581501
rect 85435 581436 85436 581500
rect 85500 581436 85501 581500
rect 85435 581435 85501 581436
rect 85034 209750 85314 209810
rect 85438 209130 85498 581435
rect 84702 209070 85498 209130
rect 83414 203630 84210 203690
rect 83046 203086 83290 203146
rect 82491 203083 82557 203084
rect 82491 203012 82557 203013
rect 82491 202948 82492 203012
rect 82556 203010 82557 203012
rect 83230 203010 83290 203086
rect 82556 202950 83106 203010
rect 83230 202950 83658 203010
rect 82556 202948 82557 202950
rect 82491 202947 82557 202948
rect 82491 202060 82557 202061
rect 82491 201996 82492 202060
rect 82556 202058 82557 202060
rect 83046 202058 83106 202950
rect 82556 201998 83106 202058
rect 82556 201996 82557 201998
rect 82491 201995 82557 201996
rect 82491 201924 82557 201925
rect 82491 201860 82492 201924
rect 82556 201922 82557 201924
rect 82556 201862 82738 201922
rect 82556 201860 82557 201862
rect 82491 201859 82557 201860
rect 82491 201788 82557 201789
rect 82491 201724 82492 201788
rect 82556 201724 82557 201788
rect 82678 201786 82738 201862
rect 83598 201786 83658 202950
rect 82678 201726 83658 201786
rect 82491 201723 82557 201724
rect 82307 201516 82373 201517
rect 82307 201452 82308 201516
rect 82372 201452 82373 201516
rect 82307 201451 82373 201452
rect 82307 201244 82373 201245
rect 82307 201180 82308 201244
rect 82372 201180 82373 201244
rect 82307 201179 82373 201180
rect 82310 200970 82370 201179
rect 82494 201109 82554 201723
rect 82629 201652 82695 201653
rect 82629 201588 82630 201652
rect 82694 201650 82695 201652
rect 82694 201590 83106 201650
rect 82694 201588 82695 201590
rect 82629 201587 82695 201588
rect 82491 201108 82557 201109
rect 82491 201044 82492 201108
rect 82556 201044 82557 201108
rect 82491 201043 82557 201044
rect 82310 200910 82922 200970
rect 82307 200836 82373 200837
rect 82307 200772 82308 200836
rect 82372 200772 82373 200836
rect 82307 200771 82373 200772
rect 82310 192266 82370 200771
rect 82491 199612 82557 199613
rect 82491 199548 82492 199612
rect 82556 199610 82557 199612
rect 82556 199550 82738 199610
rect 82556 199548 82557 199550
rect 82491 199547 82557 199548
rect 82678 196978 82738 199550
rect 82862 198250 82922 200910
rect 83046 198930 83106 201590
rect 83046 198870 84026 198930
rect 82862 198190 83842 198250
rect 82632 195470 82774 195530
rect 82632 195397 82692 195470
rect 82629 195396 82695 195397
rect 82629 195332 82630 195396
rect 82694 195332 82695 195396
rect 82629 195331 82695 195332
rect 82491 195260 82557 195261
rect 82491 195196 82492 195260
rect 82556 195196 82557 195260
rect 83230 195258 83290 196062
rect 83782 195258 83842 198190
rect 83966 196210 84026 198870
rect 84150 196890 84210 203630
rect 84702 203010 84762 209070
rect 85622 208450 85682 581707
rect 86355 581636 86421 581637
rect 86355 581572 86356 581636
rect 86420 581572 86421 581636
rect 86355 581571 86421 581572
rect 85803 581092 85869 581093
rect 85803 581028 85804 581092
rect 85868 581028 85869 581092
rect 85803 581027 85869 581028
rect 85806 209130 85866 581027
rect 86358 580957 86418 581571
rect 86355 580956 86421 580957
rect 86355 580892 86356 580956
rect 86420 580892 86421 580956
rect 86355 580891 86421 580892
rect 86726 580005 86786 582387
rect 86907 580412 86973 580413
rect 86907 580348 86908 580412
rect 86972 580348 86973 580412
rect 86907 580347 86973 580348
rect 86723 580004 86789 580005
rect 86723 579940 86724 580004
rect 86788 579940 86789 580004
rect 86723 579939 86789 579940
rect 86910 570890 86970 580347
rect 86726 570830 86970 570890
rect 85990 569910 86270 569970
rect 85990 470610 86050 569910
rect 86726 565538 86786 570830
rect 87278 568850 87338 584291
rect 87459 581364 87525 581365
rect 87459 581300 87460 581364
rect 87524 581300 87525 581364
rect 87459 581299 87525 581300
rect 87094 568790 87338 568850
rect 87094 562050 87154 568790
rect 86726 561990 87154 562050
rect 86726 548450 86786 561990
rect 86726 548390 86970 548450
rect 86910 534850 86970 548390
rect 86726 534790 86970 534850
rect 86726 530178 86786 534790
rect 87094 526010 87154 557822
rect 87462 554570 87522 581299
rect 87646 580410 87706 585651
rect 89667 585036 89733 585037
rect 89667 584972 89668 585036
rect 89732 584972 89733 585036
rect 89667 584971 89733 584972
rect 88195 584900 88261 584901
rect 88195 584836 88196 584900
rect 88260 584836 88261 584900
rect 88195 584835 88261 584836
rect 88011 581772 88077 581773
rect 88011 581708 88012 581772
rect 88076 581708 88077 581772
rect 88011 581707 88077 581708
rect 87646 580350 87890 580410
rect 87643 580004 87709 580005
rect 87643 579940 87644 580004
rect 87708 579940 87709 580004
rect 87643 579939 87709 579940
rect 86726 525950 87154 526010
rect 87278 554510 87522 554570
rect 87278 526010 87338 554510
rect 87278 525950 87522 526010
rect 86726 520658 86786 525950
rect 86874 519830 87154 519890
rect 86726 512410 86786 519062
rect 87094 518802 87154 519830
rect 86910 518742 87154 518802
rect 86910 515130 86970 518742
rect 86910 515070 87338 515130
rect 86726 512350 87154 512410
rect 87094 511050 87154 512350
rect 86910 510990 87154 511050
rect 86910 502298 86970 510990
rect 87278 510370 87338 515070
rect 87094 510310 87338 510370
rect 87094 509010 87154 510310
rect 87094 508950 87338 509010
rect 87278 507650 87338 508950
rect 87462 507650 87522 525950
rect 87094 507590 87522 507650
rect 87094 506970 87154 507590
rect 87278 506970 87338 507590
rect 87094 506910 87522 506970
rect 87278 499490 87338 506910
rect 87094 499430 87338 499490
rect 86726 492778 86786 496622
rect 87094 490650 87154 499430
rect 87462 498810 87522 506910
rect 87278 498750 87522 498810
rect 87278 490650 87338 498750
rect 86910 490590 87338 490650
rect 86910 487250 86970 490590
rect 87094 489970 87154 490590
rect 87094 489910 87522 489970
rect 86910 487190 87338 487250
rect 86874 483110 87154 483170
rect 87094 481810 87154 483110
rect 86874 481750 87154 481810
rect 85990 470550 86602 470610
rect 86542 467530 86602 470550
rect 85990 467470 86602 467530
rect 85990 258770 86050 467470
rect 86726 419930 86786 472142
rect 87278 455970 87338 487190
rect 86910 455910 87338 455970
rect 86910 442370 86970 455910
rect 86910 442310 87154 442370
rect 87094 440330 87154 442310
rect 87094 440270 87338 440330
rect 86726 419870 87154 419930
rect 87094 415850 87154 419870
rect 86726 415790 87154 415850
rect 86726 402930 86786 415790
rect 87278 407690 87338 440270
rect 87094 407630 87338 407690
rect 86726 402870 86970 402930
rect 86910 398170 86970 402870
rect 86726 398110 86970 398170
rect 86726 349978 86786 398110
rect 87094 389330 87154 407630
rect 87094 389270 87338 389330
rect 87278 350570 87338 389270
rect 87094 350510 87338 350570
rect 87094 349210 87154 350510
rect 87094 349150 87338 349210
rect 86726 328898 86786 349062
rect 87278 343650 87338 349150
rect 86910 343590 87338 343650
rect 86910 329490 86970 343590
rect 87462 340370 87522 489910
rect 87646 340370 87706 579939
rect 87830 340370 87890 580350
rect 88014 340370 88074 581707
rect 87094 340310 88074 340370
rect 87094 331258 87154 340310
rect 87462 331258 87522 340310
rect 87646 331258 87706 340310
rect 87830 331258 87890 340310
rect 88198 331258 88258 584835
rect 88379 584628 88445 584629
rect 88379 584564 88380 584628
rect 88444 584564 88445 584628
rect 88379 584563 88445 584564
rect 88382 575650 88442 584563
rect 88563 584220 88629 584221
rect 88563 584156 88564 584220
rect 88628 584156 88629 584220
rect 88563 584155 88629 584156
rect 88336 575590 88442 575650
rect 88336 574970 88396 575590
rect 88336 574910 88442 574970
rect 88382 331258 88442 574910
rect 88566 526010 88626 584155
rect 89483 582860 89549 582861
rect 89483 582796 89484 582860
rect 89548 582796 89549 582860
rect 89483 582795 89549 582796
rect 89115 582180 89181 582181
rect 89115 582116 89116 582180
rect 89180 582116 89181 582180
rect 89115 582115 89181 582116
rect 88931 580004 88997 580005
rect 88931 579940 88932 580004
rect 88996 579940 88997 580004
rect 88931 579939 88997 579940
rect 88566 525950 88810 526010
rect 88750 509010 88810 525950
rect 88566 508950 88810 509010
rect 88566 497450 88626 508950
rect 88934 500170 88994 579939
rect 88750 500110 88994 500170
rect 88750 497450 88810 500110
rect 88566 497390 88994 497450
rect 88750 496090 88810 497390
rect 88566 496030 88810 496090
rect 88566 486570 88626 496030
rect 88934 487930 88994 497390
rect 88750 487870 88994 487930
rect 88750 486570 88810 487870
rect 88566 486510 88994 486570
rect 88750 485890 88810 486510
rect 88566 485830 88810 485890
rect 88566 331258 88626 485830
rect 87094 331198 88810 331258
rect 86910 329430 87154 329490
rect 87094 328130 87154 329430
rect 87462 328130 87522 331198
rect 86874 328070 87154 328130
rect 87278 328070 87522 328130
rect 87278 327858 87338 328070
rect 87646 327858 87706 331198
rect 87830 330850 87890 331198
rect 87830 330790 88074 330850
rect 88014 330170 88074 330790
rect 88198 330170 88258 331198
rect 88382 330170 88442 331198
rect 88566 330170 88626 331198
rect 88750 330170 88810 331198
rect 87094 327798 87338 327858
rect 87462 327798 87706 327858
rect 87830 330110 88810 330170
rect 86174 320130 86270 320190
rect 86174 318610 86234 320130
rect 86174 318550 86270 318610
rect 86726 302378 86786 327302
rect 87094 326090 87154 327798
rect 86910 326030 87154 326090
rect 86910 319970 86970 326030
rect 87462 325410 87522 327798
rect 87830 327450 87890 330110
rect 88014 329850 88074 330110
rect 88198 329850 88258 330110
rect 88382 329850 88442 330110
rect 88566 329850 88626 330110
rect 88014 329790 88626 329850
rect 88198 329490 88258 329790
rect 88382 329490 88442 329790
rect 88566 329490 88626 329790
rect 87426 325350 87522 325410
rect 87646 327390 87890 327450
rect 88014 329430 88626 329490
rect 86910 319910 87154 319970
rect 87094 317250 87154 319910
rect 87278 317430 87338 324582
rect 87646 324138 87706 327390
rect 88014 323370 88074 329430
rect 88198 325410 88258 329430
rect 88382 326770 88442 329430
rect 88566 326770 88626 329430
rect 88934 328810 88994 486510
rect 88750 328750 88994 328810
rect 88750 327450 88810 328750
rect 88750 327390 88994 327450
rect 88382 326710 88626 326770
rect 88566 326090 88626 326710
rect 88566 326030 88810 326090
rect 88566 325710 88626 326030
rect 88382 325650 88626 325710
rect 88382 325410 88442 325650
rect 88198 325350 88626 325410
rect 87462 323310 88074 323370
rect 87462 320190 87522 323310
rect 87462 320130 87706 320190
rect 87646 318810 87706 320130
rect 88014 318810 88074 322542
rect 88382 320650 88442 325350
rect 88290 320590 88442 320650
rect 88290 320190 88350 320590
rect 88198 320130 88350 320190
rect 88198 318810 88258 320130
rect 87646 318750 88442 318810
rect 88014 318610 88074 318750
rect 87830 318550 88074 318610
rect 87278 317370 87522 317430
rect 87094 317190 87338 317250
rect 87278 316050 87338 317190
rect 87462 316050 87522 317370
rect 87242 315990 87706 316050
rect 87278 300250 87338 315990
rect 87058 300190 87338 300250
rect 87462 299570 87522 315990
rect 86726 299510 87522 299570
rect 86726 296730 86786 299510
rect 87646 298890 87706 315990
rect 86358 296670 86786 296730
rect 87094 298830 87706 298890
rect 86358 294810 86418 296670
rect 86358 294750 86602 294810
rect 86542 290050 86602 294750
rect 86726 290050 86786 296022
rect 87094 292590 87154 298830
rect 86910 292530 87154 292590
rect 86910 290050 86970 292530
rect 87462 290050 87522 298062
rect 86542 289990 87154 290050
rect 86726 288450 86786 289990
rect 86910 288690 86970 289990
rect 87094 289370 87154 289990
rect 87278 289990 87522 290050
rect 87278 289370 87338 289990
rect 87094 289310 87522 289370
rect 86910 288630 87154 288690
rect 87094 288450 87154 288630
rect 86506 288390 87154 288450
rect 86358 278578 86418 279702
rect 85990 258710 86234 258770
rect 86174 256730 86234 258710
rect 85990 256670 86234 256730
rect 85990 209790 86050 256670
rect 86726 255330 86786 288390
rect 87278 288010 87338 289310
rect 86910 287950 87338 288010
rect 86910 283250 86970 287950
rect 87462 287070 87522 289310
rect 87830 287330 87890 318550
rect 88198 317250 88258 318750
rect 88014 317190 88258 317250
rect 88382 317930 88442 318750
rect 88566 317930 88626 325350
rect 88382 317870 88626 317930
rect 88014 316050 88074 317190
rect 88382 316570 88442 317870
rect 88566 316570 88626 317870
rect 88750 316570 88810 326030
rect 88198 316510 88810 316570
rect 88198 316050 88258 316510
rect 88382 316050 88442 316510
rect 88014 315990 88442 316050
rect 88014 293450 88074 315990
rect 88198 293450 88258 315990
rect 88382 311810 88442 315990
rect 88566 311810 88626 316510
rect 88382 311750 88810 311810
rect 88566 300930 88626 311750
rect 88750 300930 88810 311750
rect 88382 300870 88810 300930
rect 88382 300250 88442 300870
rect 88566 300250 88626 300870
rect 88382 300190 88626 300250
rect 88382 293970 88442 300190
rect 88566 293970 88626 300190
rect 88382 293910 88810 293970
rect 88566 293450 88626 293910
rect 88750 293450 88810 293910
rect 88014 293390 88810 293450
rect 88198 288450 88258 293390
rect 88566 292770 88626 293390
rect 88750 292770 88810 293390
rect 87278 287010 87522 287070
rect 87646 287270 87890 287330
rect 88014 288390 88258 288450
rect 88382 292710 88810 292770
rect 87646 287070 87706 287270
rect 88014 287070 88074 288390
rect 87646 287010 88258 287070
rect 87278 283250 87338 287010
rect 86910 283190 87522 283250
rect 87278 281890 87338 283190
rect 86910 281830 87338 281890
rect 86910 276030 86970 281830
rect 87462 281210 87522 283190
rect 87278 281150 87522 281210
rect 86910 275970 87154 276030
rect 87094 274650 87154 275970
rect 87278 274650 87338 281150
rect 87646 277810 87706 286502
rect 88014 285290 88074 287010
rect 88198 285290 88258 287010
rect 87462 277750 87706 277810
rect 87830 285230 88258 285290
rect 87462 274650 87522 277750
rect 87094 274590 87706 274650
rect 86726 255270 86970 255330
rect 86910 247050 86970 255270
rect 87278 247050 87338 274590
rect 87462 247050 87522 274590
rect 87646 247050 87706 274590
rect 87830 247050 87890 285230
rect 88014 277410 88074 285230
rect 88382 277410 88442 292710
rect 88566 277410 88626 292710
rect 88750 277410 88810 292710
rect 88014 277350 88810 277410
rect 88014 247050 88074 277350
rect 88198 262170 88258 277350
rect 88382 262170 88442 277350
rect 88566 262170 88626 277350
rect 88198 262110 88810 262170
rect 88382 258090 88442 262110
rect 86726 246990 88074 247050
rect 88198 258030 88442 258090
rect 88198 255330 88258 258030
rect 88566 255330 88626 262110
rect 88198 255270 88626 255330
rect 88198 251290 88258 255270
rect 88382 254690 88442 255270
rect 88750 254690 88810 262110
rect 88382 254630 88810 254690
rect 88750 252650 88810 254630
rect 88382 252590 88810 252650
rect 88382 251290 88442 252590
rect 88198 251230 88442 251290
rect 86726 243810 86786 246990
rect 86910 243810 86970 246990
rect 87278 246530 87338 246990
rect 87462 246530 87522 246990
rect 87278 246470 87522 246530
rect 87278 245170 87338 246470
rect 87462 245170 87522 246470
rect 87830 245170 87890 246990
rect 88198 246530 88258 251230
rect 88290 251190 88350 251230
rect 88290 251130 88442 251190
rect 88382 247890 88442 251130
rect 88750 248029 88810 252590
rect 88747 248028 88813 248029
rect 88747 247964 88748 248028
rect 88812 247964 88813 248028
rect 88747 247963 88813 247964
rect 88382 247830 88810 247890
rect 88379 247756 88445 247757
rect 88379 247692 88380 247756
rect 88444 247692 88445 247756
rect 88379 247691 88445 247692
rect 88382 246530 88442 247691
rect 88198 246470 88442 246530
rect 87278 245110 87706 245170
rect 87830 245110 88074 245170
rect 87278 244490 87338 245110
rect 87462 244490 87522 245110
rect 87646 244490 87706 245110
rect 87278 244430 87890 244490
rect 87278 243810 87338 244430
rect 86726 243750 87522 243810
rect 86910 242910 86970 243750
rect 86726 242850 86970 242910
rect 86358 232658 86418 232782
rect 86174 232598 86418 232658
rect 86174 230890 86234 232598
rect 86726 232250 86786 242850
rect 87278 241770 87338 243750
rect 87242 241710 87338 241770
rect 87462 239594 87522 243750
rect 87278 239534 87522 239594
rect 87278 238370 87338 239534
rect 87646 239138 87706 244430
rect 87830 238770 87890 244430
rect 87646 238710 87890 238770
rect 87646 238458 87706 238710
rect 86690 232190 86786 232250
rect 86910 238310 87338 238370
rect 86910 231570 86970 238310
rect 88014 237690 88074 245110
rect 88198 243810 88258 246470
rect 88198 243750 88442 243810
rect 88198 243130 88258 243750
rect 88382 243130 88442 243750
rect 88750 243130 88810 247830
rect 88198 243070 88810 243130
rect 87278 237630 88074 237690
rect 87278 234378 87338 237630
rect 88382 237010 88442 243070
rect 88750 242910 88810 243070
rect 88566 242850 88810 242910
rect 88566 238370 88626 242850
rect 88750 238370 88810 242850
rect 88934 238370 88994 327390
rect 89118 238370 89178 582115
rect 89299 581364 89365 581365
rect 89299 581300 89300 581364
rect 89364 581300 89365 581364
rect 89299 581299 89365 581300
rect 89302 238370 89362 581299
rect 88566 238310 89362 238370
rect 88566 237010 88626 238310
rect 88750 237010 88810 238310
rect 88014 236950 88810 237010
rect 87646 234834 87706 236862
rect 88014 234834 88074 236950
rect 87462 234774 88074 234834
rect 88382 236330 88442 236950
rect 88566 236330 88626 236950
rect 88382 236270 88810 236330
rect 87462 233018 87522 234774
rect 87646 233250 87706 234774
rect 88382 233610 88442 236270
rect 88566 233610 88626 236270
rect 88014 233550 88626 233610
rect 87646 233190 87890 233250
rect 87830 232930 87890 233190
rect 87610 232870 87890 232930
rect 87827 232796 87893 232797
rect 87462 232658 87522 232782
rect 87827 232732 87828 232796
rect 87892 232732 87893 232796
rect 87827 232731 87893 232732
rect 87462 232598 87706 232658
rect 87646 232250 87706 232598
rect 87830 232250 87890 232731
rect 86874 231510 86970 231570
rect 87462 232190 87890 232250
rect 86174 230830 86970 230890
rect 86910 230210 86970 230830
rect 87462 230754 87522 232190
rect 87646 231870 87706 232190
rect 87646 231810 87890 231870
rect 87830 230754 87890 231810
rect 88014 230890 88074 233550
rect 88382 231658 88442 233550
rect 88750 233069 88810 236270
rect 88747 233068 88813 233069
rect 88747 233004 88748 233068
rect 88812 233004 88813 233068
rect 88747 233003 88813 233004
rect 88014 230830 88810 230890
rect 87462 230694 88442 230754
rect 87830 230210 87890 230694
rect 88382 230490 88442 230694
rect 88382 230430 88626 230490
rect 86690 230150 86786 230210
rect 86910 230150 87338 230210
rect 87830 230150 88074 230210
rect 86726 229530 86786 230150
rect 87278 229530 87338 230150
rect 88014 229530 88074 230150
rect 86506 229470 86970 229530
rect 87278 229470 87890 229530
rect 88014 229470 88258 229530
rect 86726 228850 86786 229470
rect 86910 228850 86970 229470
rect 86726 228790 87522 228850
rect 86910 228170 86970 228790
rect 87462 228170 87522 228790
rect 87830 228170 87890 229470
rect 86910 228110 88074 228170
rect 86506 227430 87338 227490
rect 86171 226812 86237 226813
rect 86171 226748 86172 226812
rect 86236 226810 86237 226812
rect 86236 226750 86786 226810
rect 86236 226748 86237 226750
rect 86171 226747 86237 226748
rect 86726 224090 86786 226750
rect 86726 224030 87154 224090
rect 87094 223410 87154 224030
rect 87278 223410 87338 227430
rect 87462 226538 87522 228110
rect 87830 226538 87890 228110
rect 88014 226538 88074 228110
rect 88198 226538 88258 229470
rect 88566 226538 88626 230430
rect 87462 226478 88626 226538
rect 88750 226538 88810 230830
rect 88934 226538 88994 238310
rect 89118 226538 89178 238310
rect 88750 226478 89362 226538
rect 86874 223350 87706 223410
rect 86874 222670 86970 222730
rect 86910 222050 86970 222670
rect 87094 222050 87154 223350
rect 87278 222050 87338 223350
rect 87646 222050 87706 223350
rect 86726 221990 87706 222050
rect 86726 220690 86786 221990
rect 86910 220690 86970 221990
rect 87094 220690 87154 221990
rect 86174 220630 87154 220690
rect 86174 218070 86234 220630
rect 86174 218010 86602 218070
rect 86542 217290 86602 218010
rect 86726 217290 86786 220630
rect 86910 218650 86970 220630
rect 87278 220010 87338 221990
rect 87830 221370 87890 226478
rect 88014 226350 88074 226478
rect 88198 226350 88258 226478
rect 88566 226350 88626 226478
rect 88014 226290 88442 226350
rect 88198 226130 88258 226290
rect 88382 226130 88442 226290
rect 87646 221310 87890 221370
rect 88014 226070 88442 226130
rect 88566 226290 88810 226350
rect 87646 220690 87706 221310
rect 88014 220690 88074 226070
rect 88198 220690 88258 226070
rect 88566 225450 88626 226290
rect 87094 219950 87338 220010
rect 87462 220630 87706 220690
rect 87830 220630 88258 220690
rect 88382 225390 88626 225450
rect 87094 218786 87154 219950
rect 87462 219418 87522 220630
rect 87830 218786 87890 220630
rect 88014 220010 88074 220630
rect 88014 219950 88258 220010
rect 88198 218786 88258 219950
rect 88382 219330 88442 225390
rect 88750 222210 88810 226290
rect 87094 218726 87338 218786
rect 86910 218590 87154 218650
rect 86174 217230 86786 217290
rect 86174 216610 86234 217230
rect 86174 216550 86418 216610
rect 86358 214658 86418 216550
rect 86726 211850 86786 217230
rect 87094 213210 87154 218590
rect 87278 213930 87338 218726
rect 87462 218726 87890 218786
rect 88014 218726 88258 218786
rect 88336 219270 88442 219330
rect 88566 222150 88810 222210
rect 88566 220690 88626 222150
rect 88934 221370 88994 226478
rect 88750 221310 88994 221370
rect 88750 220690 88810 221310
rect 88566 220630 88994 220690
rect 87462 218514 87522 218726
rect 88014 218514 88074 218726
rect 88336 218650 88396 219270
rect 87462 218454 87706 218514
rect 87646 218070 87706 218454
rect 87462 218010 87706 218070
rect 87830 218454 88074 218514
rect 88244 218590 88396 218650
rect 88566 218650 88626 220630
rect 88566 218590 88810 218650
rect 87462 215250 87522 218010
rect 87830 216018 87890 218454
rect 88244 218070 88304 218590
rect 88244 218010 88442 218070
rect 87462 215190 87706 215250
rect 87646 214658 87706 215190
rect 88382 214658 88442 218010
rect 87278 213870 88626 213930
rect 87094 213150 87522 213210
rect 87462 212530 87522 213150
rect 87462 212470 87890 212530
rect 86726 211790 87338 211850
rect 86726 211110 87154 211170
rect 86726 210578 86786 211110
rect 85990 209730 86786 209790
rect 85806 209070 86050 209130
rect 85990 208538 86050 209070
rect 84518 202950 84762 203010
rect 84886 208390 85682 208450
rect 84518 198250 84578 202950
rect 84886 202418 84946 208390
rect 85254 202058 85314 205582
rect 84886 201998 85314 202058
rect 84886 199018 84946 201998
rect 85622 201650 85682 204902
rect 85990 202418 86050 206262
rect 86726 205818 86786 209730
rect 86174 205670 86270 205730
rect 86174 203690 86234 205670
rect 87094 205730 87154 211110
rect 87278 208410 87338 211790
rect 87278 208350 87522 208410
rect 87462 207030 87522 208350
rect 87278 206970 87522 207030
rect 87278 206274 87338 206970
rect 87278 206214 87374 206274
rect 87094 205670 87338 205730
rect 86174 203630 86786 203690
rect 85622 201590 85902 201650
rect 84518 198190 85130 198250
rect 84150 196830 84762 196890
rect 84702 196298 84762 196830
rect 83966 196150 84394 196210
rect 82491 195195 82557 195196
rect 82632 195198 83290 195258
rect 83414 195198 83842 195258
rect 82494 192405 82554 195195
rect 82632 194989 82692 195198
rect 82629 194988 82695 194989
rect 82629 194924 82630 194988
rect 82694 194924 82695 194988
rect 82629 194923 82695 194924
rect 82629 194852 82695 194853
rect 82629 194788 82630 194852
rect 82694 194850 82695 194852
rect 82694 194790 82774 194850
rect 82694 194788 82695 194790
rect 82629 194787 82695 194788
rect 83414 194850 83474 195198
rect 84334 194938 84394 196150
rect 85070 195258 85130 198190
rect 85254 196890 85314 201502
rect 85990 198250 86050 198782
rect 85806 198190 86050 198250
rect 85254 196830 85682 196890
rect 84702 195198 85130 195258
rect 83230 194790 83474 194850
rect 82491 192404 82557 192405
rect 82491 192340 82492 192404
rect 82556 192340 82557 192404
rect 82491 192339 82557 192340
rect 82629 192404 82695 192405
rect 82629 192340 82630 192404
rect 82694 192402 82695 192404
rect 82862 192402 82922 194022
rect 82694 192342 82922 192402
rect 82694 192340 82695 192342
rect 82629 192339 82695 192340
rect 82310 192206 82738 192266
rect 82491 191996 82557 191997
rect 82491 191932 82492 191996
rect 82556 191932 82557 191996
rect 82491 191931 82557 191932
rect 82494 191181 82554 191931
rect 82678 191453 82738 192206
rect 82629 191452 82738 191453
rect 82629 191388 82630 191452
rect 82694 191390 82738 191452
rect 83230 191450 83290 194790
rect 83598 191538 83658 194022
rect 83046 191390 83290 191450
rect 82694 191388 82695 191390
rect 82629 191387 82695 191388
rect 82491 191180 82557 191181
rect 82491 191116 82492 191180
rect 82556 191116 82557 191180
rect 82491 191115 82557 191116
rect 82491 190908 82557 190909
rect 82491 190858 82492 190908
rect 82556 190858 82557 190908
rect 82307 190500 82373 190501
rect 82307 190436 82308 190500
rect 82372 190436 82373 190500
rect 82307 190435 82373 190436
rect 82310 181250 82370 190435
rect 82629 190364 82695 190365
rect 82629 190300 82630 190364
rect 82694 190362 82695 190364
rect 83046 190362 83106 191390
rect 83966 191178 84026 191982
rect 82694 190302 83106 190362
rect 83782 191118 84026 191178
rect 82694 190300 82695 190302
rect 82629 190299 82695 190300
rect 82491 188732 82557 188733
rect 82491 188668 82492 188732
rect 82556 188730 82557 188732
rect 82556 188670 82738 188730
rect 82556 188668 82557 188670
rect 82491 188667 82557 188668
rect 82678 188138 82738 188670
rect 83782 187458 83842 191118
rect 82491 187372 82557 187373
rect 82491 187308 82492 187372
rect 82556 187370 82557 187372
rect 82556 187310 83290 187370
rect 82556 187308 82557 187310
rect 82491 187307 82557 187308
rect 82629 187100 82695 187101
rect 82629 187036 82630 187100
rect 82694 187036 82695 187100
rect 82629 187035 82695 187036
rect 82491 186964 82557 186965
rect 82491 186900 82492 186964
rect 82556 186900 82557 186964
rect 82632 186962 82692 187035
rect 82632 186902 83106 186962
rect 82491 186899 82557 186900
rect 82494 181389 82554 186899
rect 82491 181388 82557 181389
rect 82491 181324 82492 181388
rect 82556 181324 82557 181388
rect 82491 181323 82557 181324
rect 82310 181190 82738 181250
rect 82307 181116 82373 181117
rect 82307 181052 82308 181116
rect 82372 181052 82373 181116
rect 82307 181051 82373 181052
rect 82310 174589 82370 181051
rect 82491 179892 82557 179893
rect 82491 179828 82492 179892
rect 82556 179890 82557 179892
rect 82678 179890 82738 181190
rect 82556 179830 82738 179890
rect 82556 179828 82557 179830
rect 82491 179827 82557 179828
rect 83046 179210 83106 186902
rect 83230 186690 83290 187310
rect 83230 186630 83878 186690
rect 84334 183970 84394 191302
rect 84702 191178 84762 195198
rect 84702 191118 85498 191178
rect 84886 190498 84946 190622
rect 84518 190438 84946 190498
rect 84518 186962 84578 190438
rect 84886 187370 84946 187902
rect 84886 187310 85314 187370
rect 84518 186902 85130 186962
rect 84702 185330 84762 186542
rect 84702 185270 84946 185330
rect 84150 183910 84394 183970
rect 83414 179978 83474 183142
rect 84150 179978 84210 183910
rect 84518 181386 84578 183142
rect 84518 181326 84762 181386
rect 83046 179150 83842 179210
rect 82491 178668 82557 178669
rect 82491 178604 82492 178668
rect 82556 178604 82557 178668
rect 82678 178666 82738 179062
rect 82678 178606 83106 178666
rect 82491 178603 82557 178604
rect 82494 178530 82554 178603
rect 82494 178470 82738 178530
rect 82491 178396 82557 178397
rect 82491 178332 82492 178396
rect 82556 178332 82557 178396
rect 82491 178331 82557 178332
rect 82307 174588 82373 174589
rect 82307 174524 82308 174588
rect 82372 174524 82373 174588
rect 82307 174523 82373 174524
rect 82494 174450 82554 178331
rect 82678 175133 82738 178470
rect 82629 175132 82738 175133
rect 82629 175068 82630 175132
rect 82694 175070 82738 175132
rect 83046 175130 83106 178606
rect 83782 178530 83842 179150
rect 84334 178666 84394 179062
rect 84334 178606 84578 178666
rect 83782 178470 84394 178530
rect 83414 177850 83474 178382
rect 83414 177790 84026 177850
rect 83598 176490 83658 177022
rect 83598 176430 83842 176490
rect 83046 175070 83474 175130
rect 82694 175068 82695 175070
rect 82629 175067 82695 175068
rect 82310 174390 82554 174450
rect 82123 170644 82189 170645
rect 82123 170580 82124 170644
rect 82188 170580 82189 170644
rect 82123 170579 82189 170580
rect 82123 169828 82189 169829
rect 82123 169764 82124 169828
rect 82188 169764 82189 169828
rect 82123 169763 82189 169764
rect 82126 11797 82186 169763
rect 82310 159085 82370 174390
rect 82491 173908 82557 173909
rect 82491 173844 82492 173908
rect 82556 173844 82557 173908
rect 82491 173843 82557 173844
rect 82678 173846 82922 173906
rect 82494 171869 82554 173843
rect 82678 173773 82738 173846
rect 82629 173772 82738 173773
rect 82629 173708 82630 173772
rect 82694 173710 82738 173772
rect 82694 173708 82695 173710
rect 82629 173707 82695 173708
rect 82629 172412 82695 172413
rect 82629 172348 82630 172412
rect 82694 172410 82695 172412
rect 82862 172410 82922 173846
rect 83414 172498 83474 175070
rect 82694 172350 82922 172410
rect 82694 172348 82695 172350
rect 82629 172347 82695 172348
rect 82491 171868 82557 171869
rect 82491 171804 82492 171868
rect 82556 171804 82557 171868
rect 83782 171866 83842 176430
rect 82491 171803 82557 171804
rect 83046 171806 83842 171866
rect 83046 171730 83106 171806
rect 82862 171670 83106 171730
rect 82491 171596 82557 171597
rect 82491 171532 82492 171596
rect 82556 171532 82557 171596
rect 82862 171594 82922 171670
rect 82491 171531 82557 171532
rect 82632 171534 82922 171594
rect 82494 170642 82554 171531
rect 82632 171461 82692 171534
rect 82629 171460 82695 171461
rect 82629 171396 82630 171460
rect 82694 171396 82695 171460
rect 82629 171395 82695 171396
rect 82629 171052 82695 171053
rect 82629 170988 82630 171052
rect 82694 171050 82695 171052
rect 82694 170990 83290 171050
rect 82694 170988 82695 170990
rect 82629 170987 82695 170988
rect 82494 170582 83106 170642
rect 82491 170508 82557 170509
rect 82491 170444 82492 170508
rect 82556 170444 82557 170508
rect 82491 170443 82557 170444
rect 82629 170508 82695 170509
rect 82629 170444 82630 170508
rect 82694 170506 82695 170508
rect 82694 170446 82922 170506
rect 82694 170444 82695 170446
rect 82629 170443 82695 170444
rect 82494 170370 82554 170443
rect 82494 170310 82738 170370
rect 82491 170100 82557 170101
rect 82491 170036 82492 170100
rect 82556 170036 82557 170100
rect 82491 170035 82557 170036
rect 82494 162213 82554 170035
rect 82491 162212 82557 162213
rect 82491 162148 82492 162212
rect 82556 162148 82557 162212
rect 82491 162147 82557 162148
rect 82491 160852 82557 160853
rect 82491 160788 82492 160852
rect 82556 160850 82557 160852
rect 82678 160850 82738 170310
rect 82556 160790 82738 160850
rect 82556 160788 82557 160790
rect 82491 160787 82557 160788
rect 82307 159084 82373 159085
rect 82307 159020 82308 159084
rect 82372 159020 82373 159084
rect 82307 159019 82373 159020
rect 82862 158946 82922 170446
rect 82310 158886 82922 158946
rect 82310 156773 82370 158886
rect 83046 158810 83106 170582
rect 82494 158750 83106 158810
rect 82494 157450 82554 158750
rect 83230 158538 83290 170990
rect 83966 170458 84026 177790
rect 84334 170098 84394 178470
rect 84150 170038 84394 170098
rect 84150 169778 84210 170038
rect 83046 158478 83290 158538
rect 83414 168814 84026 168874
rect 83046 157450 83106 158478
rect 82494 157390 82922 157450
rect 83046 157390 83290 157450
rect 82491 157316 82557 157317
rect 82491 157252 82492 157316
rect 82556 157252 82557 157316
rect 82862 157314 82922 157390
rect 82862 157254 83106 157314
rect 82491 157251 82557 157252
rect 82307 156772 82373 156773
rect 82307 156708 82308 156772
rect 82372 156708 82373 156772
rect 82307 156707 82373 156708
rect 82494 149701 82554 157251
rect 82629 156772 82695 156773
rect 82629 156708 82630 156772
rect 82694 156770 82695 156772
rect 82694 156710 82922 156770
rect 82694 156708 82695 156710
rect 82629 156707 82695 156708
rect 82491 149700 82557 149701
rect 82491 149636 82492 149700
rect 82556 149636 82557 149700
rect 82491 149635 82557 149636
rect 82307 146844 82373 146845
rect 82307 146780 82308 146844
rect 82372 146780 82373 146844
rect 82307 146779 82373 146780
rect 82310 144533 82370 146779
rect 82307 144532 82373 144533
rect 82307 144468 82308 144532
rect 82372 144468 82373 144532
rect 82862 144530 82922 156710
rect 82307 144467 82373 144468
rect 82494 144470 82922 144530
rect 82494 143850 82554 144470
rect 82310 143790 82554 143850
rect 82310 138410 82370 143790
rect 82491 143172 82557 143173
rect 82491 143108 82492 143172
rect 82556 143108 82557 143172
rect 82491 143107 82557 143108
rect 82494 141949 82554 143107
rect 82491 141948 82557 141949
rect 82491 141884 82492 141948
rect 82556 141884 82557 141948
rect 82491 141883 82557 141884
rect 82310 138350 82922 138410
rect 82491 137460 82557 137461
rect 82491 137396 82492 137460
rect 82556 137396 82557 137460
rect 82491 137395 82557 137396
rect 82307 137324 82373 137325
rect 82307 137260 82308 137324
rect 82372 137260 82373 137324
rect 82307 137259 82373 137260
rect 82310 136101 82370 137259
rect 82494 136370 82554 137395
rect 82494 136310 82738 136370
rect 82307 136100 82373 136101
rect 82307 136036 82308 136100
rect 82372 136036 82373 136100
rect 82307 136035 82373 136036
rect 82491 136100 82557 136101
rect 82491 136036 82492 136100
rect 82556 136036 82557 136100
rect 82491 136035 82557 136036
rect 82307 135964 82373 135965
rect 82307 135900 82308 135964
rect 82372 135900 82373 135964
rect 82307 135899 82373 135900
rect 82310 116517 82370 135899
rect 82494 129029 82554 136035
rect 82491 129028 82557 129029
rect 82491 128964 82492 129028
rect 82556 128964 82557 129028
rect 82491 128963 82557 128964
rect 82678 123589 82738 136310
rect 82675 123588 82741 123589
rect 82675 123524 82676 123588
rect 82740 123524 82741 123588
rect 82675 123523 82741 123524
rect 82862 120733 82922 138350
rect 82859 120732 82925 120733
rect 82859 120668 82860 120732
rect 82924 120668 82925 120732
rect 82859 120667 82925 120668
rect 82307 116516 82373 116517
rect 82307 116452 82308 116516
rect 82372 116452 82373 116516
rect 82307 116451 82373 116452
rect 82859 106996 82925 106997
rect 82859 106932 82860 106996
rect 82924 106932 82925 106996
rect 82859 106931 82925 106932
rect 82862 98021 82922 106931
rect 82859 98020 82925 98021
rect 82859 97956 82860 98020
rect 82924 97956 82925 98020
rect 82859 97955 82925 97956
rect 82859 84964 82925 84965
rect 82859 84900 82860 84964
rect 82924 84900 82925 84964
rect 82859 84899 82925 84900
rect 82862 78709 82922 84899
rect 82859 78708 82925 78709
rect 82859 78644 82860 78708
rect 82924 78644 82925 78708
rect 82859 78643 82925 78644
rect 82859 65516 82925 65517
rect 82859 65452 82860 65516
rect 82924 65452 82925 65516
rect 82859 65451 82925 65452
rect 82862 55861 82922 65451
rect 82859 55860 82925 55861
rect 82859 55796 82860 55860
rect 82924 55796 82925 55860
rect 82859 55795 82925 55796
rect 83046 13021 83106 157254
rect 83230 118013 83290 157390
rect 83414 153370 83474 168814
rect 83966 168738 84026 168814
rect 84518 168738 84578 178606
rect 83966 168678 84578 168738
rect 83966 164930 84026 165462
rect 83966 164870 84210 164930
rect 83782 158898 83842 162742
rect 84150 161530 84210 164870
rect 83966 161470 84210 161530
rect 83966 160170 84026 161470
rect 84334 160938 84394 166822
rect 83966 160110 84210 160170
rect 84150 158810 84210 160110
rect 84150 158750 84578 158810
rect 83966 157314 84026 157982
rect 83966 157254 84394 157314
rect 83782 154050 83842 155262
rect 83782 153990 84210 154050
rect 83414 153310 84026 153370
rect 83598 150738 83658 151862
rect 83966 149698 84026 153310
rect 83414 149638 84026 149698
rect 83414 140858 83474 149638
rect 84150 149290 84210 153990
rect 83966 149230 84210 149290
rect 83966 145890 84026 149230
rect 84334 147250 84394 157254
rect 83782 145830 84026 145890
rect 84150 147190 84394 147250
rect 83782 141898 83842 145830
rect 84150 144618 84210 147190
rect 84518 141130 84578 158750
rect 84114 141070 84578 141130
rect 83414 140798 84026 140858
rect 83598 130338 83658 140302
rect 83966 131018 84026 140798
rect 84334 133058 84394 140302
rect 84702 130930 84762 181326
rect 84518 130870 84762 130930
rect 83414 129510 84062 129570
rect 83414 127530 83474 129510
rect 83368 127470 83474 127530
rect 83368 126170 83428 127470
rect 83368 126110 83474 126170
rect 83227 118012 83293 118013
rect 83227 117948 83228 118012
rect 83292 117948 83293 118012
rect 83227 117947 83293 117948
rect 83414 106997 83474 126110
rect 83779 123996 83845 123997
rect 83779 123932 83780 123996
rect 83844 123932 83845 123996
rect 83779 123931 83845 123932
rect 84331 123996 84397 123997
rect 84331 123932 84332 123996
rect 84396 123932 84397 123996
rect 84331 123931 84397 123932
rect 83782 122229 83842 123931
rect 83779 122228 83845 122229
rect 83779 122164 83780 122228
rect 83844 122164 83845 122228
rect 83779 122163 83845 122164
rect 83604 121254 84204 122000
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83411 106996 83477 106997
rect 83411 106932 83412 106996
rect 83476 106932 83477 106996
rect 83411 106931 83477 106932
rect 83227 106316 83293 106317
rect 83227 106252 83228 106316
rect 83292 106252 83293 106316
rect 83227 106251 83293 106252
rect 83230 104821 83290 106251
rect 83227 104820 83293 104821
rect 83227 104756 83228 104820
rect 83292 104756 83293 104820
rect 83227 104755 83293 104756
rect 83411 98020 83477 98021
rect 83411 97956 83412 98020
rect 83476 97956 83477 98020
rect 83411 97955 83477 97956
rect 83227 95300 83293 95301
rect 83227 95236 83228 95300
rect 83292 95236 83293 95300
rect 83227 95235 83293 95236
rect 83230 86869 83290 95235
rect 83227 86868 83293 86869
rect 83227 86804 83228 86868
rect 83292 86804 83293 86868
rect 83227 86803 83293 86804
rect 83414 84965 83474 97955
rect 83604 85254 84204 120698
rect 84334 106997 84394 123931
rect 84518 122093 84578 130870
rect 84699 123180 84765 123181
rect 84699 123116 84700 123180
rect 84764 123116 84765 123180
rect 84699 123115 84765 123116
rect 84515 122092 84581 122093
rect 84515 122028 84516 122092
rect 84580 122028 84581 122092
rect 84515 122027 84581 122028
rect 84331 106996 84397 106997
rect 84331 106932 84332 106996
rect 84396 106932 84397 106996
rect 84331 106931 84397 106932
rect 84331 98700 84397 98701
rect 84331 98636 84332 98700
rect 84396 98636 84397 98700
rect 84331 98635 84397 98636
rect 84334 86325 84394 98635
rect 84331 86324 84397 86325
rect 84331 86260 84332 86324
rect 84396 86260 84397 86324
rect 84331 86259 84397 86260
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83411 84964 83477 84965
rect 83411 84900 83412 84964
rect 83476 84900 83477 84964
rect 83411 84899 83477 84900
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83411 78708 83477 78709
rect 83411 78644 83412 78708
rect 83476 78644 83477 78708
rect 83411 78643 83477 78644
rect 83227 77348 83293 77349
rect 83227 77284 83228 77348
rect 83292 77284 83293 77348
rect 83227 77283 83293 77284
rect 83230 77210 83290 77283
rect 83230 77150 83336 77210
rect 83276 77077 83336 77150
rect 83273 77076 83339 77077
rect 83273 77012 83274 77076
rect 83338 77012 83339 77076
rect 83273 77011 83339 77012
rect 83227 67692 83293 67693
rect 83227 67628 83228 67692
rect 83292 67628 83293 67692
rect 83227 67627 83293 67628
rect 83230 57901 83290 67627
rect 83414 65517 83474 78643
rect 83411 65516 83477 65517
rect 83411 65452 83412 65516
rect 83476 65452 83477 65516
rect 83411 65451 83477 65452
rect 83227 57900 83293 57901
rect 83227 57836 83228 57900
rect 83292 57836 83293 57900
rect 83227 57835 83293 57836
rect 83411 55860 83477 55861
rect 83411 55796 83412 55860
rect 83476 55796 83477 55860
rect 83411 55795 83477 55796
rect 83227 48380 83293 48381
rect 83227 48316 83228 48380
rect 83292 48316 83293 48380
rect 83227 48315 83293 48316
rect 83230 38589 83290 48315
rect 83227 38588 83293 38589
rect 83227 38524 83228 38588
rect 83292 38524 83293 38588
rect 83227 38523 83293 38524
rect 83414 35189 83474 55795
rect 83604 49254 84204 84698
rect 84331 78028 84397 78029
rect 84331 77964 84332 78028
rect 84396 77964 84397 78028
rect 84331 77963 84397 77964
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83411 35188 83477 35189
rect 83411 35124 83412 35188
rect 83476 35124 83477 35188
rect 83411 35123 83477 35124
rect 83227 29068 83293 29069
rect 83227 29004 83228 29068
rect 83292 29004 83293 29068
rect 83227 29003 83293 29004
rect 83230 19277 83290 29003
rect 83227 19276 83293 19277
rect 83227 19212 83228 19276
rect 83292 19212 83293 19276
rect 83227 19211 83293 19212
rect 83604 13254 84204 48698
rect 84334 39949 84394 77963
rect 84331 39948 84397 39949
rect 84331 39884 84332 39948
rect 84396 39884 84397 39948
rect 84331 39883 84397 39884
rect 84515 39948 84581 39949
rect 84515 39884 84516 39948
rect 84580 39884 84581 39948
rect 84515 39883 84581 39884
rect 84518 23493 84578 39883
rect 84331 23492 84397 23493
rect 84331 23428 84332 23492
rect 84396 23428 84397 23492
rect 84331 23427 84397 23428
rect 84515 23492 84581 23493
rect 84515 23428 84516 23492
rect 84580 23428 84581 23492
rect 84515 23427 84581 23428
rect 84334 23357 84394 23427
rect 84331 23356 84397 23357
rect 84331 23292 84332 23356
rect 84396 23292 84397 23356
rect 84331 23291 84397 23292
rect 84331 13836 84397 13837
rect 84331 13772 84332 13836
rect 84396 13772 84397 13836
rect 84331 13771 84397 13772
rect 84334 13701 84394 13771
rect 84331 13700 84397 13701
rect 84331 13636 84332 13700
rect 84396 13636 84397 13700
rect 84331 13635 84397 13636
rect 83043 13020 83109 13021
rect 83043 12956 83044 13020
rect 83108 12956 83109 13020
rect 83043 12955 83109 12956
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 82123 11796 82189 11797
rect 82123 11732 82124 11796
rect 82188 11732 82189 11796
rect 82123 11731 82189 11732
rect 81939 6220 82005 6221
rect 81939 6156 81940 6220
rect 82004 6156 82005 6220
rect 81939 6155 82005 6156
rect 80835 3364 80901 3365
rect 80835 3300 80836 3364
rect 80900 3300 80901 3364
rect 80835 3299 80901 3300
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 84331 4180 84397 4181
rect 84331 4116 84332 4180
rect 84396 4116 84397 4180
rect 84331 4115 84397 4116
rect 84334 3909 84394 4115
rect 84331 3908 84397 3909
rect 84331 3844 84332 3908
rect 84396 3844 84397 3908
rect 84331 3843 84397 3844
rect 84702 3093 84762 123115
rect 84886 122229 84946 185270
rect 84883 122228 84949 122229
rect 84883 122164 84884 122228
rect 84948 122164 84949 122228
rect 84883 122163 84949 122164
rect 85070 121413 85130 186902
rect 85067 121412 85133 121413
rect 85067 121348 85068 121412
rect 85132 121348 85133 121412
rect 85067 121347 85133 121348
rect 85254 119917 85314 187310
rect 85251 119916 85317 119917
rect 85251 119852 85252 119916
rect 85316 119852 85317 119916
rect 85251 119851 85317 119852
rect 85438 6765 85498 191118
rect 85622 118965 85682 196830
rect 85619 118964 85685 118965
rect 85619 118900 85620 118964
rect 85684 118900 85685 118964
rect 85619 118899 85685 118900
rect 85806 62797 85866 198190
rect 86726 197370 86786 203630
rect 86910 197570 86970 204902
rect 87278 204778 87338 205670
rect 87830 205138 87890 212470
rect 88014 208410 88074 213062
rect 88014 208350 88258 208410
rect 87278 204718 87706 204778
rect 86910 197510 87154 197570
rect 85990 197310 86786 197370
rect 85990 116925 86050 197310
rect 86174 195470 86270 195530
rect 86174 192810 86234 195470
rect 86726 194258 86786 196742
rect 86174 192750 86786 192810
rect 86726 192218 86786 192750
rect 87094 191450 87154 197510
rect 86910 191390 87154 191450
rect 86910 186690 86970 191390
rect 87278 191178 87338 202182
rect 87646 202058 87706 204718
rect 87462 201998 87706 202058
rect 87462 201242 87522 201998
rect 87462 201182 87706 201242
rect 87646 196890 87706 201182
rect 86726 186630 86970 186690
rect 87094 191118 87338 191178
rect 87462 196830 87706 196890
rect 86726 186330 86786 186630
rect 86726 186270 86970 186330
rect 86910 186010 86970 186270
rect 87094 186010 87154 191118
rect 87462 186330 87522 196830
rect 87830 196298 87890 201502
rect 88198 195990 88258 208350
rect 88382 195990 88442 212382
rect 88566 195990 88626 213870
rect 87830 195930 88626 195990
rect 88750 213210 88810 218590
rect 88934 213210 88994 220630
rect 88750 213150 88994 213210
rect 87830 195258 87890 195930
rect 88198 195258 88258 195930
rect 88382 195258 88442 195930
rect 87646 195198 88442 195258
rect 87646 190498 87706 195198
rect 87830 190770 87890 195198
rect 88198 192218 88258 195198
rect 87830 190710 88294 190770
rect 87646 190438 88626 190498
rect 88346 190030 88442 190090
rect 86726 185950 87154 186010
rect 87278 186270 87522 186330
rect 86726 181338 86786 185950
rect 86910 184950 86970 185950
rect 87278 184950 87338 186270
rect 88014 186010 88074 187222
rect 88014 185950 88258 186010
rect 86910 184890 87154 184950
rect 87278 184890 87522 184950
rect 87094 180810 87154 184890
rect 87462 180810 87522 184890
rect 88198 184650 88258 185950
rect 88382 184950 88442 190030
rect 88566 184950 88626 190438
rect 88382 184890 88626 184950
rect 88382 184650 88442 184890
rect 87646 184590 88442 184650
rect 87646 181250 87706 184590
rect 88198 182610 88258 184590
rect 88014 182550 88258 182610
rect 88014 181930 88074 182550
rect 88382 181930 88442 184590
rect 87830 181870 88074 181930
rect 88198 181870 88442 181930
rect 87830 181250 87890 181870
rect 88198 181250 88258 181870
rect 87646 181190 88442 181250
rect 87830 180810 87890 181190
rect 88198 180810 88258 181190
rect 86358 180750 87522 180810
rect 87646 180750 88258 180810
rect 86358 175130 86418 180750
rect 87094 180658 87154 180750
rect 87646 180570 87706 180750
rect 87462 180510 87706 180570
rect 86358 175070 86602 175130
rect 86542 173910 86602 175070
rect 86358 173850 86602 173910
rect 86358 171730 86418 173850
rect 86726 173770 86786 180422
rect 87321 179892 87387 179893
rect 87321 179890 87322 179892
rect 86910 179830 87322 179890
rect 86910 174450 86970 179830
rect 87321 179828 87322 179830
rect 87386 179828 87387 179892
rect 87321 179827 87387 179828
rect 87462 178530 87522 180510
rect 87324 178470 87522 178530
rect 87830 178530 87890 180750
rect 87830 178470 88074 178530
rect 87324 177170 87384 178470
rect 88014 177258 88074 178470
rect 87324 177110 87706 177170
rect 87646 176490 87706 177110
rect 87426 176430 87890 176490
rect 87278 174538 87338 175662
rect 86910 174390 87016 174450
rect 86956 173910 87016 174390
rect 86956 173850 87154 173910
rect 86542 173710 86786 173770
rect 87094 173770 87154 173850
rect 87646 173770 87706 176430
rect 87830 173770 87890 176430
rect 88382 174450 88442 181190
rect 88750 180810 88810 213150
rect 88934 180810 88994 213150
rect 88566 180750 88994 180810
rect 88566 179210 88626 180750
rect 88750 179893 88810 180750
rect 88747 179892 88813 179893
rect 88747 179828 88748 179892
rect 88812 179828 88813 179892
rect 88747 179827 88813 179828
rect 88566 179150 88810 179210
rect 88198 174390 88442 174450
rect 88198 173770 88258 174390
rect 87094 173710 88442 173770
rect 86542 172530 86602 173710
rect 86542 172470 86970 172530
rect 86358 171670 86602 171730
rect 86542 171150 86602 171670
rect 86174 171090 86602 171150
rect 86174 170370 86234 171090
rect 86910 171050 86970 172470
rect 87094 171150 87154 172942
rect 87472 172262 87522 172410
rect 87462 171866 87522 172262
rect 87324 171806 87522 171866
rect 87324 171597 87384 171806
rect 87646 171730 87706 173710
rect 87462 171670 87706 171730
rect 87321 171596 87387 171597
rect 87321 171532 87322 171596
rect 87386 171532 87387 171596
rect 87321 171531 87387 171532
rect 87094 171090 87292 171150
rect 86910 170990 87016 171050
rect 86956 170370 87016 170990
rect 87232 170370 87292 171090
rect 87462 170370 87522 171670
rect 87643 171596 87709 171597
rect 87643 171532 87644 171596
rect 87708 171532 87709 171596
rect 87643 171531 87709 171532
rect 87646 170370 87706 171531
rect 87830 170370 87890 173710
rect 88198 172410 88258 173710
rect 88014 172350 88258 172410
rect 88014 170370 88074 172350
rect 88382 170458 88442 173710
rect 88750 173090 88810 179150
rect 89118 177170 89178 226478
rect 88934 177110 89178 177170
rect 88934 175810 88994 177110
rect 89302 176670 89362 226478
rect 89486 176670 89546 582795
rect 89118 176610 89546 176670
rect 89118 175810 89178 176610
rect 89302 176490 89362 176610
rect 89302 176430 89546 176490
rect 88934 175750 89362 175810
rect 89118 173858 89178 175750
rect 88750 173030 89132 173090
rect 89072 172410 89132 173030
rect 89072 172350 89178 172410
rect 86174 170310 87154 170370
rect 87232 170310 87338 170370
rect 87462 170310 88212 170370
rect 86956 170098 87016 170310
rect 86910 170038 87016 170098
rect 86910 169282 86970 170038
rect 86358 169222 86970 169282
rect 86358 163658 86418 169222
rect 87094 169010 87154 170310
rect 86956 168950 87154 169010
rect 86726 155410 86786 168862
rect 86956 168738 87016 168950
rect 86956 168678 87154 168738
rect 87094 166290 87154 168678
rect 87278 166290 87338 170310
rect 87646 169282 87706 170310
rect 87830 170098 87890 170310
rect 88014 170098 88074 170310
rect 88152 170098 88212 170310
rect 87830 170038 88442 170098
rect 87508 169222 87706 169282
rect 87508 169146 87568 169222
rect 88014 169146 88074 170038
rect 88152 169770 88212 170038
rect 88152 169710 88258 169770
rect 87462 169086 88074 169146
rect 88198 169146 88258 169710
rect 88382 169282 88442 170038
rect 88750 169778 88810 172262
rect 88382 169222 88994 169282
rect 88198 169086 88442 169146
rect 87462 169010 87568 169086
rect 87462 168950 88074 169010
rect 87462 168738 87522 168950
rect 87462 168678 87890 168738
rect 87462 166378 87522 168182
rect 86910 166230 87338 166290
rect 86910 156090 86970 166230
rect 87094 165610 87154 166230
rect 87094 165550 87522 165610
rect 87094 164782 87144 164930
rect 87094 162890 87154 164782
rect 87462 164658 87522 165550
rect 87830 164930 87890 168678
rect 87278 164598 87522 164658
rect 87646 164870 87890 164930
rect 87278 163026 87338 164598
rect 87646 163658 87706 164870
rect 87278 162966 87522 163026
rect 87462 162890 87522 162966
rect 88014 162890 88074 168950
rect 88382 167650 88442 169086
rect 88336 167590 88442 167650
rect 88566 168862 88616 169010
rect 88336 166426 88396 167590
rect 88198 166366 88396 166426
rect 88566 166378 88626 168862
rect 88198 162890 88258 166366
rect 88934 165610 88994 169222
rect 88796 165550 88994 165610
rect 88566 164930 88626 165462
rect 88336 164870 88626 164930
rect 88336 164658 88396 164870
rect 88796 164658 88856 165550
rect 89118 164930 89178 172350
rect 88336 164598 88442 164658
rect 88382 162890 88442 164598
rect 88566 164598 88856 164658
rect 88934 164870 89178 164930
rect 88566 163658 88626 164598
rect 88566 163510 88616 163658
rect 88934 163026 88994 164870
rect 89302 164658 89362 175750
rect 89118 164598 89362 164658
rect 89118 163570 89178 164598
rect 89486 163570 89546 176430
rect 89072 163510 89178 163570
rect 89348 163510 89546 163570
rect 89072 163026 89132 163510
rect 89348 163026 89408 163510
rect 88566 162966 89546 163026
rect 88566 162890 88626 162966
rect 87094 162830 88626 162890
rect 87462 162210 87522 162830
rect 87462 162150 87890 162210
rect 87278 160850 87338 161382
rect 87094 160790 87338 160850
rect 87094 157450 87154 160790
rect 87610 160110 87706 160170
rect 87094 157390 87338 157450
rect 87278 156090 87338 157390
rect 86910 156030 87338 156090
rect 86910 155410 86970 156030
rect 87094 155410 87154 156030
rect 86726 155350 87522 155410
rect 86910 154590 86970 155350
rect 86726 154530 86970 154590
rect 86726 137818 86786 154530
rect 87094 143938 87154 155350
rect 87462 153210 87522 155350
rect 87646 153210 87706 160110
rect 87830 153210 87890 162150
rect 88014 153210 88074 162830
rect 88198 153210 88258 162830
rect 88382 153210 88442 162830
rect 88750 154730 88810 162062
rect 88566 154670 88810 154730
rect 88566 153210 88626 154670
rect 87462 153150 88810 153210
rect 87094 141946 87154 142342
rect 87094 141886 87338 141946
rect 87278 137594 87338 141886
rect 87094 137534 87338 137594
rect 87094 137322 87154 137534
rect 86726 137262 87154 137322
rect 86726 135690 86786 137262
rect 87094 136370 87154 136902
rect 87094 136310 87522 136370
rect 86726 135630 87338 135690
rect 86726 123997 86786 132822
rect 86723 123996 86789 123997
rect 86723 123932 86724 123996
rect 86788 123932 86789 123996
rect 86723 123931 86789 123932
rect 86171 123452 86237 123453
rect 86171 123388 86172 123452
rect 86236 123388 86237 123452
rect 87278 123450 87338 135630
rect 87462 123589 87522 136310
rect 87459 123588 87525 123589
rect 87459 123524 87460 123588
rect 87524 123524 87525 123588
rect 87459 123523 87525 123524
rect 87278 123390 87522 123450
rect 86171 123387 86237 123388
rect 85987 116924 86053 116925
rect 85987 116860 85988 116924
rect 86052 116860 86053 116924
rect 85987 116859 86053 116860
rect 85987 106452 86053 106453
rect 85987 106388 85988 106452
rect 86052 106388 86053 106452
rect 85987 106387 86053 106388
rect 85990 105909 86050 106387
rect 85987 105908 86053 105909
rect 85987 105844 85988 105908
rect 86052 105844 86053 105908
rect 85987 105843 86053 105844
rect 85987 105772 86053 105773
rect 85987 105708 85988 105772
rect 86052 105708 86053 105772
rect 85987 105707 86053 105708
rect 85990 67285 86050 105707
rect 85987 67284 86053 67285
rect 85987 67220 85988 67284
rect 86052 67220 86053 67284
rect 85987 67219 86053 67220
rect 85987 67148 86053 67149
rect 85987 67084 85988 67148
rect 86052 67084 86053 67148
rect 85987 67083 86053 67084
rect 85803 62796 85869 62797
rect 85803 62732 85804 62796
rect 85868 62732 85869 62796
rect 85803 62731 85869 62732
rect 85803 48380 85869 48381
rect 85803 48316 85804 48380
rect 85868 48316 85869 48380
rect 85803 48315 85869 48316
rect 85806 43485 85866 48315
rect 85990 48109 86050 67083
rect 85987 48108 86053 48109
rect 85987 48044 85988 48108
rect 86052 48044 86053 48108
rect 85987 48043 86053 48044
rect 85987 47836 86053 47837
rect 85987 47772 85988 47836
rect 86052 47772 86053 47836
rect 85987 47771 86053 47772
rect 85803 43484 85869 43485
rect 85803 43420 85804 43484
rect 85868 43420 85869 43484
rect 85803 43419 85869 43420
rect 85803 37364 85869 37365
rect 85803 37300 85804 37364
rect 85868 37300 85869 37364
rect 85803 37299 85869 37300
rect 85806 27573 85866 37299
rect 85803 27572 85869 27573
rect 85803 27508 85804 27572
rect 85868 27508 85869 27572
rect 85803 27507 85869 27508
rect 85990 19277 86050 47771
rect 85987 19276 86053 19277
rect 85987 19212 85988 19276
rect 86052 19212 86053 19276
rect 85987 19211 86053 19212
rect 85619 18052 85685 18053
rect 85619 17988 85620 18052
rect 85684 17988 85685 18052
rect 85619 17987 85685 17988
rect 85622 9893 85682 17987
rect 85619 9892 85685 9893
rect 85619 9828 85620 9892
rect 85684 9828 85685 9892
rect 85619 9827 85685 9828
rect 85803 9756 85869 9757
rect 85803 9692 85804 9756
rect 85868 9692 85869 9756
rect 85803 9691 85869 9692
rect 85987 9756 86053 9757
rect 85987 9692 85988 9756
rect 86052 9692 86053 9756
rect 85987 9691 86053 9692
rect 85806 8261 85866 9691
rect 85990 9485 86050 9691
rect 85987 9484 86053 9485
rect 85987 9420 85988 9484
rect 86052 9420 86053 9484
rect 85987 9419 86053 9420
rect 85803 8260 85869 8261
rect 85803 8196 85804 8260
rect 85868 8196 85869 8260
rect 85803 8195 85869 8196
rect 85435 6764 85501 6765
rect 85435 6700 85436 6764
rect 85500 6700 85501 6764
rect 85435 6699 85501 6700
rect 86174 4725 86234 123387
rect 86907 123044 86973 123045
rect 86907 122980 86908 123044
rect 86972 122980 86973 123044
rect 86907 122979 86973 122980
rect 86910 116789 86970 122979
rect 87275 122092 87341 122093
rect 87275 122028 87276 122092
rect 87340 122028 87341 122092
rect 87275 122027 87341 122028
rect 86907 116788 86973 116789
rect 86907 116724 86908 116788
rect 86972 116724 86973 116788
rect 86907 116723 86973 116724
rect 87278 111213 87338 122027
rect 87275 111212 87341 111213
rect 87275 111148 87276 111212
rect 87340 111148 87341 111212
rect 87275 111147 87341 111148
rect 86723 106996 86789 106997
rect 86723 106932 86724 106996
rect 86788 106932 86789 106996
rect 86723 106931 86789 106932
rect 86726 40221 86786 106931
rect 87091 105908 87157 105909
rect 87091 105844 87092 105908
rect 87156 105844 87157 105908
rect 87091 105843 87157 105844
rect 87094 86325 87154 105843
rect 87091 86324 87157 86325
rect 87091 86260 87092 86324
rect 87156 86260 87157 86324
rect 87091 86259 87157 86260
rect 87462 84285 87522 123390
rect 87646 121410 87706 153150
rect 87830 122637 87890 153150
rect 87827 122636 87893 122637
rect 87827 122572 87828 122636
rect 87892 122572 87893 122636
rect 87827 122571 87893 122572
rect 87646 121350 87890 121410
rect 87830 119237 87890 121350
rect 87827 119236 87893 119237
rect 87827 119172 87828 119236
rect 87892 119172 87893 119236
rect 87827 119171 87893 119172
rect 88014 115429 88074 153150
rect 88198 120733 88258 153150
rect 88382 123997 88442 153150
rect 88379 123996 88445 123997
rect 88379 123932 88380 123996
rect 88444 123932 88445 123996
rect 88379 123931 88445 123932
rect 88566 123317 88626 153150
rect 88563 123316 88629 123317
rect 88563 123252 88564 123316
rect 88628 123252 88629 123316
rect 88563 123251 88629 123252
rect 88750 122770 88810 153150
rect 88934 123045 88994 162966
rect 89072 162890 89132 162966
rect 89348 162890 89408 162966
rect 89072 162830 89178 162890
rect 88931 123044 88997 123045
rect 88931 122980 88932 123044
rect 88996 122980 88997 123044
rect 88931 122979 88997 122980
rect 88931 122772 88997 122773
rect 88931 122770 88932 122772
rect 88750 122710 88932 122770
rect 88931 122708 88932 122710
rect 88996 122708 88997 122772
rect 88931 122707 88997 122708
rect 88195 120732 88261 120733
rect 88195 120668 88196 120732
rect 88260 120668 88261 120732
rect 88195 120667 88261 120668
rect 88011 115428 88077 115429
rect 88011 115364 88012 115428
rect 88076 115364 88077 115428
rect 88011 115363 88077 115364
rect 88379 115428 88445 115429
rect 88379 115364 88380 115428
rect 88444 115364 88445 115428
rect 88379 115363 88445 115364
rect 88382 106538 88442 115363
rect 88382 101690 88442 105622
rect 88014 101630 88442 101690
rect 88014 96389 88074 101630
rect 88195 101556 88261 101557
rect 88195 101492 88196 101556
rect 88260 101492 88261 101556
rect 88195 101491 88261 101492
rect 88198 96525 88258 101491
rect 88195 96524 88261 96525
rect 88195 96460 88196 96524
rect 88260 96460 88261 96524
rect 88195 96459 88261 96460
rect 88011 96388 88077 96389
rect 88011 96324 88012 96388
rect 88076 96324 88077 96388
rect 88011 96323 88077 96324
rect 88195 94620 88261 94621
rect 88195 94556 88196 94620
rect 88260 94556 88261 94620
rect 88195 94555 88261 94556
rect 88011 92716 88077 92717
rect 88011 92652 88012 92716
rect 88076 92652 88077 92716
rect 88011 92651 88077 92652
rect 88014 92445 88074 92651
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88198 92170 88258 94555
rect 87646 92110 88258 92170
rect 87646 88365 87706 92110
rect 88011 92036 88077 92037
rect 88011 91972 88012 92036
rect 88076 91972 88077 92036
rect 88011 91971 88077 91972
rect 87643 88364 87709 88365
rect 87643 88300 87644 88364
rect 87708 88300 87709 88364
rect 87643 88299 87709 88300
rect 87459 84284 87525 84285
rect 87459 84220 87460 84284
rect 87524 84220 87525 84284
rect 87459 84219 87525 84220
rect 87643 84284 87709 84285
rect 87643 84220 87644 84284
rect 87708 84220 87709 84284
rect 87643 84219 87709 84220
rect 87646 78029 87706 84219
rect 88014 84149 88074 91971
rect 88195 88364 88261 88365
rect 88195 88300 88196 88364
rect 88260 88300 88261 88364
rect 88195 88299 88261 88300
rect 88011 84148 88077 84149
rect 88011 84084 88012 84148
rect 88076 84084 88077 84148
rect 88011 84083 88077 84084
rect 88011 83876 88077 83877
rect 88011 83812 88012 83876
rect 88076 83812 88077 83876
rect 88011 83811 88077 83812
rect 87091 78028 87157 78029
rect 87091 77964 87092 78028
rect 87156 77964 87157 78028
rect 87091 77963 87157 77964
rect 87643 78028 87709 78029
rect 87643 77964 87644 78028
rect 87708 77964 87709 78028
rect 87643 77963 87709 77964
rect 86723 40220 86789 40221
rect 86723 40156 86724 40220
rect 86788 40156 86789 40220
rect 86723 40155 86789 40156
rect 86539 39948 86605 39949
rect 86539 39884 86540 39948
rect 86604 39884 86605 39948
rect 86539 39883 86605 39884
rect 86542 22813 86602 39883
rect 86539 22812 86605 22813
rect 86539 22748 86540 22812
rect 86604 22748 86605 22812
rect 86539 22747 86605 22748
rect 86171 4724 86237 4725
rect 86171 4660 86172 4724
rect 86236 4660 86237 4724
rect 86171 4659 86237 4660
rect 86355 4180 86421 4181
rect 86355 4116 86356 4180
rect 86420 4116 86421 4180
rect 86355 4115 86421 4116
rect 86358 3773 86418 4115
rect 87094 3773 87154 77963
rect 87643 67692 87709 67693
rect 87643 67628 87644 67692
rect 87708 67628 87709 67692
rect 87643 67627 87709 67628
rect 87646 62253 87706 67627
rect 87643 62252 87709 62253
rect 87643 62188 87644 62252
rect 87708 62188 87709 62252
rect 87643 62187 87709 62188
rect 87459 61980 87525 61981
rect 87459 61916 87460 61980
rect 87524 61916 87525 61980
rect 87459 61915 87525 61916
rect 87462 57901 87522 61915
rect 87459 57900 87525 57901
rect 87459 57836 87460 57900
rect 87524 57836 87525 57900
rect 87459 57835 87525 57836
rect 87459 48380 87525 48381
rect 87459 48316 87460 48380
rect 87524 48316 87525 48380
rect 87459 48315 87525 48316
rect 87462 40221 87522 48315
rect 87459 40220 87525 40221
rect 87459 40156 87460 40220
rect 87524 40156 87525 40220
rect 87459 40155 87525 40156
rect 87275 39948 87341 39949
rect 87275 39884 87276 39948
rect 87340 39884 87341 39948
rect 87275 39883 87341 39884
rect 87278 35325 87338 39883
rect 87275 35324 87341 35325
rect 87275 35260 87276 35324
rect 87340 35260 87341 35324
rect 87275 35259 87341 35260
rect 87459 23492 87525 23493
rect 87459 23428 87460 23492
rect 87524 23428 87525 23492
rect 87459 23427 87525 23428
rect 87462 18733 87522 23427
rect 87459 18732 87525 18733
rect 87459 18668 87460 18732
rect 87524 18668 87525 18732
rect 87459 18667 87525 18668
rect 88014 6085 88074 83811
rect 88198 78029 88258 88299
rect 88195 78028 88261 78029
rect 88195 77964 88196 78028
rect 88260 77964 88261 78028
rect 88195 77963 88261 77964
rect 88195 69188 88261 69189
rect 88195 69124 88196 69188
rect 88260 69124 88261 69188
rect 88195 69123 88261 69124
rect 88011 6084 88077 6085
rect 88011 6020 88012 6084
rect 88076 6020 88077 6084
rect 88011 6019 88077 6020
rect 86355 3772 86421 3773
rect 86355 3708 86356 3772
rect 86420 3708 86421 3772
rect 86355 3707 86421 3708
rect 87091 3772 87157 3773
rect 87091 3708 87092 3772
rect 87156 3708 87157 3772
rect 87091 3707 87157 3708
rect 88198 3637 88258 69123
rect 89118 3909 89178 162830
rect 89302 162830 89408 162890
rect 89302 122773 89362 162830
rect 89299 122772 89365 122773
rect 89299 122708 89300 122772
rect 89364 122708 89365 122772
rect 89299 122707 89365 122708
rect 89486 122637 89546 162966
rect 89483 122636 89549 122637
rect 89483 122572 89484 122636
rect 89548 122572 89549 122636
rect 89483 122571 89549 122572
rect 89299 122364 89365 122365
rect 89299 122300 89300 122364
rect 89364 122300 89365 122364
rect 89299 122299 89365 122300
rect 89302 5269 89362 122299
rect 89670 121549 89730 584971
rect 89851 582044 89917 582045
rect 89851 581980 89852 582044
rect 89916 581980 89917 582044
rect 89851 581979 89917 581980
rect 89667 121548 89733 121549
rect 89667 121484 89668 121548
rect 89732 121484 89733 121548
rect 89667 121483 89733 121484
rect 89854 119101 89914 581979
rect 90035 581364 90101 581365
rect 90035 581300 90036 581364
rect 90100 581300 90101 581364
rect 90035 581299 90101 581300
rect 90038 122501 90098 581299
rect 90035 122500 90101 122501
rect 90035 122436 90036 122500
rect 90100 122436 90101 122500
rect 90035 122435 90101 122436
rect 90222 121277 90282 699755
rect 90804 668454 91404 705202
rect 92243 700772 92309 700773
rect 92243 700708 92244 700772
rect 92308 700708 92309 700772
rect 92243 700707 92309 700708
rect 91875 700364 91941 700365
rect 91875 700300 91876 700364
rect 91940 700300 91941 700364
rect 91875 700299 91941 700300
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 582000 91404 595898
rect 91691 584764 91757 584765
rect 91691 584700 91692 584764
rect 91756 584700 91757 584764
rect 91691 584699 91757 584700
rect 91694 581909 91754 584699
rect 91323 581908 91389 581909
rect 91323 581844 91324 581908
rect 91388 581844 91389 581908
rect 91323 581843 91389 581844
rect 91691 581908 91757 581909
rect 91691 581844 91692 581908
rect 91756 581844 91757 581908
rect 91691 581843 91757 581844
rect 90587 581364 90653 581365
rect 90587 581300 90588 581364
rect 90652 581300 90653 581364
rect 90587 581299 90653 581300
rect 90403 579868 90469 579869
rect 90403 579804 90404 579868
rect 90468 579804 90469 579868
rect 90403 579803 90469 579804
rect 90406 545130 90466 579803
rect 90590 545130 90650 581299
rect 91139 580276 91205 580277
rect 91139 580212 91140 580276
rect 91204 580212 91205 580276
rect 91139 580211 91205 580212
rect 90406 545070 90834 545130
rect 90590 526010 90650 545070
rect 90774 526010 90834 545070
rect 90406 525950 90834 526010
rect 90406 216610 90466 525950
rect 90590 263530 90650 525950
rect 90590 263470 91018 263530
rect 90958 254690 91018 263470
rect 90774 254630 91018 254690
rect 90774 254010 90834 254630
rect 90590 253950 90834 254010
rect 90590 217970 90650 253950
rect 90590 217910 90834 217970
rect 90406 216550 90650 216610
rect 90590 215338 90650 216550
rect 90774 215930 90834 217910
rect 90774 215870 91018 215930
rect 90958 214570 91018 215870
rect 90406 214510 91018 214570
rect 90406 213210 90466 214510
rect 90406 213150 90650 213210
rect 90590 201650 90650 213150
rect 90774 201650 90834 213742
rect 90406 201590 90834 201650
rect 90406 181930 90466 201590
rect 90590 190362 90650 201590
rect 90590 190302 90834 190362
rect 90774 181930 90834 190302
rect 90406 181870 90650 181930
rect 90774 181870 91018 181930
rect 90590 181338 90650 181870
rect 90958 179890 91018 181870
rect 90406 179830 91018 179890
rect 90406 170370 90466 179830
rect 90774 177170 90834 178382
rect 90774 177110 91018 177170
rect 90406 170310 90502 170370
rect 90958 170098 91018 177110
rect 90406 170038 91018 170098
rect 90219 121276 90285 121277
rect 90219 121212 90220 121276
rect 90284 121212 90285 121276
rect 90219 121211 90285 121212
rect 89851 119100 89917 119101
rect 89851 119036 89852 119100
rect 89916 119036 89917 119100
rect 89851 119035 89917 119036
rect 89299 5268 89365 5269
rect 89299 5204 89300 5268
rect 89364 5204 89365 5268
rect 89299 5203 89365 5204
rect 90406 5133 90466 170038
rect 90774 164930 90834 169542
rect 90590 164870 90834 164930
rect 90590 122637 90650 164870
rect 90771 123996 90837 123997
rect 90771 123932 90772 123996
rect 90836 123932 90837 123996
rect 90771 123931 90837 123932
rect 90955 123996 91021 123997
rect 90955 123932 90956 123996
rect 91020 123932 91021 123996
rect 90955 123931 91021 123932
rect 90587 122636 90653 122637
rect 90587 122572 90588 122636
rect 90652 122572 90653 122636
rect 90587 122571 90653 122572
rect 90774 122498 90834 123931
rect 90958 123725 91018 123931
rect 91142 123725 91202 580211
rect 90955 123724 91021 123725
rect 90955 123660 90956 123724
rect 91020 123660 91021 123724
rect 90955 123659 91021 123660
rect 91139 123724 91205 123725
rect 91139 123660 91140 123724
rect 91204 123660 91205 123724
rect 91139 123659 91205 123660
rect 91326 122773 91386 581843
rect 91691 581364 91757 581365
rect 91691 581300 91692 581364
rect 91756 581300 91757 581364
rect 91691 581299 91757 581300
rect 91507 580140 91573 580141
rect 91507 580076 91508 580140
rect 91572 580076 91573 580140
rect 91507 580075 91573 580076
rect 91323 122772 91389 122773
rect 91323 122708 91324 122772
rect 91388 122708 91389 122772
rect 91323 122707 91389 122708
rect 90590 122438 90834 122498
rect 90590 121957 90650 122438
rect 91510 122093 91570 580075
rect 91507 122092 91573 122093
rect 91507 122028 91508 122092
rect 91572 122028 91573 122092
rect 91507 122027 91573 122028
rect 90587 121956 90653 121957
rect 90587 121892 90588 121956
rect 90652 121892 90653 121956
rect 90587 121891 90653 121892
rect 90804 92454 91404 122000
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90403 5132 90469 5133
rect 90403 5068 90404 5132
rect 90468 5068 90469 5132
rect 90403 5067 90469 5068
rect 89115 3908 89181 3909
rect 89115 3844 89116 3908
rect 89180 3844 89181 3908
rect 89115 3843 89181 3844
rect 88195 3636 88261 3637
rect 88195 3572 88196 3636
rect 88260 3572 88261 3636
rect 88195 3571 88261 3572
rect 84699 3092 84765 3093
rect 84699 3028 84700 3092
rect 84764 3028 84765 3092
rect 84699 3027 84765 3028
rect 90804 -1266 91404 19898
rect 91694 8941 91754 581299
rect 91878 122637 91938 700299
rect 92059 583812 92125 583813
rect 92059 583748 92060 583812
rect 92124 583748 92125 583812
rect 92059 583747 92125 583748
rect 91875 122636 91941 122637
rect 91875 122572 91876 122636
rect 91940 122572 91941 122636
rect 91875 122571 91941 122572
rect 91691 8940 91757 8941
rect 91691 8876 91692 8940
rect 91756 8876 91757 8940
rect 91691 8875 91757 8876
rect 92062 5949 92122 583747
rect 92246 119645 92306 700707
rect 93347 700500 93413 700501
rect 93347 700436 93348 700500
rect 93412 700436 93413 700500
rect 93347 700435 93413 700436
rect 92611 584084 92677 584085
rect 92611 584020 92612 584084
rect 92676 584020 92677 584084
rect 92611 584019 92677 584020
rect 92427 581364 92493 581365
rect 92427 581300 92428 581364
rect 92492 581300 92493 581364
rect 92427 581299 92493 581300
rect 92243 119644 92309 119645
rect 92243 119580 92244 119644
rect 92308 119580 92309 119644
rect 92243 119579 92309 119580
rect 92059 5948 92125 5949
rect 92059 5884 92060 5948
rect 92124 5884 92125 5948
rect 92059 5883 92125 5884
rect 92430 3909 92490 581299
rect 92614 580410 92674 584019
rect 92614 580350 92858 580410
rect 92611 579868 92677 579869
rect 92611 579804 92612 579868
rect 92676 579804 92677 579868
rect 92611 579803 92677 579804
rect 92614 123453 92674 579803
rect 92611 123452 92677 123453
rect 92611 123388 92612 123452
rect 92676 123388 92677 123452
rect 92611 123387 92677 123388
rect 92611 123044 92677 123045
rect 92611 122980 92612 123044
rect 92676 122980 92677 123044
rect 92611 122979 92677 122980
rect 92614 118829 92674 122979
rect 92798 122365 92858 580350
rect 92795 122364 92861 122365
rect 92795 122300 92796 122364
rect 92860 122300 92861 122364
rect 92795 122299 92861 122300
rect 92611 118828 92677 118829
rect 92611 118764 92612 118828
rect 92676 118764 92677 118828
rect 92611 118763 92677 118764
rect 92982 5405 93042 583662
rect 93163 581364 93229 581365
rect 93163 581300 93164 581364
rect 93228 581300 93229 581364
rect 93163 581299 93229 581300
rect 93166 6901 93226 581299
rect 93350 119781 93410 700435
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 93531 583812 93597 583813
rect 93531 583748 93532 583812
rect 93596 583748 93597 583812
rect 93531 583747 93597 583748
rect 93347 119780 93413 119781
rect 93347 119716 93348 119780
rect 93412 119716 93413 119780
rect 93347 119715 93413 119716
rect 93163 6900 93229 6901
rect 93163 6836 93164 6900
rect 93228 6836 93229 6900
rect 93163 6835 93229 6836
rect 92979 5404 93045 5405
rect 92979 5340 92980 5404
rect 93044 5340 93045 5404
rect 92979 5339 93045 5340
rect 93534 3909 93594 583747
rect 93718 580141 93778 584342
rect 94404 582000 95004 599498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 97763 584492 97829 584493
rect 97763 584428 97764 584492
rect 97828 584428 97829 584492
rect 97763 584427 97829 584428
rect 94267 581228 94333 581229
rect 94267 581164 94268 581228
rect 94332 581164 94333 581228
rect 94267 581163 94333 581164
rect 94270 580957 94330 581163
rect 94267 580956 94333 580957
rect 94267 580892 94268 580956
rect 94332 580892 94333 580956
rect 94267 580891 94333 580892
rect 93715 580140 93781 580141
rect 93715 580076 93716 580140
rect 93780 580076 93781 580140
rect 93715 580075 93781 580076
rect 94086 580005 94146 580262
rect 94083 580004 94149 580005
rect 94083 579940 94084 580004
rect 94148 579940 94149 580004
rect 94083 579939 94149 579940
rect 97766 579869 97826 584427
rect 98004 582000 98604 603098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 582000 102204 606698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 106043 582860 106109 582861
rect 106043 582796 106044 582860
rect 106108 582796 106109 582860
rect 106043 582795 106109 582796
rect 104387 581228 104453 581229
rect 104387 581164 104388 581228
rect 104452 581164 104453 581228
rect 104387 581163 104453 581164
rect 104390 580957 104450 581163
rect 104387 580956 104453 580957
rect 104387 580892 104388 580956
rect 104452 580892 104453 580956
rect 104387 580891 104453 580892
rect 99971 580548 100037 580549
rect 99971 580498 99972 580548
rect 100036 580498 100037 580548
rect 106046 580498 106106 582795
rect 108804 582000 109404 613898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582000 113004 617498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 113771 582316 113837 582317
rect 113771 582252 113772 582316
rect 113836 582252 113837 582316
rect 113771 582251 113837 582252
rect 108806 581710 109234 581770
rect 108806 581229 108866 581710
rect 108987 581636 109053 581637
rect 108987 581572 108988 581636
rect 109052 581572 109053 581636
rect 108987 581571 109053 581572
rect 108803 581228 108869 581229
rect 108803 581164 108804 581228
rect 108868 581164 108869 581228
rect 108803 581163 108869 581164
rect 108990 581090 109050 581571
rect 109174 581362 109234 581710
rect 113587 581500 113653 581501
rect 113587 581436 113588 581500
rect 113652 581436 113653 581500
rect 113587 581435 113653 581436
rect 109355 581364 109421 581365
rect 109355 581362 109356 581364
rect 109174 581302 109356 581362
rect 109355 581300 109356 581302
rect 109420 581300 109421 581364
rect 109355 581299 109421 581300
rect 113590 581093 113650 581435
rect 113774 581093 113834 582251
rect 116004 582000 116604 585098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 582000 120204 588698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 582000 127404 595898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 582000 131004 599498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 582000 134604 603098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 582000 138204 606698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 582000 145404 613898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582000 149004 617498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 151675 582044 151741 582045
rect 151675 581980 151676 582044
rect 151740 581980 151741 582044
rect 152004 582000 152604 585098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 582000 156204 588698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162347 582316 162413 582317
rect 162347 582252 162348 582316
rect 162412 582252 162413 582316
rect 162347 582251 162413 582252
rect 156459 582044 156525 582045
rect 151675 581979 151741 581980
rect 156459 581980 156460 582044
rect 156524 581980 156525 582044
rect 156459 581979 156525 581980
rect 128123 581636 128189 581637
rect 128123 581572 128124 581636
rect 128188 581572 128189 581636
rect 128123 581571 128189 581572
rect 128307 581636 128373 581637
rect 128307 581572 128308 581636
rect 128372 581572 128373 581636
rect 128307 581571 128373 581572
rect 137875 581636 137941 581637
rect 137875 581572 137876 581636
rect 137940 581572 137941 581636
rect 137875 581571 137941 581572
rect 123339 581500 123405 581501
rect 123339 581436 123340 581500
rect 123404 581436 123405 581500
rect 123339 581435 123405 581436
rect 118555 581228 118621 581229
rect 118555 581164 118556 581228
rect 118620 581164 118621 581228
rect 118555 581163 118621 581164
rect 109355 581092 109421 581093
rect 109355 581090 109356 581092
rect 108990 581030 109356 581090
rect 109355 581028 109356 581030
rect 109420 581028 109421 581092
rect 109355 581027 109421 581028
rect 113587 581092 113653 581093
rect 113587 581028 113588 581092
rect 113652 581028 113653 581092
rect 113587 581027 113653 581028
rect 113771 581092 113837 581093
rect 113771 581028 113772 581092
rect 113836 581028 113837 581092
rect 113771 581027 113837 581028
rect 118558 580821 118618 581163
rect 123342 581093 123402 581435
rect 128126 581093 128186 581571
rect 128310 581093 128370 581571
rect 137323 581228 137389 581229
rect 137323 581164 137324 581228
rect 137388 581164 137389 581228
rect 137323 581163 137389 581164
rect 123339 581092 123405 581093
rect 123339 581028 123340 581092
rect 123404 581028 123405 581092
rect 123339 581027 123405 581028
rect 128123 581092 128189 581093
rect 128123 581028 128124 581092
rect 128188 581028 128189 581092
rect 128123 581027 128189 581028
rect 128307 581092 128373 581093
rect 128307 581028 128308 581092
rect 128372 581028 128373 581092
rect 128307 581027 128373 581028
rect 137326 580957 137386 581163
rect 137507 581092 137573 581093
rect 137507 581028 137508 581092
rect 137572 581090 137573 581092
rect 137878 581090 137938 581571
rect 151678 581229 151738 581979
rect 156091 581364 156157 581365
rect 156091 581300 156092 581364
rect 156156 581300 156157 581364
rect 156091 581299 156157 581300
rect 151675 581228 151741 581229
rect 151675 581164 151676 581228
rect 151740 581164 151741 581228
rect 151675 581163 151741 581164
rect 156094 581093 156154 581299
rect 156462 581229 156522 581979
rect 157195 581636 157261 581637
rect 157195 581572 157196 581636
rect 157260 581572 157261 581636
rect 157195 581571 157261 581572
rect 156459 581228 156525 581229
rect 156459 581164 156460 581228
rect 156524 581164 156525 581228
rect 156459 581163 156525 581164
rect 157198 581093 157258 581571
rect 162350 581229 162410 582251
rect 162804 582000 163404 595898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 582000 167004 599498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 582000 170604 603098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 172470 585110 172714 585170
rect 172470 584901 172530 585110
rect 172467 584900 172533 584901
rect 172467 584836 172468 584900
rect 172532 584836 172533 584900
rect 172467 584835 172533 584836
rect 172654 584765 172714 585110
rect 172651 584764 172717 584765
rect 172651 584700 172652 584764
rect 172716 584700 172717 584764
rect 172651 584699 172717 584700
rect 173604 582000 174204 606698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 582000 181404 613898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 181667 582316 181733 582317
rect 181667 582252 181668 582316
rect 181732 582252 181733 582316
rect 181667 582251 181733 582252
rect 181670 581229 181730 582251
rect 184404 582000 185004 617498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 582000 188604 585098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 190683 582316 190749 582317
rect 190683 582252 190684 582316
rect 190748 582252 190749 582316
rect 190683 582251 190749 582252
rect 186267 581636 186333 581637
rect 186267 581572 186268 581636
rect 186332 581572 186333 581636
rect 186267 581571 186333 581572
rect 186270 581229 186330 581571
rect 190686 581229 190746 582251
rect 191604 582000 192204 588698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 582000 199404 595898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 200987 582316 201053 582317
rect 200987 582252 200988 582316
rect 201052 582252 201053 582316
rect 200987 582251 201053 582252
rect 195835 581636 195901 581637
rect 195835 581572 195836 581636
rect 195900 581572 195901 581636
rect 195835 581571 195901 581572
rect 191051 581500 191117 581501
rect 191051 581436 191052 581500
rect 191116 581436 191117 581500
rect 191051 581435 191117 581436
rect 161427 581228 161493 581229
rect 161427 581164 161428 581228
rect 161492 581164 161493 581228
rect 161427 581163 161493 581164
rect 162347 581228 162413 581229
rect 162347 581164 162348 581228
rect 162412 581164 162413 581228
rect 162347 581163 162413 581164
rect 181667 581228 181733 581229
rect 181667 581164 181668 581228
rect 181732 581164 181733 581228
rect 181667 581163 181733 581164
rect 186267 581228 186333 581229
rect 186267 581164 186268 581228
rect 186332 581164 186333 581228
rect 186267 581163 186333 581164
rect 190499 581228 190565 581229
rect 190499 581164 190500 581228
rect 190564 581164 190565 581228
rect 190499 581163 190565 581164
rect 190683 581228 190749 581229
rect 190683 581164 190684 581228
rect 190748 581164 190749 581228
rect 190683 581163 190749 581164
rect 137572 581030 137938 581090
rect 138059 581092 138125 581093
rect 137572 581028 137573 581030
rect 137507 581027 137573 581028
rect 138059 581028 138060 581092
rect 138124 581090 138125 581092
rect 138427 581092 138493 581093
rect 138427 581090 138428 581092
rect 138124 581030 138428 581090
rect 138124 581028 138125 581030
rect 138059 581027 138125 581028
rect 138427 581028 138428 581030
rect 138492 581028 138493 581092
rect 138427 581027 138493 581028
rect 156091 581092 156157 581093
rect 156091 581028 156092 581092
rect 156156 581028 156157 581092
rect 156091 581027 156157 581028
rect 157195 581092 157261 581093
rect 157195 581028 157196 581092
rect 157260 581028 157261 581092
rect 157195 581027 157261 581028
rect 137323 580956 137389 580957
rect 137323 580892 137324 580956
rect 137388 580892 137389 580956
rect 137323 580891 137389 580892
rect 118555 580820 118621 580821
rect 118555 580756 118556 580820
rect 118620 580756 118621 580820
rect 118555 580755 118621 580756
rect 161430 580685 161490 581163
rect 190502 581090 190562 581163
rect 191054 581090 191114 581435
rect 190502 581030 191114 581090
rect 195838 580957 195898 581571
rect 200990 581229 201050 582251
rect 202404 582000 203004 599498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 582000 206604 603098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 582000 210204 606698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 210371 582180 210437 582181
rect 210371 582116 210372 582180
rect 210436 582116 210437 582180
rect 210371 582115 210437 582116
rect 205587 581636 205653 581637
rect 205587 581572 205588 581636
rect 205652 581572 205653 581636
rect 205587 581571 205653 581572
rect 205590 581229 205650 581571
rect 200987 581228 201053 581229
rect 200987 581164 200988 581228
rect 201052 581164 201053 581228
rect 200987 581163 201053 581164
rect 205587 581228 205653 581229
rect 205587 581164 205588 581228
rect 205652 581164 205653 581228
rect 205587 581163 205653 581164
rect 210374 581093 210434 582115
rect 216804 582000 217404 613898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582000 221004 617498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 221227 582044 221293 582045
rect 221227 581980 221228 582044
rect 221292 581980 221293 582044
rect 224004 582000 224604 585098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 582000 228204 588698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 233923 584492 233989 584493
rect 233923 584428 233924 584492
rect 233988 584428 233989 584492
rect 233923 584427 233989 584428
rect 233926 583898 233986 584427
rect 229323 582044 229389 582045
rect 221227 581979 221293 581980
rect 229323 581980 229324 582044
rect 229388 581980 229389 582044
rect 234804 582000 235404 595898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 582000 239004 599498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 582000 242604 603098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 582000 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 249747 582044 249813 582045
rect 229323 581979 229389 581980
rect 249747 581980 249748 582044
rect 249812 581980 249813 582044
rect 252804 582000 253404 613898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582000 257004 617498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 582000 260604 585098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 260787 582180 260853 582181
rect 260787 582116 260788 582180
rect 260852 582116 260853 582180
rect 260787 582115 260853 582116
rect 249747 581979 249813 581980
rect 221230 581093 221290 581979
rect 224907 581636 224973 581637
rect 224907 581572 224908 581636
rect 224972 581572 224973 581636
rect 224907 581571 224973 581572
rect 224910 581229 224970 581571
rect 224907 581228 224973 581229
rect 224907 581164 224908 581228
rect 224972 581164 224973 581228
rect 224907 581163 224973 581164
rect 229326 581093 229386 581979
rect 249011 581908 249077 581909
rect 249011 581844 249012 581908
rect 249076 581844 249077 581908
rect 249011 581843 249077 581844
rect 244227 581636 244293 581637
rect 244227 581572 244228 581636
rect 244292 581572 244293 581636
rect 244227 581571 244293 581572
rect 231899 581364 231965 581365
rect 231899 581300 231900 581364
rect 231964 581300 231965 581364
rect 231899 581299 231965 581300
rect 210371 581092 210437 581093
rect 210371 581028 210372 581092
rect 210436 581028 210437 581092
rect 210371 581027 210437 581028
rect 221227 581092 221293 581093
rect 221227 581028 221228 581092
rect 221292 581028 221293 581092
rect 221227 581027 221293 581028
rect 229323 581092 229389 581093
rect 229323 581028 229324 581092
rect 229388 581028 229389 581092
rect 229323 581027 229389 581028
rect 179275 580956 179341 580957
rect 179275 580892 179276 580956
rect 179340 580892 179341 580956
rect 179275 580891 179341 580892
rect 195835 580956 195901 580957
rect 195835 580892 195836 580956
rect 195900 580892 195901 580956
rect 195835 580891 195901 580892
rect 161427 580684 161493 580685
rect 161427 580620 161428 580684
rect 161492 580620 161493 580684
rect 161427 580619 161493 580620
rect 169707 580684 169773 580685
rect 169707 580620 169708 580684
rect 169772 580620 169773 580684
rect 169707 580619 169773 580620
rect 113771 580548 113837 580549
rect 113771 580498 113772 580548
rect 113836 580498 113837 580548
rect 114507 580548 114573 580549
rect 114507 580498 114508 580548
rect 114572 580498 114573 580548
rect 123707 580548 123773 580549
rect 123707 580498 123708 580548
rect 123772 580498 123773 580548
rect 124259 580548 124325 580549
rect 124259 580498 124260 580548
rect 124324 580498 124325 580548
rect 137139 580548 137205 580549
rect 137139 580498 137140 580548
rect 137204 580498 137205 580548
rect 142107 580548 142173 580549
rect 142107 580498 142108 580548
rect 142172 580498 142173 580548
rect 151491 580548 151557 580549
rect 151491 580498 151492 580548
rect 151556 580498 151557 580548
rect 151859 580548 151925 580549
rect 151859 580498 151860 580548
rect 151924 580498 151925 580548
rect 161243 580548 161309 580549
rect 161243 580498 161244 580548
rect 161308 580498 161309 580548
rect 166211 580548 166277 580549
rect 166211 580498 166212 580548
rect 166276 580498 166277 580548
rect 167683 580548 167749 580549
rect 167683 580498 167684 580548
rect 167748 580498 167749 580548
rect 169710 580141 169770 580619
rect 179278 580141 179338 580891
rect 197307 580548 197373 580549
rect 197307 580498 197308 580548
rect 197372 580498 197373 580548
rect 206875 580548 206941 580549
rect 206875 580498 206876 580548
rect 206940 580498 206941 580548
rect 216627 580548 216693 580549
rect 216627 580498 216628 580548
rect 216692 580498 216693 580548
rect 226195 580548 226261 580549
rect 226195 580498 226196 580548
rect 226260 580498 226261 580548
rect 215306 580350 215806 580410
rect 227082 580350 227582 580410
rect 231902 580413 231962 581299
rect 244230 581229 244290 581571
rect 244227 581228 244293 581229
rect 244227 581164 244228 581228
rect 244292 581164 244293 581228
rect 244227 581163 244293 581164
rect 249014 581093 249074 581843
rect 249750 581229 249810 581979
rect 258947 581908 259013 581909
rect 258947 581844 258948 581908
rect 259012 581844 259013 581908
rect 258947 581843 259013 581844
rect 249747 581228 249813 581229
rect 249747 581164 249748 581228
rect 249812 581164 249813 581228
rect 249747 581163 249813 581164
rect 258950 581093 259010 581843
rect 260603 581636 260669 581637
rect 260603 581572 260604 581636
rect 260668 581572 260669 581636
rect 260603 581571 260669 581572
rect 260606 581229 260666 581571
rect 260790 581229 260850 582115
rect 263604 582000 264204 588698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 268515 582044 268581 582045
rect 268515 581980 268516 582044
rect 268580 581980 268581 582044
rect 270804 582000 271404 595898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 582000 275004 599498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 277531 582180 277597 582181
rect 277531 582116 277532 582180
rect 277596 582116 277597 582180
rect 277531 582115 277597 582116
rect 268515 581979 268581 581980
rect 268331 581908 268397 581909
rect 268331 581844 268332 581908
rect 268396 581844 268397 581908
rect 268331 581843 268397 581844
rect 260603 581228 260669 581229
rect 260603 581164 260604 581228
rect 260668 581164 260669 581228
rect 260603 581163 260669 581164
rect 260787 581228 260853 581229
rect 260787 581164 260788 581228
rect 260852 581164 260853 581228
rect 260787 581163 260853 581164
rect 268334 581093 268394 581843
rect 268518 581229 268578 581979
rect 277534 581229 277594 582115
rect 277715 582044 277781 582045
rect 277715 581980 277716 582044
rect 277780 581980 277781 582044
rect 278004 582000 278604 603098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 582000 282204 606698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 287835 582180 287901 582181
rect 287835 582116 287836 582180
rect 287900 582116 287901 582180
rect 287835 582115 287901 582116
rect 287651 582044 287717 582045
rect 277715 581979 277781 581980
rect 287651 581980 287652 582044
rect 287716 581980 287717 582044
rect 287651 581979 287717 581980
rect 268515 581228 268581 581229
rect 268515 581164 268516 581228
rect 268580 581164 268581 581228
rect 268515 581163 268581 581164
rect 277531 581228 277597 581229
rect 277531 581164 277532 581228
rect 277596 581164 277597 581228
rect 277531 581163 277597 581164
rect 277718 581093 277778 581979
rect 287654 581093 287714 581979
rect 287838 581229 287898 582115
rect 288804 582000 289404 613898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582000 293004 617498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 582000 296604 585098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 298142 583813 298202 584342
rect 298139 583812 298205 583813
rect 298139 583748 298140 583812
rect 298204 583748 298205 583812
rect 298139 583747 298205 583748
rect 297219 582180 297285 582181
rect 297219 582116 297220 582180
rect 297284 582116 297285 582180
rect 297219 582115 297285 582116
rect 297222 581229 297282 582115
rect 297403 582044 297469 582045
rect 297403 581980 297404 582044
rect 297468 581980 297469 582044
rect 299604 582000 300204 588698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306603 582180 306669 582181
rect 306603 582116 306604 582180
rect 306668 582116 306669 582180
rect 306603 582115 306669 582116
rect 306051 582044 306117 582045
rect 297403 581979 297469 581980
rect 306051 581980 306052 582044
rect 306116 581980 306117 582044
rect 306051 581979 306117 581980
rect 287835 581228 287901 581229
rect 287835 581164 287836 581228
rect 287900 581164 287901 581228
rect 287835 581163 287901 581164
rect 297219 581228 297285 581229
rect 297219 581164 297220 581228
rect 297284 581164 297285 581228
rect 297219 581163 297285 581164
rect 297406 581093 297466 581979
rect 306054 581093 306114 581979
rect 306606 581229 306666 582115
rect 306804 582000 307404 595898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 582000 311004 599498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 582000 314604 603098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 316539 582316 316605 582317
rect 316539 582252 316540 582316
rect 316604 582252 316605 582316
rect 316539 582251 316605 582252
rect 306603 581228 306669 581229
rect 306603 581164 306604 581228
rect 306668 581164 306669 581228
rect 306603 581163 306669 581164
rect 316542 581093 316602 582251
rect 316723 582180 316789 582181
rect 316723 582116 316724 582180
rect 316788 582116 316789 582180
rect 316723 582115 316789 582116
rect 316726 581229 316786 582115
rect 317604 582000 318204 606698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 582000 325404 613898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 326475 582316 326541 582317
rect 326475 582252 326476 582316
rect 326540 582252 326541 582316
rect 326475 582251 326541 582252
rect 326291 582180 326357 582181
rect 326291 582116 326292 582180
rect 326356 582116 326357 582180
rect 326291 582115 326357 582116
rect 321875 581636 321941 581637
rect 321875 581572 321876 581636
rect 321940 581572 321941 581636
rect 321875 581571 321941 581572
rect 316723 581228 316789 581229
rect 316723 581164 316724 581228
rect 316788 581164 316789 581228
rect 316723 581163 316789 581164
rect 249011 581092 249077 581093
rect 249011 581028 249012 581092
rect 249076 581028 249077 581092
rect 249011 581027 249077 581028
rect 258947 581092 259013 581093
rect 258947 581028 258948 581092
rect 259012 581028 259013 581092
rect 258947 581027 259013 581028
rect 268331 581092 268397 581093
rect 268331 581028 268332 581092
rect 268396 581028 268397 581092
rect 268331 581027 268397 581028
rect 277715 581092 277781 581093
rect 277715 581028 277716 581092
rect 277780 581028 277781 581092
rect 277715 581027 277781 581028
rect 287651 581092 287717 581093
rect 287651 581028 287652 581092
rect 287716 581028 287717 581092
rect 287651 581027 287717 581028
rect 297403 581092 297469 581093
rect 297403 581028 297404 581092
rect 297468 581028 297469 581092
rect 297403 581027 297469 581028
rect 306051 581092 306117 581093
rect 306051 581028 306052 581092
rect 306116 581028 306117 581092
rect 306051 581027 306117 581028
rect 316539 581092 316605 581093
rect 316539 581028 316540 581092
rect 316604 581028 316605 581092
rect 316539 581027 316605 581028
rect 231899 580412 231965 580413
rect 231899 580348 231900 580412
rect 231964 580348 231965 580412
rect 231899 580347 231965 580348
rect 311906 580350 312406 580410
rect 169707 580140 169773 580141
rect 169707 580076 169708 580140
rect 169772 580076 169773 580140
rect 169707 580075 169773 580076
rect 179275 580140 179341 580141
rect 179275 580076 179276 580140
rect 179340 580076 179341 580140
rect 321878 580277 321938 581571
rect 326294 581229 326354 582115
rect 326291 581228 326357 581229
rect 326291 581164 326292 581228
rect 326356 581164 326357 581228
rect 326291 581163 326357 581164
rect 326478 581093 326538 582251
rect 328404 582000 329004 617498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 582000 332604 585098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 582000 336204 588698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 582000 343404 595898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 582000 347004 599498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 582000 350604 603098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 582000 354204 606698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 582000 361404 613898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582000 365004 617498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 582000 368604 585098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 582000 372204 588698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 582000 379404 595898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 582000 383004 599498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 582000 386604 603098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 582000 390204 606698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 393451 582180 393517 582181
rect 393451 582116 393452 582180
rect 393516 582116 393517 582180
rect 393451 582115 393517 582116
rect 335859 581772 335925 581773
rect 335859 581708 335860 581772
rect 335924 581708 335925 581772
rect 335859 581707 335925 581708
rect 350395 581772 350461 581773
rect 350395 581708 350396 581772
rect 350460 581708 350461 581772
rect 350395 581707 350461 581708
rect 355363 581772 355429 581773
rect 355363 581708 355364 581772
rect 355428 581708 355429 581772
rect 355363 581707 355429 581708
rect 364747 581772 364813 581773
rect 364747 581708 364748 581772
rect 364812 581708 364813 581772
rect 364747 581707 364813 581708
rect 374131 581772 374197 581773
rect 374131 581708 374132 581772
rect 374196 581708 374197 581772
rect 374131 581707 374197 581708
rect 384435 581772 384501 581773
rect 384435 581708 384436 581772
rect 384500 581708 384501 581772
rect 384435 581707 384501 581708
rect 393267 581772 393333 581773
rect 393267 581708 393268 581772
rect 393332 581708 393333 581772
rect 393267 581707 393333 581708
rect 335862 581229 335922 581707
rect 336043 581636 336109 581637
rect 336043 581572 336044 581636
rect 336108 581572 336109 581636
rect 336043 581571 336109 581572
rect 345611 581636 345677 581637
rect 345611 581572 345612 581636
rect 345676 581572 345677 581636
rect 345611 581571 345677 581572
rect 346899 581636 346965 581637
rect 346899 581572 346900 581636
rect 346964 581572 346965 581636
rect 346899 581571 346965 581572
rect 335859 581228 335925 581229
rect 335859 581164 335860 581228
rect 335924 581164 335925 581228
rect 335859 581163 335925 581164
rect 336046 581093 336106 581571
rect 345614 581093 345674 581571
rect 326475 581092 326541 581093
rect 326475 581028 326476 581092
rect 326540 581028 326541 581092
rect 326475 581027 326541 581028
rect 336043 581092 336109 581093
rect 336043 581028 336044 581092
rect 336108 581028 336109 581092
rect 336043 581027 336109 581028
rect 345611 581092 345677 581093
rect 345611 581028 345612 581092
rect 345676 581028 345677 581092
rect 345611 581027 345677 581028
rect 321875 580276 321941 580277
rect 321875 580212 321876 580276
rect 321940 580212 321941 580276
rect 346902 580413 346962 581571
rect 350398 581229 350458 581707
rect 351683 581636 351749 581637
rect 351683 581572 351684 581636
rect 351748 581572 351749 581636
rect 351683 581571 351749 581572
rect 355179 581636 355245 581637
rect 355179 581572 355180 581636
rect 355244 581572 355245 581636
rect 355179 581571 355245 581572
rect 350395 581228 350461 581229
rect 350395 581164 350396 581228
rect 350460 581164 350461 581228
rect 350395 581163 350461 581164
rect 346899 580412 346965 580413
rect 346899 580348 346900 580412
rect 346964 580348 346965 580412
rect 346899 580347 346965 580348
rect 351686 580277 351746 581571
rect 355182 581229 355242 581571
rect 355179 581228 355245 581229
rect 355179 581164 355180 581228
rect 355244 581164 355245 581228
rect 355179 581163 355245 581164
rect 355366 581093 355426 581707
rect 360147 581636 360213 581637
rect 360147 581572 360148 581636
rect 360212 581572 360213 581636
rect 360147 581571 360213 581572
rect 358675 581364 358741 581365
rect 358675 581300 358676 581364
rect 358740 581300 358741 581364
rect 358675 581299 358741 581300
rect 355363 581092 355429 581093
rect 355363 581028 355364 581092
rect 355428 581028 355429 581092
rect 355363 581027 355429 581028
rect 358678 580549 358738 581299
rect 360150 581229 360210 581571
rect 360147 581228 360213 581229
rect 360147 581164 360148 581228
rect 360212 581164 360213 581228
rect 360147 581163 360213 581164
rect 364750 581093 364810 581707
rect 365115 581636 365181 581637
rect 365115 581572 365116 581636
rect 365180 581572 365181 581636
rect 365115 581571 365181 581572
rect 373947 581636 374013 581637
rect 373947 581572 373948 581636
rect 374012 581572 374013 581636
rect 373947 581571 374013 581572
rect 364747 581092 364813 581093
rect 364747 581028 364748 581092
rect 364812 581028 364813 581092
rect 364747 581027 364813 581028
rect 358675 580548 358741 580549
rect 358675 580484 358676 580548
rect 358740 580484 358741 580548
rect 365118 580498 365178 581571
rect 373950 581093 374010 581571
rect 374134 581229 374194 581707
rect 384251 581636 384317 581637
rect 384251 581572 384252 581636
rect 384316 581572 384317 581636
rect 384251 581571 384317 581572
rect 374131 581228 374197 581229
rect 374131 581164 374132 581228
rect 374196 581164 374197 581228
rect 374131 581163 374197 581164
rect 384254 581093 384314 581571
rect 384438 581229 384498 581707
rect 384803 581636 384869 581637
rect 384803 581572 384804 581636
rect 384868 581572 384869 581636
rect 384803 581571 384869 581572
rect 389771 581636 389837 581637
rect 389771 581572 389772 581636
rect 389836 581572 389837 581636
rect 389771 581571 389837 581572
rect 391795 581636 391861 581637
rect 391795 581572 391796 581636
rect 391860 581572 391861 581636
rect 391795 581571 391861 581572
rect 384435 581228 384501 581229
rect 384435 581164 384436 581228
rect 384500 581164 384501 581228
rect 384435 581163 384501 581164
rect 373947 581092 374013 581093
rect 373947 581028 373948 581092
rect 374012 581028 374013 581092
rect 373947 581027 374013 581028
rect 384251 581092 384317 581093
rect 384251 581028 384252 581092
rect 384316 581028 384317 581092
rect 384251 581027 384317 581028
rect 384806 580821 384866 581571
rect 389774 580957 389834 581571
rect 389771 580956 389837 580957
rect 389771 580892 389772 580956
rect 389836 580892 389837 580956
rect 389771 580891 389837 580892
rect 384803 580820 384869 580821
rect 384803 580756 384804 580820
rect 384868 580756 384869 580820
rect 384803 580755 384869 580756
rect 391798 580685 391858 581571
rect 393270 581093 393330 581707
rect 393454 581229 393514 582115
rect 396804 582000 397404 613898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582000 401004 617498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 403755 582180 403821 582181
rect 403755 582116 403756 582180
rect 403820 582116 403821 582180
rect 403755 582115 403821 582116
rect 403571 581772 403637 581773
rect 403571 581708 403572 581772
rect 403636 581708 403637 581772
rect 403571 581707 403637 581708
rect 393451 581228 393517 581229
rect 393451 581164 393452 581228
rect 393516 581164 393517 581228
rect 393451 581163 393517 581164
rect 403574 581093 403634 581707
rect 403758 581229 403818 582115
rect 404004 582000 404604 585098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 582000 408204 588698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 412771 582316 412837 582317
rect 412771 582252 412772 582316
rect 412836 582252 412837 582316
rect 412771 582251 412837 582252
rect 412587 582180 412653 582181
rect 412587 582116 412588 582180
rect 412652 582116 412653 582180
rect 412587 582115 412653 582116
rect 403755 581228 403821 581229
rect 403755 581164 403756 581228
rect 403820 581164 403821 581228
rect 403755 581163 403821 581164
rect 412590 581093 412650 582115
rect 412774 581229 412834 582251
rect 414804 582000 415404 595898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 582000 419004 599498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 582000 422604 603098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 423075 582316 423141 582317
rect 423075 582252 423076 582316
rect 423140 582252 423141 582316
rect 423075 582251 423141 582252
rect 422891 582180 422957 582181
rect 422891 582116 422892 582180
rect 422956 582116 422957 582180
rect 422891 582115 422957 582116
rect 412771 581228 412837 581229
rect 412771 581164 412772 581228
rect 412836 581164 412837 581228
rect 412771 581163 412837 581164
rect 422894 581093 422954 582115
rect 423078 581229 423138 582251
rect 425604 582000 426204 606698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 431907 582316 431973 582317
rect 431907 582252 431908 582316
rect 431972 582252 431973 582316
rect 431907 582251 431973 582252
rect 423075 581228 423141 581229
rect 423075 581164 423076 581228
rect 423140 581164 423141 581228
rect 423075 581163 423141 581164
rect 431910 581093 431970 582251
rect 432804 582000 433404 613898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582000 437004 617498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 582000 440604 585098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 442211 582316 442277 582317
rect 442211 582252 442212 582316
rect 442276 582252 442277 582316
rect 442211 582251 442277 582252
rect 432091 581228 432157 581229
rect 432091 581164 432092 581228
rect 432156 581164 432157 581228
rect 432091 581163 432157 581164
rect 437427 581228 437493 581229
rect 437427 581164 437428 581228
rect 437492 581164 437493 581228
rect 437427 581163 437493 581164
rect 393267 581092 393333 581093
rect 393267 581028 393268 581092
rect 393332 581028 393333 581092
rect 393267 581027 393333 581028
rect 403571 581092 403637 581093
rect 403571 581028 403572 581092
rect 403636 581028 403637 581092
rect 403571 581027 403637 581028
rect 412587 581092 412653 581093
rect 412587 581028 412588 581092
rect 412652 581028 412653 581092
rect 412587 581027 412653 581028
rect 422891 581092 422957 581093
rect 422891 581028 422892 581092
rect 422956 581028 422957 581092
rect 422891 581027 422957 581028
rect 431907 581092 431973 581093
rect 431907 581028 431908 581092
rect 431972 581028 431973 581092
rect 431907 581027 431973 581028
rect 391795 580684 391861 580685
rect 391795 580620 391796 580684
rect 391860 580620 391861 580684
rect 391795 580619 391861 580620
rect 358675 580483 358741 580484
rect 351683 580276 351749 580277
rect 321875 580211 321941 580212
rect 328318 580141 328378 580262
rect 351683 580212 351684 580276
rect 351748 580212 351749 580276
rect 351683 580211 351749 580212
rect 432094 580141 432154 581163
rect 437430 580141 437490 581163
rect 442214 581093 442274 582251
rect 443604 582000 444204 588698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 582000 451404 595898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 451963 582316 452029 582317
rect 451963 582252 451964 582316
rect 452028 582252 452029 582316
rect 451963 582251 452029 582252
rect 451966 581093 452026 582251
rect 454404 582000 455004 599498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 582000 458604 603098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461347 582316 461413 582317
rect 461347 582252 461348 582316
rect 461412 582252 461413 582316
rect 461347 582251 461413 582252
rect 456563 581228 456629 581229
rect 456563 581164 456564 581228
rect 456628 581164 456629 581228
rect 456563 581163 456629 581164
rect 456747 581228 456813 581229
rect 456747 581164 456748 581228
rect 456812 581164 456813 581228
rect 456747 581163 456813 581164
rect 442211 581092 442277 581093
rect 442211 581028 442212 581092
rect 442276 581028 442277 581092
rect 442211 581027 442277 581028
rect 451963 581092 452029 581093
rect 451963 581028 451964 581092
rect 452028 581028 452029 581092
rect 451963 581027 452029 581028
rect 456566 580141 456626 581163
rect 456750 580141 456810 581163
rect 461350 581093 461410 582251
rect 461604 582000 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 582000 469404 613898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 470547 582316 470613 582317
rect 470547 582252 470548 582316
rect 470612 582252 470613 582316
rect 470547 582251 470613 582252
rect 470550 581093 470610 582251
rect 472404 582000 473004 617498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 582000 476604 585098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 582000 480204 588698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 480851 582316 480917 582317
rect 480851 582252 480852 582316
rect 480916 582252 480917 582316
rect 480851 582251 480917 582252
rect 470731 581228 470797 581229
rect 470731 581164 470732 581228
rect 470796 581164 470797 581228
rect 470731 581163 470797 581164
rect 476067 581228 476133 581229
rect 476067 581164 476068 581228
rect 476132 581164 476133 581228
rect 476067 581163 476133 581164
rect 461347 581092 461413 581093
rect 461347 581028 461348 581092
rect 461412 581028 461413 581092
rect 461347 581027 461413 581028
rect 470547 581092 470613 581093
rect 470547 581028 470548 581092
rect 470612 581028 470613 581092
rect 470547 581027 470613 581028
rect 470734 580141 470794 581163
rect 476070 580141 476130 581163
rect 480854 581093 480914 582251
rect 486804 582000 487404 595898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 489867 582316 489933 582317
rect 489867 582252 489868 582316
rect 489932 582252 489933 582316
rect 489867 582251 489933 582252
rect 489870 581229 489930 582251
rect 490404 582000 491004 599498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 491707 582180 491773 582181
rect 491707 582116 491708 582180
rect 491772 582116 491773 582180
rect 491707 582115 491773 582116
rect 489867 581228 489933 581229
rect 489867 581164 489868 581228
rect 489932 581164 489933 581228
rect 489867 581163 489933 581164
rect 480851 581092 480917 581093
rect 480851 581028 480852 581092
rect 480916 581028 480917 581092
rect 480851 581027 480917 581028
rect 489867 581092 489933 581093
rect 489867 581028 489868 581092
rect 489932 581028 489933 581092
rect 489867 581027 489933 581028
rect 328315 580140 328381 580141
rect 179275 580075 179341 580076
rect 318747 580076 318748 580126
rect 318812 580076 318813 580126
rect 318747 580075 318813 580076
rect 328315 580076 328316 580140
rect 328380 580076 328381 580140
rect 328315 580075 328381 580076
rect 432091 580140 432157 580141
rect 432091 580076 432092 580140
rect 432156 580076 432157 580140
rect 432091 580075 432157 580076
rect 437427 580140 437493 580141
rect 437427 580076 437428 580140
rect 437492 580076 437493 580140
rect 437427 580075 437493 580076
rect 456563 580140 456629 580141
rect 456563 580076 456564 580140
rect 456628 580076 456629 580140
rect 456563 580075 456629 580076
rect 456747 580140 456813 580141
rect 456747 580076 456748 580140
rect 456812 580076 456813 580140
rect 456747 580075 456813 580076
rect 470731 580140 470797 580141
rect 470731 580076 470732 580140
rect 470796 580076 470797 580140
rect 470731 580075 470797 580076
rect 476067 580140 476133 580141
rect 476067 580076 476068 580140
rect 476132 580076 476133 580140
rect 476067 580075 476133 580076
rect 489870 580005 489930 581027
rect 491710 580141 491770 582115
rect 494004 582000 494604 603098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497411 582044 497477 582045
rect 497411 581980 497412 582044
rect 497476 581980 497477 582044
rect 497604 582000 498204 606698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 505691 696964 505757 696965
rect 505691 696900 505692 696964
rect 505756 696900 505757 696964
rect 505691 696899 505757 696900
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 501643 584900 501709 584901
rect 501643 584836 501644 584900
rect 501708 584836 501709 584900
rect 501643 584835 501709 584836
rect 499435 583948 499501 583949
rect 499435 583898 499436 583948
rect 499500 583898 499501 583948
rect 499067 583812 499133 583813
rect 499067 583748 499068 583812
rect 499132 583748 499133 583812
rect 499067 583747 499133 583748
rect 497411 581979 497477 581980
rect 497414 581770 497474 581979
rect 498147 581908 498213 581909
rect 498147 581844 498148 581908
rect 498212 581844 498213 581908
rect 498147 581843 498213 581844
rect 497414 581710 497658 581770
rect 495387 581228 495453 581229
rect 495387 581164 495388 581228
rect 495452 581164 495453 581228
rect 495387 581163 495453 581164
rect 491707 580140 491773 580141
rect 491707 580076 491708 580140
rect 491772 580076 491773 580140
rect 491707 580075 491773 580076
rect 495390 580005 495450 581163
rect 489867 580004 489933 580005
rect 489867 579940 489868 580004
rect 489932 579940 489933 580004
rect 489867 579939 489933 579940
rect 495387 580004 495453 580005
rect 495387 579940 495388 580004
rect 495452 579940 495453 580004
rect 495387 579939 495453 579940
rect 97763 579868 97829 579869
rect 97763 579804 97764 579868
rect 97828 579804 97829 579868
rect 97763 579803 97829 579804
rect 101814 576418 101874 578902
rect 101814 571570 101874 573462
rect 101630 571510 101874 571570
rect 101630 541058 101690 571510
rect 497598 540970 497658 581710
rect 497598 540910 497842 540970
rect 101814 521930 101874 535382
rect 497782 531450 497842 540910
rect 101630 521870 101874 521930
rect 497598 531390 497842 531450
rect 101630 521338 101690 521870
rect 101630 517850 101690 519742
rect 101630 517790 101874 517850
rect 101814 487338 101874 517790
rect 101726 487298 101962 487338
rect 101726 487022 101962 487062
rect 101814 483850 101874 487022
rect 101630 483790 101874 483850
rect 101630 471610 101690 483790
rect 101630 471550 101874 471610
rect 101814 458778 101874 471550
rect 101627 456452 101628 456502
rect 101692 456452 101693 456502
rect 101627 456451 101693 456452
rect 101630 446450 101690 446982
rect 101630 446390 101874 446450
rect 101814 445090 101874 446390
rect 101630 445030 101874 445090
rect 101630 414490 101690 445030
rect 101630 414430 101874 414490
rect 101814 402930 101874 414430
rect 497598 409050 497658 531390
rect 497598 408990 497842 409050
rect 101630 402870 101874 402930
rect 101630 394770 101690 402870
rect 497782 396130 497842 408990
rect 497598 396070 497842 396130
rect 101630 394710 101726 394770
rect 101778 392670 101874 392730
rect 101814 378450 101874 392670
rect 101778 378390 101874 378450
rect 101778 376350 101874 376410
rect 101814 374370 101874 376350
rect 101630 374310 101874 374370
rect 101630 327450 101690 374310
rect 101630 327390 101874 327450
rect 101814 324730 101874 327390
rect 101778 324670 101874 324730
rect 101630 322630 101726 322690
rect 101630 318610 101690 322630
rect 101630 318550 101874 318610
rect 101814 307050 101874 318550
rect 101630 306990 101874 307050
rect 101630 305778 101690 306990
rect 101814 302290 101874 303502
rect 101630 302230 101874 302290
rect 101630 281890 101690 302230
rect 497598 291410 497658 396070
rect 498150 390690 498210 581843
rect 498331 581772 498397 581773
rect 498331 581708 498332 581772
rect 498396 581708 498397 581772
rect 498331 581707 498397 581708
rect 497782 390630 498210 390690
rect 497782 293450 497842 390630
rect 498334 390010 498394 581707
rect 498699 581636 498765 581637
rect 498699 581572 498700 581636
rect 498764 581572 498765 581636
rect 498699 581571 498765 581572
rect 498702 573746 498762 581571
rect 498702 573686 498946 573746
rect 498886 572250 498946 573686
rect 498702 572190 498946 572250
rect 499070 572250 499130 583747
rect 500355 582996 500421 582997
rect 500355 582932 500356 582996
rect 500420 582932 500421 582996
rect 500355 582931 500421 582932
rect 499987 581636 500053 581637
rect 499987 581572 499988 581636
rect 500052 581572 500053 581636
rect 499987 581571 500053 581572
rect 499990 581229 500050 581571
rect 499987 581228 500053 581229
rect 499987 581164 499988 581228
rect 500052 581164 500053 581228
rect 499987 581163 500053 581164
rect 499070 572190 499314 572250
rect 498702 568938 498762 572190
rect 499254 568170 499314 572190
rect 499070 568110 499314 568170
rect 499070 418298 499130 568110
rect 499622 545050 499682 568702
rect 499438 544990 499682 545050
rect 499438 536890 499498 544990
rect 499438 536830 499682 536890
rect 499622 535530 499682 536830
rect 499438 535470 499682 535530
rect 499438 527370 499498 535470
rect 499254 527310 499498 527370
rect 499254 517850 499314 527310
rect 500358 522610 500418 582931
rect 501275 582724 501341 582725
rect 501275 582660 501276 582724
rect 501340 582660 501341 582724
rect 501275 582659 501341 582660
rect 501091 580820 501157 580821
rect 501091 580756 501092 580820
rect 501156 580756 501157 580820
rect 501091 580755 501157 580756
rect 501094 573610 501154 580755
rect 501278 573749 501338 582659
rect 501275 573748 501341 573749
rect 501275 573684 501276 573748
rect 501340 573684 501341 573748
rect 501275 573683 501341 573684
rect 501275 573612 501341 573613
rect 501275 573610 501276 573612
rect 501094 573550 501276 573610
rect 501275 573548 501276 573550
rect 501340 573548 501341 573612
rect 501275 573547 501341 573548
rect 501459 572252 501525 572253
rect 501459 572250 501460 572252
rect 500174 522550 500418 522610
rect 501278 572190 501460 572250
rect 499254 517790 499682 517850
rect 499622 500850 499682 517790
rect 500174 512410 500234 522550
rect 501278 517309 501338 572190
rect 501459 572188 501460 572190
rect 501524 572188 501525 572252
rect 501459 572187 501525 572188
rect 501459 571980 501525 571981
rect 501459 571916 501460 571980
rect 501524 571916 501525 571980
rect 501459 571915 501525 571916
rect 501462 557157 501522 571915
rect 501459 557156 501525 557157
rect 501459 557092 501460 557156
rect 501524 557092 501525 557156
rect 501459 557091 501525 557092
rect 501459 547908 501525 547909
rect 501459 547844 501460 547908
rect 501524 547844 501525 547908
rect 501459 547843 501525 547844
rect 501275 517308 501341 517309
rect 501275 517244 501276 517308
rect 501340 517244 501341 517308
rect 501275 517243 501341 517244
rect 501275 513772 501341 513773
rect 501275 513708 501276 513772
rect 501340 513708 501341 513772
rect 501275 513707 501341 513708
rect 500174 512350 500418 512410
rect 500358 504930 500418 512350
rect 501278 512005 501338 513707
rect 501275 512004 501341 512005
rect 501275 511940 501276 512004
rect 501340 511940 501341 512004
rect 501275 511939 501341 511940
rect 501462 511730 501522 547843
rect 501646 520165 501706 584835
rect 502011 580548 502077 580549
rect 502011 580484 502012 580548
rect 502076 580484 502077 580548
rect 502011 580483 502077 580484
rect 501827 573612 501893 573613
rect 501827 573548 501828 573612
rect 501892 573548 501893 573612
rect 501827 573547 501893 573548
rect 501830 571981 501890 573547
rect 501827 571980 501893 571981
rect 501827 571916 501828 571980
rect 501892 571916 501893 571980
rect 501827 571915 501893 571916
rect 502014 559058 502074 580483
rect 501830 558998 502074 559058
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 501643 520164 501709 520165
rect 501643 520100 501644 520164
rect 501708 520100 501709 520164
rect 501643 520099 501709 520100
rect 501643 519620 501709 519621
rect 501643 519556 501644 519620
rect 501708 519556 501709 519620
rect 501643 519555 501709 519556
rect 501646 512410 501706 519555
rect 501830 517306 501890 558998
rect 504804 542454 505404 577898
rect 505507 570076 505573 570077
rect 505507 570012 505508 570076
rect 505572 570012 505573 570076
rect 505507 570011 505573 570012
rect 502563 542332 502629 542333
rect 502563 542268 502564 542332
rect 502628 542268 502629 542332
rect 502563 542267 502629 542268
rect 502011 517308 502077 517309
rect 502011 517306 502012 517308
rect 501830 517246 502012 517306
rect 502011 517244 502012 517246
rect 502076 517244 502077 517308
rect 502011 517243 502077 517244
rect 502195 517308 502261 517309
rect 502195 517244 502196 517308
rect 502260 517244 502261 517308
rect 502195 517243 502261 517244
rect 501646 512350 501890 512410
rect 500726 511670 501522 511730
rect 500726 507738 500786 511670
rect 501275 506972 501341 506973
rect 501275 506908 501276 506972
rect 501340 506908 501341 506972
rect 501275 506907 501341 506908
rect 500358 504870 500602 504930
rect 499622 500790 500050 500850
rect 499990 499490 500050 500790
rect 499806 499430 500050 499490
rect 499806 491330 499866 499430
rect 500542 492010 500602 504870
rect 499622 491270 499866 491330
rect 499990 491950 500602 492010
rect 499622 474330 499682 491270
rect 499990 488610 500050 491950
rect 499990 488550 500418 488610
rect 500358 475010 500418 488550
rect 499254 474270 499682 474330
rect 499806 474950 500418 475010
rect 499254 458690 499314 474270
rect 499806 469570 499866 474950
rect 500910 473650 500970 500022
rect 501278 474877 501338 506907
rect 501275 474876 501341 474877
rect 501275 474812 501276 474876
rect 501340 474812 501341 474876
rect 501275 474811 501341 474812
rect 500174 473590 500970 473650
rect 500174 473058 500234 473590
rect 499622 469510 499866 469570
rect 499622 463450 499682 469510
rect 501094 467530 501154 472822
rect 501094 467470 501338 467530
rect 499622 463390 499866 463450
rect 499806 462770 499866 463390
rect 499806 462710 500050 462770
rect 499254 458630 499866 458690
rect 499806 441690 499866 458630
rect 499990 449850 500050 462710
rect 501278 456650 501338 467470
rect 501462 464541 501522 507502
rect 501830 506970 501890 512350
rect 502011 512004 502077 512005
rect 502011 511940 502012 512004
rect 502076 511940 502077 512004
rect 502011 511939 502077 511940
rect 501646 506910 501890 506970
rect 501459 464540 501525 464541
rect 501459 464476 501460 464540
rect 501524 464476 501525 464540
rect 501459 464475 501525 464476
rect 501646 464405 501706 506910
rect 501827 506836 501893 506837
rect 501827 506772 501828 506836
rect 501892 506772 501893 506836
rect 501827 506771 501893 506772
rect 501830 500853 501890 506771
rect 501827 500852 501893 500853
rect 501827 500788 501828 500852
rect 501892 500788 501893 500852
rect 501827 500787 501893 500788
rect 502014 500258 502074 511939
rect 502198 506837 502258 517243
rect 502195 506836 502261 506837
rect 502195 506772 502196 506836
rect 502260 506772 502261 506836
rect 502195 506771 502261 506772
rect 502379 503708 502445 503709
rect 502379 503644 502380 503708
rect 502444 503644 502445 503708
rect 502379 503643 502445 503644
rect 501827 493372 501893 493373
rect 501827 493308 501828 493372
rect 501892 493308 501893 493372
rect 501827 493307 501893 493308
rect 501830 478685 501890 493307
rect 501827 478684 501893 478685
rect 501827 478620 501828 478684
rect 501892 478620 501893 478684
rect 501827 478619 501893 478620
rect 502011 478684 502077 478685
rect 502011 478620 502012 478684
rect 502076 478620 502077 478684
rect 502011 478619 502077 478620
rect 501643 464404 501709 464405
rect 501643 464340 501644 464404
rect 501708 464340 501709 464404
rect 501643 464339 501709 464340
rect 501459 464268 501525 464269
rect 501459 464204 501460 464268
rect 501524 464204 501525 464268
rect 501459 464203 501525 464204
rect 500910 456590 501338 456650
rect 499990 449790 500234 449850
rect 499622 441630 499866 441690
rect 499622 439650 499682 441630
rect 499438 439590 499682 439650
rect 499438 432850 499498 439590
rect 500174 436930 500234 449790
rect 500174 436870 500418 436930
rect 499438 432790 499682 432850
rect 499622 427954 499682 432790
rect 499622 427894 499866 427954
rect 499070 418238 499314 418298
rect 499254 417210 499314 418238
rect 499806 417298 499866 427894
rect 500358 423874 500418 436870
rect 500358 423814 500602 423874
rect 499070 417150 499314 417210
rect 498702 411858 498762 417062
rect 499070 407010 499130 417150
rect 500542 413898 500602 423814
rect 499990 408506 500050 411622
rect 499438 408446 500050 408506
rect 499070 406950 499314 407010
rect 499254 405650 499314 406950
rect 499070 405590 499314 405650
rect 499070 390690 499130 405590
rect 499438 403746 499498 408446
rect 500358 407690 500418 412302
rect 500910 408370 500970 456590
rect 501462 454610 501522 464203
rect 501643 454884 501709 454885
rect 501643 454820 501644 454884
rect 501708 454820 501709 454884
rect 501643 454819 501709 454820
rect 501278 454550 501522 454610
rect 501278 442509 501338 454550
rect 501459 443324 501525 443325
rect 501459 443260 501460 443324
rect 501524 443260 501525 443324
rect 501459 443259 501525 443260
rect 501462 442509 501522 443259
rect 501275 442508 501341 442509
rect 501275 442444 501276 442508
rect 501340 442444 501341 442508
rect 501275 442443 501341 442444
rect 501459 442508 501525 442509
rect 501459 442444 501460 442508
rect 501524 442444 501525 442508
rect 501459 442443 501525 442444
rect 501459 442236 501525 442237
rect 501459 442172 501460 442236
rect 501524 442172 501525 442236
rect 501459 442171 501525 442172
rect 501275 439788 501341 439789
rect 501275 439724 501276 439788
rect 501340 439724 501341 439788
rect 501275 439723 501341 439724
rect 501278 438970 501338 439723
rect 499990 407630 500418 407690
rect 500726 408310 500970 408370
rect 501094 438910 501338 438970
rect 499438 403686 499866 403746
rect 499070 390630 499498 390690
rect 497966 389950 498394 390010
rect 497966 379130 498026 389950
rect 498518 385250 498578 388502
rect 499438 387970 499498 390630
rect 498334 385190 498578 385250
rect 499070 387910 499498 387970
rect 498334 383890 498394 385190
rect 498334 383830 498762 383890
rect 498702 383210 498762 383830
rect 498150 383150 498762 383210
rect 498150 381850 498210 383150
rect 498150 381790 498394 381850
rect 498334 379810 498394 381790
rect 498334 379750 498578 379810
rect 497966 379070 498394 379130
rect 498334 370970 498394 379070
rect 498150 370910 498394 370970
rect 498150 366978 498210 370910
rect 498518 366210 498578 379750
rect 498150 366150 498578 366210
rect 498150 360858 498210 366150
rect 498702 365530 498762 381022
rect 499070 377770 499130 387910
rect 499806 386610 499866 403686
rect 499990 398850 500050 407630
rect 499990 398790 500602 398850
rect 500542 395450 500602 398790
rect 500174 395390 500602 395450
rect 500174 387970 500234 395390
rect 500726 394770 500786 408310
rect 500542 394710 500786 394770
rect 500542 387970 500602 394710
rect 500174 387910 500418 387970
rect 500542 387910 500970 387970
rect 500358 386610 500418 387910
rect 499806 386550 500234 386610
rect 500358 386550 500602 386610
rect 499438 382618 499498 386462
rect 500174 385930 500234 386550
rect 500174 385870 500418 385930
rect 499990 381170 500050 385102
rect 499806 381110 500050 381170
rect 499438 380490 499498 381022
rect 499806 380490 499866 381110
rect 499438 380430 499866 380490
rect 500358 379810 500418 385870
rect 499622 379750 500418 379810
rect 499070 377710 499498 377770
rect 499438 376410 499498 377710
rect 499070 376350 499498 376410
rect 498702 365470 498946 365530
rect 498518 360090 498578 364702
rect 498886 364170 498946 365470
rect 498150 360030 498578 360090
rect 498702 364110 498946 364170
rect 498150 355330 498210 360030
rect 498702 358818 498762 364110
rect 499070 358594 499130 376350
rect 499622 367570 499682 379750
rect 500542 379130 500602 386550
rect 499438 367510 499682 367570
rect 500358 379070 500602 379130
rect 499438 366210 499498 367510
rect 499438 366150 499682 366210
rect 499070 358534 499498 358594
rect 499438 357370 499498 358534
rect 498702 357310 499498 357370
rect 498150 355270 498394 355330
rect 498334 311130 498394 355270
rect 498702 346354 498762 357310
rect 499254 355738 499314 356542
rect 499254 355678 499498 355738
rect 499438 354650 499498 355678
rect 499070 354590 499498 354650
rect 499070 354058 499130 354590
rect 499622 353970 499682 366150
rect 499990 364938 500050 366742
rect 500358 363490 500418 379070
rect 500174 363430 500418 363490
rect 500174 362810 500234 363430
rect 499438 353910 499682 353970
rect 499990 362750 500234 362810
rect 499438 353290 499498 353910
rect 499254 353230 499498 353290
rect 499254 349618 499314 353230
rect 499622 349978 499682 352462
rect 499990 349890 500050 362750
rect 500910 358050 500970 387910
rect 500174 357990 500970 358050
rect 500174 355330 500234 357990
rect 500174 355270 500418 355330
rect 500358 350658 500418 355270
rect 500726 349890 500786 357222
rect 501094 350570 501154 438910
rect 501462 438290 501522 442171
rect 501278 438230 501522 438290
rect 501278 427821 501338 438230
rect 501459 438156 501525 438157
rect 501459 438092 501460 438156
rect 501524 438092 501525 438156
rect 501459 438091 501525 438092
rect 501275 427820 501341 427821
rect 501275 427756 501276 427820
rect 501340 427756 501341 427820
rect 501275 427755 501341 427756
rect 501275 418300 501341 418301
rect 501275 418236 501276 418300
rect 501340 418236 501341 418300
rect 501275 418235 501341 418236
rect 501278 411501 501338 418235
rect 501275 411500 501341 411501
rect 501275 411436 501276 411500
rect 501340 411436 501341 411500
rect 501275 411435 501341 411436
rect 501275 410004 501341 410005
rect 501275 409940 501276 410004
rect 501340 409940 501341 410004
rect 501275 409939 501341 409940
rect 501278 351661 501338 409939
rect 501462 403749 501522 438091
rect 501646 408506 501706 454819
rect 502014 454749 502074 478619
rect 502195 464540 502261 464541
rect 502195 464476 502196 464540
rect 502260 464476 502261 464540
rect 502195 464475 502261 464476
rect 502011 454748 502077 454749
rect 502011 454684 502012 454748
rect 502076 454684 502077 454748
rect 502011 454683 502077 454684
rect 502198 449170 502258 464475
rect 502014 449110 502258 449170
rect 502014 438157 502074 449110
rect 502195 449036 502261 449037
rect 502195 448972 502196 449036
rect 502260 448972 502261 449036
rect 502195 448971 502261 448972
rect 502011 438156 502077 438157
rect 502011 438092 502012 438156
rect 502076 438092 502077 438156
rect 502011 438091 502077 438092
rect 502198 427954 502258 448971
rect 502014 427894 502258 427954
rect 502014 423877 502074 427894
rect 502011 423876 502077 423877
rect 502011 423812 502012 423876
rect 502076 423812 502077 423876
rect 502011 423811 502077 423812
rect 501827 423740 501893 423741
rect 501827 423676 501828 423740
rect 501892 423676 501893 423740
rect 501827 423675 501893 423676
rect 501830 423469 501890 423675
rect 501827 423468 501893 423469
rect 501827 423404 501828 423468
rect 501892 423404 501893 423468
rect 501827 423403 501893 423404
rect 502011 414084 502077 414085
rect 502011 414020 502012 414084
rect 502076 414020 502077 414084
rect 502011 414019 502077 414020
rect 502014 413810 502074 414019
rect 502195 413812 502261 413813
rect 502195 413810 502196 413812
rect 502014 413750 502196 413810
rect 502195 413748 502196 413750
rect 502260 413748 502261 413812
rect 502195 413747 502261 413748
rect 501646 408446 501890 408506
rect 501830 405789 501890 408446
rect 501827 405788 501893 405789
rect 501827 405724 501828 405788
rect 501892 405724 501893 405788
rect 501827 405723 501893 405724
rect 501827 405652 501893 405653
rect 501827 405588 501828 405652
rect 501892 405588 501893 405652
rect 501827 405587 501893 405588
rect 501459 403748 501525 403749
rect 501459 403684 501460 403748
rect 501524 403684 501525 403748
rect 501459 403683 501525 403684
rect 501830 400893 501890 405587
rect 501827 400892 501893 400893
rect 501827 400828 501828 400892
rect 501892 400828 501893 400892
rect 501827 400827 501893 400828
rect 502195 400892 502261 400893
rect 502195 400828 502196 400892
rect 502260 400828 502261 400892
rect 502195 400827 502261 400828
rect 501827 400756 501893 400757
rect 501827 400692 501828 400756
rect 501892 400692 501893 400756
rect 501827 400691 501893 400692
rect 501830 398170 501890 400691
rect 502011 398716 502077 398717
rect 502011 398652 502012 398716
rect 502076 398652 502077 398716
rect 502011 398651 502077 398652
rect 501646 398110 501890 398170
rect 501646 391917 501706 398110
rect 501643 391916 501709 391917
rect 501643 391852 501644 391916
rect 501708 391852 501709 391916
rect 501643 391851 501709 391852
rect 501827 391780 501893 391781
rect 501827 391716 501828 391780
rect 501892 391716 501893 391780
rect 501827 391715 501893 391716
rect 501459 385116 501525 385117
rect 501459 385052 501460 385116
rect 501524 385052 501525 385116
rect 501459 385051 501525 385052
rect 501462 358597 501522 385051
rect 501830 379130 501890 391715
rect 502014 385117 502074 398651
rect 502198 394637 502258 400827
rect 502195 394636 502261 394637
rect 502195 394572 502196 394636
rect 502260 394572 502261 394636
rect 502195 394571 502261 394572
rect 502195 387156 502261 387157
rect 502195 387092 502196 387156
rect 502260 387092 502261 387156
rect 502195 387091 502261 387092
rect 502011 385116 502077 385117
rect 502011 385052 502012 385116
rect 502076 385052 502077 385116
rect 502011 385051 502077 385052
rect 502198 379810 502258 387091
rect 501646 379070 501890 379130
rect 502014 379750 502258 379810
rect 501459 358596 501525 358597
rect 501459 358532 501460 358596
rect 501524 358532 501525 358596
rect 501459 358531 501525 358532
rect 501275 351660 501341 351661
rect 501275 351596 501276 351660
rect 501340 351596 501341 351660
rect 501275 351595 501341 351596
rect 501459 350572 501525 350573
rect 501459 350570 501460 350572
rect 501094 350510 501460 350570
rect 501459 350508 501460 350510
rect 501524 350508 501525 350572
rect 501459 350507 501525 350508
rect 501459 349892 501525 349893
rect 501459 349890 501460 349892
rect 499990 349830 500234 349890
rect 499254 349558 500050 349618
rect 498886 349150 499166 349210
rect 498886 347170 498946 349150
rect 499990 348530 500050 349558
rect 499806 348470 500050 348530
rect 498886 347110 499314 347170
rect 498702 346294 499130 346354
rect 498702 345130 498762 345662
rect 498702 345070 498946 345130
rect 498886 344450 498946 345070
rect 497966 311070 498394 311130
rect 498702 344390 498946 344450
rect 497966 305010 498026 311070
rect 497966 304950 498246 305010
rect 498702 304330 498762 344390
rect 499070 324138 499130 346294
rect 499254 330850 499314 347110
rect 499806 346490 499866 348470
rect 500174 347850 500234 349830
rect 499622 346430 499866 346490
rect 499990 347790 500234 347850
rect 500542 349830 500786 349890
rect 500910 349830 501460 349890
rect 499254 330790 499498 330850
rect 499438 322690 499498 330790
rect 499622 326770 499682 346430
rect 499990 341818 500050 347790
rect 500542 347170 500602 349830
rect 500910 349618 500970 349830
rect 501459 349828 501460 349830
rect 501524 349828 501525 349892
rect 501459 349827 501525 349828
rect 500358 347110 500602 347170
rect 500726 349558 500970 349618
rect 500358 345898 500418 347110
rect 500726 341730 500786 349558
rect 501278 348530 501338 349062
rect 500358 341670 500786 341730
rect 500910 348470 501338 348530
rect 500358 341050 500418 341670
rect 499806 340990 500418 341050
rect 499806 332890 499866 340990
rect 499806 332830 500234 332890
rect 499622 326710 500050 326770
rect 498886 322630 499498 322690
rect 498886 320650 498946 322630
rect 498886 320590 499130 320650
rect 499070 319970 499130 320590
rect 498518 304270 498762 304330
rect 498886 319910 499130 319970
rect 498518 300930 498578 304270
rect 498886 303738 498946 319910
rect 499438 312490 499498 321862
rect 499990 319290 500050 326710
rect 499070 312430 499498 312490
rect 499622 319230 500050 319290
rect 499070 304330 499130 312430
rect 499070 304270 499498 304330
rect 499438 302970 499498 304270
rect 498334 300870 498578 300930
rect 498886 302910 499498 302970
rect 498334 298210 498394 300870
rect 498334 298150 498578 298210
rect 497782 293390 498026 293450
rect 497598 291350 497842 291410
rect 497782 290730 497842 291350
rect 497598 290670 497842 290730
rect 101630 281830 101874 281890
rect 101814 254010 101874 281830
rect 497598 269738 497658 290670
rect 497966 290186 498026 293390
rect 497782 290126 498026 290186
rect 497782 282570 497842 290126
rect 498150 285970 498210 294662
rect 498518 287418 498578 298150
rect 498886 286650 498946 302910
rect 499254 289458 499314 302142
rect 499622 300250 499682 319230
rect 499622 300190 500050 300250
rect 499990 293450 500050 300190
rect 499622 293390 500050 293450
rect 499622 288690 499682 293390
rect 499254 288630 499682 288690
rect 499254 287418 499314 288630
rect 498886 286590 499682 286650
rect 498150 285910 498946 285970
rect 497782 282510 498026 282570
rect 497598 260218 497658 266102
rect 497966 264298 498026 282510
rect 498150 266250 498210 285142
rect 498886 284018 498946 285910
rect 498518 280618 498578 283782
rect 499254 281978 499314 285822
rect 499622 281482 499682 286590
rect 498886 281422 499682 281482
rect 498886 277810 498946 281422
rect 499254 278578 499314 281062
rect 499806 279170 499866 287862
rect 500174 285378 500234 332830
rect 500358 322690 500418 340222
rect 500358 322630 500786 322690
rect 500726 311130 500786 322630
rect 500542 311070 500786 311130
rect 500542 292770 500602 311070
rect 500542 292710 500786 292770
rect 500726 292090 500786 292710
rect 500358 292030 500786 292090
rect 500358 285970 500418 292030
rect 500910 288690 500970 348470
rect 501459 346492 501525 346493
rect 501459 346490 501460 346492
rect 501094 346430 501460 346490
rect 501094 289370 501154 346430
rect 501459 346428 501460 346430
rect 501524 346428 501525 346492
rect 501459 346427 501525 346428
rect 501459 346356 501525 346357
rect 501459 346292 501460 346356
rect 501524 346292 501525 346356
rect 501459 346291 501525 346292
rect 501462 345810 501522 346291
rect 501278 345750 501522 345810
rect 501278 344861 501338 345750
rect 501275 344860 501341 344861
rect 501275 344796 501276 344860
rect 501340 344796 501341 344860
rect 501275 344795 501341 344796
rect 501459 344316 501525 344317
rect 501459 344252 501460 344316
rect 501524 344252 501525 344316
rect 501459 344251 501525 344252
rect 501462 339690 501522 344251
rect 501278 339630 501522 339690
rect 501278 307730 501338 339630
rect 501459 339012 501525 339013
rect 501459 338948 501460 339012
rect 501524 338948 501525 339012
rect 501459 338947 501525 338948
rect 501462 308410 501522 338947
rect 501646 325685 501706 379070
rect 502014 358730 502074 379750
rect 502014 358670 502258 358730
rect 502011 358596 502077 358597
rect 502011 358532 502012 358596
rect 502076 358532 502077 358596
rect 502011 358531 502077 358532
rect 502014 339013 502074 358531
rect 502198 344997 502258 358670
rect 502195 344996 502261 344997
rect 502195 344932 502196 344996
rect 502260 344932 502261 344996
rect 502195 344931 502261 344932
rect 502011 339012 502077 339013
rect 502011 338948 502012 339012
rect 502076 338948 502077 339012
rect 502011 338947 502077 338948
rect 502011 338876 502077 338877
rect 502011 338812 502012 338876
rect 502076 338812 502077 338876
rect 502011 338811 502077 338812
rect 501643 325684 501709 325685
rect 501643 325620 501644 325684
rect 501708 325620 501709 325684
rect 501643 325619 501709 325620
rect 501827 315892 501893 315893
rect 501827 315828 501828 315892
rect 501892 315828 501893 315892
rect 501827 315827 501893 315828
rect 501830 313170 501890 315827
rect 502014 313850 502074 338811
rect 501968 313790 502074 313850
rect 501968 313306 502028 313790
rect 501968 313246 502074 313306
rect 501646 313110 501890 313170
rect 501646 308549 501706 313110
rect 501643 308548 501709 308549
rect 501643 308484 501644 308548
rect 501708 308484 501709 308548
rect 501643 308483 501709 308484
rect 502014 308410 502074 313246
rect 501462 308350 501706 308410
rect 502014 308350 502258 308410
rect 501278 307670 501522 307730
rect 501462 307050 501522 307670
rect 501278 306990 501522 307050
rect 501278 290050 501338 306990
rect 501646 306917 501706 308350
rect 501459 306916 501525 306917
rect 501459 306852 501460 306916
rect 501524 306852 501525 306916
rect 501459 306851 501525 306852
rect 501643 306916 501709 306917
rect 501643 306852 501644 306916
rect 501708 306852 501709 306916
rect 501643 306851 501709 306852
rect 501462 290325 501522 306851
rect 501830 294898 501890 304862
rect 502011 290460 502077 290461
rect 502011 290396 502012 290460
rect 502076 290396 502077 290460
rect 502011 290395 502077 290396
rect 501459 290324 501525 290325
rect 501459 290260 501460 290324
rect 501524 290260 501525 290324
rect 501459 290259 501525 290260
rect 501459 290052 501525 290053
rect 501459 290050 501460 290052
rect 501278 289990 501460 290050
rect 501459 289988 501460 289990
rect 501524 289988 501525 290052
rect 501459 289987 501525 289988
rect 501094 289310 501522 289370
rect 501275 289100 501341 289101
rect 501275 289036 501276 289100
rect 501340 289036 501341 289100
rect 501275 289035 501341 289036
rect 501278 288690 501338 289035
rect 500910 288630 501338 288690
rect 501462 286381 501522 289310
rect 501643 289100 501709 289101
rect 501643 289036 501644 289100
rect 501708 289036 501709 289100
rect 501643 289035 501709 289036
rect 501459 286380 501525 286381
rect 501459 286316 501460 286380
rect 501524 286316 501525 286380
rect 501459 286315 501525 286316
rect 500358 285910 501522 285970
rect 501275 284748 501341 284749
rect 501275 284746 501276 284748
rect 499622 279110 499866 279170
rect 499990 284686 501276 284746
rect 499990 279170 500050 284686
rect 501275 284684 501276 284686
rect 501340 284684 501341 284748
rect 501275 284683 501341 284684
rect 501462 284610 501522 285910
rect 501278 284550 501522 284610
rect 500726 283250 500786 283782
rect 500726 283190 501154 283250
rect 499990 279110 500234 279170
rect 498886 277750 499314 277810
rect 499254 275770 499314 277750
rect 498702 275710 499314 275770
rect 498702 267882 498762 275710
rect 499622 275090 499682 279110
rect 500174 277810 500234 279110
rect 498886 275030 499682 275090
rect 499990 277750 500234 277810
rect 498886 268970 498946 275030
rect 499254 270418 499314 274262
rect 499990 274138 500050 277750
rect 500358 277130 500418 280382
rect 500174 277070 500418 277130
rect 500174 275906 500234 277070
rect 500174 275846 500418 275906
rect 500358 274410 500418 275846
rect 500726 275042 500786 278342
rect 500358 274350 500602 274410
rect 499990 274078 500418 274138
rect 500358 273322 500418 274078
rect 499622 273262 500418 273322
rect 499622 269058 499682 273262
rect 500174 270330 500234 272902
rect 500542 271098 500602 274350
rect 501094 273818 501154 283190
rect 501278 281485 501338 284550
rect 501459 282436 501525 282437
rect 501459 282372 501460 282436
rect 501524 282372 501525 282436
rect 501459 282371 501525 282372
rect 501275 281484 501341 281485
rect 501275 281420 501276 281484
rect 501340 281420 501341 281484
rect 501275 281419 501341 281420
rect 501462 276450 501522 282371
rect 501646 276589 501706 289035
rect 501827 286380 501893 286381
rect 501827 286316 501828 286380
rect 501892 286316 501893 286380
rect 501827 286315 501893 286316
rect 501643 276588 501709 276589
rect 501643 276524 501644 276588
rect 501708 276524 501709 276588
rect 501643 276523 501709 276524
rect 501462 276390 501706 276450
rect 501459 276316 501525 276317
rect 501459 276252 501460 276316
rect 501524 276252 501525 276316
rect 501459 276251 501525 276252
rect 501462 275229 501522 276251
rect 501459 275228 501525 275229
rect 501459 275164 501460 275228
rect 501524 275164 501525 275228
rect 501459 275163 501525 275164
rect 501459 275092 501525 275093
rect 501459 275090 501460 275092
rect 501278 275030 501460 275090
rect 501278 274141 501338 275030
rect 501459 275028 501460 275030
rect 501524 275028 501525 275092
rect 501459 275027 501525 275028
rect 501459 274956 501525 274957
rect 501459 274892 501460 274956
rect 501524 274892 501525 274956
rect 501459 274891 501525 274892
rect 501275 274140 501341 274141
rect 501275 274076 501276 274140
rect 501340 274076 501341 274140
rect 501275 274075 501341 274076
rect 501462 273189 501522 274891
rect 501646 273325 501706 276390
rect 501830 275909 501890 286315
rect 502014 282301 502074 290395
rect 502011 282300 502077 282301
rect 502011 282236 502012 282300
rect 502076 282236 502077 282300
rect 502011 282235 502077 282236
rect 501827 275908 501893 275909
rect 501827 275844 501828 275908
rect 501892 275844 501893 275908
rect 501827 275843 501893 275844
rect 502198 275090 502258 308350
rect 501830 275030 502258 275090
rect 501643 273324 501709 273325
rect 501643 273260 501644 273324
rect 501708 273260 501709 273324
rect 501643 273259 501709 273260
rect 501459 273188 501525 273189
rect 501459 273124 501460 273188
rect 501524 273124 501525 273188
rect 501459 273123 501525 273124
rect 501459 272916 501525 272917
rect 501459 272852 501460 272916
rect 501524 272852 501525 272916
rect 501459 272851 501525 272852
rect 501462 272642 501522 272851
rect 500910 272582 501522 272642
rect 501643 272644 501709 272645
rect 500174 270270 500786 270330
rect 498886 268910 499314 268970
rect 499254 268378 499314 268910
rect 498702 267822 499866 267882
rect 498150 266190 498578 266250
rect 497966 260130 498026 263382
rect 497966 260070 498394 260130
rect 498334 259450 498394 260070
rect 101630 253950 101874 254010
rect 497782 259390 498394 259450
rect 101630 234378 101690 253950
rect 497782 252738 497842 259390
rect 498150 253418 498210 258622
rect 498150 247210 498210 252502
rect 498518 247210 498578 266190
rect 498886 260130 498946 267462
rect 499806 263530 499866 267822
rect 499990 267610 500050 269502
rect 499990 267550 500234 267610
rect 500174 264298 500234 267550
rect 500726 266930 500786 270270
rect 500910 267066 500970 272582
rect 501643 272580 501644 272644
rect 501708 272580 501709 272644
rect 501643 272579 501709 272580
rect 501459 272508 501525 272509
rect 501459 272444 501460 272508
rect 501524 272444 501525 272508
rect 501459 272443 501525 272444
rect 501275 272372 501341 272373
rect 501275 272370 501276 272372
rect 501094 272310 501276 272370
rect 501094 268290 501154 272310
rect 501275 272308 501276 272310
rect 501340 272308 501341 272372
rect 501275 272307 501341 272308
rect 501275 270876 501341 270877
rect 501275 270812 501276 270876
rect 501340 270812 501341 270876
rect 501275 270811 501341 270812
rect 501278 270469 501338 270811
rect 501275 270468 501341 270469
rect 501275 270404 501276 270468
rect 501340 270404 501341 270468
rect 501275 270403 501341 270404
rect 501275 268292 501341 268293
rect 501275 268290 501276 268292
rect 501094 268230 501276 268290
rect 501275 268228 501276 268230
rect 501340 268228 501341 268292
rect 501275 268227 501341 268228
rect 501275 267068 501341 267069
rect 501275 267066 501276 267068
rect 500910 267006 501276 267066
rect 501275 267004 501276 267006
rect 501340 267004 501341 267068
rect 501275 267003 501341 267004
rect 500726 266870 500970 266930
rect 500542 263666 500602 266102
rect 500910 264298 500970 266870
rect 497598 247150 498210 247210
rect 498334 247150 498578 247210
rect 498702 260070 498946 260130
rect 499070 263470 499866 263530
rect 499990 263606 500602 263666
rect 101630 227490 101690 230062
rect 101630 227430 101874 227490
rect 101814 220690 101874 227430
rect 101630 220630 101874 220690
rect 101630 199610 101690 220630
rect 497598 217378 497658 247150
rect 497966 244898 498026 245022
rect 497782 244838 498026 244898
rect 497782 232930 497842 244838
rect 498334 243130 498394 247150
rect 498702 246210 498762 260070
rect 499070 245714 499130 263470
rect 499438 259538 499498 262702
rect 499990 262442 500050 263606
rect 501275 263532 501341 263533
rect 501275 263530 501276 263532
rect 499806 262382 500050 262442
rect 500174 263470 501276 263530
rect 499438 256050 499498 258622
rect 499806 256186 499866 262382
rect 500174 258858 500234 263470
rect 501275 263468 501276 263470
rect 501340 263468 501341 263532
rect 501275 263467 501341 263468
rect 499806 256126 500234 256186
rect 497966 243070 498394 243130
rect 498886 245654 499130 245714
rect 499254 255990 499498 256050
rect 497966 240410 498026 243070
rect 498334 240410 498394 240942
rect 497966 240350 498394 240410
rect 498886 239050 498946 245654
rect 499254 245170 499314 255990
rect 499070 245110 499314 245170
rect 499070 241498 499130 245110
rect 499622 241770 499682 255494
rect 500174 255098 500234 256126
rect 499990 255038 500234 255098
rect 499990 253194 500050 255038
rect 500542 254554 500602 262702
rect 501275 260268 501341 260269
rect 501275 260204 501276 260268
rect 501340 260204 501341 260268
rect 501275 260203 501341 260204
rect 501278 260130 501338 260203
rect 499806 253134 500050 253194
rect 500174 254494 500602 254554
rect 500726 260070 501338 260130
rect 499806 243810 499866 253134
rect 500174 249114 500234 254494
rect 500726 253330 500786 260070
rect 501094 258770 501154 259302
rect 501275 258772 501341 258773
rect 501275 258770 501276 258772
rect 501094 258710 501276 258770
rect 501275 258708 501276 258710
rect 501340 258708 501341 258772
rect 501275 258707 501341 258708
rect 501275 256732 501341 256733
rect 501275 256730 501276 256732
rect 501094 256670 501276 256730
rect 501094 256138 501154 256670
rect 501275 256668 501276 256670
rect 501340 256668 501341 256732
rect 501275 256667 501341 256668
rect 501462 256325 501522 272443
rect 501646 262445 501706 272579
rect 501830 262850 501890 275030
rect 502011 274956 502077 274957
rect 502011 274892 502012 274956
rect 502076 274892 502077 274956
rect 502011 274891 502077 274892
rect 502014 270605 502074 274891
rect 502195 274140 502261 274141
rect 502195 274076 502196 274140
rect 502260 274076 502261 274140
rect 502195 274075 502261 274076
rect 502011 270604 502077 270605
rect 502011 270540 502012 270604
rect 502076 270540 502077 270604
rect 502011 270539 502077 270540
rect 502011 267204 502077 267205
rect 502011 267140 502012 267204
rect 502076 267140 502077 267204
rect 502011 267139 502077 267140
rect 502014 263397 502074 267139
rect 502011 263396 502077 263397
rect 502011 263332 502012 263396
rect 502076 263332 502077 263396
rect 502011 263331 502077 263332
rect 501830 262790 502074 262850
rect 501643 262444 501709 262445
rect 501643 262380 501644 262444
rect 501708 262380 501709 262444
rect 501643 262379 501709 262380
rect 501827 259860 501893 259861
rect 501827 259796 501828 259860
rect 501892 259796 501893 259860
rect 501827 259795 501893 259796
rect 501830 256730 501890 259795
rect 501646 256670 501890 256730
rect 501459 256324 501525 256325
rect 501459 256260 501460 256324
rect 501524 256260 501525 256324
rect 501459 256259 501525 256260
rect 501459 256188 501525 256189
rect 501459 256124 501460 256188
rect 501524 256124 501525 256188
rect 501459 256123 501525 256124
rect 501462 255642 501522 256123
rect 501278 255582 501522 255642
rect 501278 254010 501338 255582
rect 501646 255509 501706 256670
rect 501827 256324 501893 256325
rect 501827 256260 501828 256324
rect 501892 256260 501893 256324
rect 501827 256259 501893 256260
rect 501643 255508 501709 255509
rect 501643 255444 501644 255508
rect 501708 255444 501709 255508
rect 501643 255443 501709 255444
rect 501643 255372 501709 255373
rect 501643 255308 501644 255372
rect 501708 255308 501709 255372
rect 501643 255307 501709 255308
rect 501646 254149 501706 255307
rect 501830 255101 501890 256259
rect 501827 255100 501893 255101
rect 501827 255036 501828 255100
rect 501892 255036 501893 255100
rect 501827 255035 501893 255036
rect 501827 254556 501893 254557
rect 501827 254492 501828 254556
rect 501892 254492 501893 254556
rect 501827 254491 501893 254492
rect 501643 254148 501709 254149
rect 501643 254084 501644 254148
rect 501708 254084 501709 254148
rect 501643 254083 501709 254084
rect 501278 253950 501706 254010
rect 500726 253270 501154 253330
rect 501094 253194 501154 253270
rect 501275 253196 501341 253197
rect 501275 253194 501276 253196
rect 501094 253134 501276 253194
rect 501275 253132 501276 253134
rect 501340 253132 501341 253196
rect 501275 253131 501341 253132
rect 501459 253196 501525 253197
rect 501459 253132 501460 253196
rect 501524 253132 501525 253196
rect 501459 253131 501525 253132
rect 501094 249658 501154 252502
rect 501275 249660 501341 249661
rect 501275 249658 501276 249660
rect 501094 249598 501276 249658
rect 501275 249596 501276 249598
rect 501340 249596 501341 249660
rect 501275 249595 501341 249596
rect 501462 249389 501522 253131
rect 501646 251973 501706 253950
rect 501643 251972 501709 251973
rect 501643 251908 501644 251972
rect 501708 251908 501709 251972
rect 501643 251907 501709 251908
rect 501643 251836 501709 251837
rect 501643 251772 501644 251836
rect 501708 251772 501709 251836
rect 501643 251771 501709 251772
rect 501459 249388 501525 249389
rect 501459 249324 501460 249388
rect 501524 249324 501525 249388
rect 501459 249323 501525 249324
rect 501459 249116 501525 249117
rect 500174 249054 500418 249114
rect 500358 245170 500418 249054
rect 501459 249052 501460 249116
rect 501524 249052 501525 249116
rect 501459 249051 501525 249052
rect 501462 246669 501522 249051
rect 501459 246668 501525 246669
rect 501459 246604 501460 246668
rect 501524 246604 501525 246668
rect 501459 246603 501525 246604
rect 501459 246124 501525 246125
rect 501459 246060 501460 246124
rect 501524 246060 501525 246124
rect 501459 246059 501525 246060
rect 501462 245714 501522 246059
rect 501094 245654 501522 245714
rect 501094 245258 501154 245654
rect 500358 245110 500786 245170
rect 500726 244626 500786 245110
rect 501459 244628 501525 244629
rect 501459 244626 501460 244628
rect 500726 244566 501460 244626
rect 501459 244564 501460 244566
rect 501524 244564 501525 244628
rect 501459 244563 501525 244564
rect 501459 244492 501525 244493
rect 501459 244490 501460 244492
rect 500910 244430 501460 244490
rect 499806 243750 500050 243810
rect 499622 241710 499866 241770
rect 499070 241438 499682 241498
rect 498518 238990 498946 239050
rect 498518 234290 498578 238990
rect 498886 235058 498946 238222
rect 498518 234230 498946 234290
rect 497782 232870 498062 232930
rect 497966 220282 498026 232102
rect 498518 227578 498578 232782
rect 498886 226810 498946 234230
rect 498334 226750 498946 226810
rect 498334 221642 498394 226750
rect 499254 226674 499314 240942
rect 499622 236330 499682 241438
rect 499438 236270 499682 236330
rect 499438 234970 499498 236270
rect 499438 234910 499682 234970
rect 499622 227490 499682 234910
rect 499806 227626 499866 241710
rect 499990 237690 500050 243750
rect 500358 238458 500418 244342
rect 500910 242722 500970 244430
rect 501459 244428 501460 244430
rect 501524 244428 501525 244492
rect 501459 244427 501525 244428
rect 501459 244356 501525 244357
rect 501459 244292 501460 244356
rect 501524 244292 501525 244356
rect 501459 244291 501525 244292
rect 500910 242662 501338 242722
rect 501278 242589 501338 242662
rect 501275 242588 501341 242589
rect 501275 242524 501276 242588
rect 501340 242524 501341 242588
rect 501275 242523 501341 242524
rect 501462 242453 501522 244291
rect 501646 242725 501706 251771
rect 501830 246530 501890 254491
rect 502014 246666 502074 262790
rect 502198 255645 502258 274075
rect 502195 255644 502261 255645
rect 502195 255580 502196 255644
rect 502260 255580 502261 255644
rect 502195 255579 502261 255580
rect 502195 255508 502261 255509
rect 502195 255444 502196 255508
rect 502260 255444 502261 255508
rect 502195 255443 502261 255444
rect 502198 251837 502258 255443
rect 502195 251836 502261 251837
rect 502195 251772 502196 251836
rect 502260 251772 502261 251836
rect 502195 251771 502261 251772
rect 502014 246606 502258 246666
rect 501830 246470 502074 246530
rect 501827 244628 501893 244629
rect 501827 244564 501828 244628
rect 501892 244564 501893 244628
rect 501827 244563 501893 244564
rect 501643 242724 501709 242725
rect 501643 242660 501644 242724
rect 501708 242660 501709 242724
rect 501643 242659 501709 242660
rect 501459 242452 501525 242453
rect 501459 242388 501460 242452
rect 501524 242388 501525 242452
rect 501830 242450 501890 244563
rect 502014 244493 502074 246470
rect 502198 244901 502258 246606
rect 502195 244900 502261 244901
rect 502195 244836 502196 244900
rect 502260 244836 502261 244900
rect 502195 244835 502261 244836
rect 502195 244764 502261 244765
rect 502195 244700 502196 244764
rect 502260 244700 502261 244764
rect 502195 244699 502261 244700
rect 502011 244492 502077 244493
rect 502011 244428 502012 244492
rect 502076 244428 502077 244492
rect 502011 244427 502077 244428
rect 502011 244220 502077 244221
rect 502011 244156 502012 244220
rect 502076 244156 502077 244220
rect 502011 244155 502077 244156
rect 501459 242387 501525 242388
rect 501646 242390 501890 242450
rect 501459 242180 501525 242181
rect 501459 242116 501460 242180
rect 501524 242116 501525 242180
rect 501459 242115 501525 242116
rect 501462 242042 501522 242115
rect 501646 242045 501706 242390
rect 501827 242316 501893 242317
rect 501827 242252 501828 242316
rect 501892 242252 501893 242316
rect 501827 242251 501893 242252
rect 501094 241982 501522 242042
rect 501643 242044 501709 242045
rect 501094 238458 501154 241982
rect 501643 241980 501644 242044
rect 501708 241980 501709 242044
rect 501643 241979 501709 241980
rect 501459 241500 501525 241501
rect 501459 241436 501460 241500
rect 501524 241436 501525 241500
rect 501459 241435 501525 241436
rect 501643 241500 501709 241501
rect 501643 241436 501644 241500
rect 501708 241436 501709 241500
rect 501643 241435 501709 241436
rect 501275 238100 501341 238101
rect 501275 238098 501276 238100
rect 500726 238038 501276 238098
rect 499990 237630 500418 237690
rect 500358 234970 500418 237630
rect 500726 234970 500786 238038
rect 501275 238036 501276 238038
rect 501340 238036 501341 238100
rect 501275 238035 501341 238036
rect 501462 237829 501522 241435
rect 501646 237829 501706 241435
rect 501830 238101 501890 242251
rect 501827 238100 501893 238101
rect 501827 238036 501828 238100
rect 501892 238036 501893 238100
rect 501827 238035 501893 238036
rect 501459 237828 501525 237829
rect 501459 237764 501460 237828
rect 501524 237764 501525 237828
rect 501459 237763 501525 237764
rect 501643 237828 501709 237829
rect 501643 237764 501644 237828
rect 501708 237764 501709 237828
rect 501643 237763 501709 237764
rect 501827 237692 501893 237693
rect 501827 237628 501828 237692
rect 501892 237628 501893 237692
rect 501827 237627 501893 237628
rect 501459 237556 501525 237557
rect 501094 237494 501338 237554
rect 501094 237098 501154 237494
rect 501278 237285 501338 237494
rect 501459 237492 501460 237556
rect 501524 237492 501525 237556
rect 501459 237491 501525 237492
rect 501643 237556 501709 237557
rect 501643 237492 501644 237556
rect 501708 237492 501709 237556
rect 501643 237491 501709 237492
rect 501275 237284 501341 237285
rect 501275 237220 501276 237284
rect 501340 237220 501341 237284
rect 501275 237219 501341 237220
rect 501275 235788 501341 235789
rect 501275 235786 501276 235788
rect 500174 234910 500418 234970
rect 500542 234910 500786 234970
rect 500910 235726 501276 235786
rect 500174 233018 500234 234910
rect 500542 234378 500602 234910
rect 500910 233610 500970 235726
rect 501275 235724 501276 235726
rect 501340 235724 501341 235788
rect 501275 235723 501341 235724
rect 501275 235652 501341 235653
rect 501275 235588 501276 235652
rect 501340 235588 501341 235652
rect 501275 235587 501341 235588
rect 500542 233550 500970 233610
rect 500542 228170 500602 233550
rect 500542 228110 500786 228170
rect 499806 227566 500602 227626
rect 499622 227430 500418 227490
rect 498886 226614 499314 226674
rect 498886 226130 498946 226614
rect 499990 226130 500050 226662
rect 498702 226070 498946 226130
rect 499438 226070 500050 226130
rect 498334 221582 498578 221642
rect 497966 220222 498394 220282
rect 497966 217290 498026 219182
rect 497966 217230 498210 217290
rect 498150 215794 498210 217230
rect 497598 215734 498210 215794
rect 497598 201650 497658 215734
rect 498334 215250 498394 220222
rect 497966 215190 498394 215250
rect 497598 201590 497842 201650
rect 101594 199550 101690 199610
rect 101630 179890 101690 196062
rect 497782 194850 497842 201590
rect 497966 195530 498026 215190
rect 498518 214570 498578 221582
rect 498150 214510 498578 214570
rect 498702 214570 498762 226070
rect 499070 220010 499130 222582
rect 499438 221506 499498 226070
rect 500358 224090 500418 227430
rect 500138 224030 500418 224090
rect 499438 221446 499682 221506
rect 499622 220778 499682 221446
rect 498886 219950 499130 220010
rect 498886 215794 498946 219950
rect 499070 219862 499350 219874
rect 499070 219814 499498 219862
rect 499070 216338 499130 219814
rect 499622 216698 499682 219182
rect 499070 216278 499866 216338
rect 498886 215734 499682 215794
rect 498702 214510 498946 214570
rect 498150 206410 498210 214510
rect 498886 213890 498946 214510
rect 498518 213830 498946 213890
rect 498518 207090 498578 213830
rect 498886 209898 498946 212382
rect 498886 207770 498946 208982
rect 499254 208450 499314 209662
rect 499622 209218 499682 215734
rect 499806 213210 499866 216278
rect 499990 214570 500050 223262
rect 500542 222594 500602 227566
rect 500726 223682 500786 228110
rect 500910 224906 500970 232782
rect 501278 225181 501338 235587
rect 501275 225180 501341 225181
rect 501275 225116 501276 225180
rect 501340 225116 501341 225180
rect 501275 225115 501341 225116
rect 501275 224908 501341 224909
rect 501275 224906 501276 224908
rect 500910 224846 501276 224906
rect 501275 224844 501276 224846
rect 501340 224844 501341 224908
rect 501275 224843 501341 224844
rect 501462 223685 501522 237491
rect 501459 223684 501525 223685
rect 500726 223622 500970 223682
rect 500910 223498 500970 223622
rect 501459 223620 501460 223684
rect 501524 223620 501525 223684
rect 501459 223619 501525 223620
rect 501459 222596 501525 222597
rect 500542 222534 501338 222594
rect 501278 222189 501338 222534
rect 501459 222532 501460 222596
rect 501524 222532 501525 222596
rect 501459 222531 501525 222532
rect 501275 222188 501341 222189
rect 501275 222124 501276 222188
rect 501340 222124 501341 222188
rect 501275 222123 501341 222124
rect 501275 221644 501341 221645
rect 501275 221642 501276 221644
rect 500174 221582 501276 221642
rect 500174 216338 500234 221582
rect 501275 221580 501276 221582
rect 501340 221580 501341 221644
rect 501275 221579 501341 221580
rect 501275 221508 501341 221509
rect 501275 221444 501276 221508
rect 501340 221444 501341 221508
rect 501275 221443 501341 221444
rect 501278 220098 501338 221443
rect 501462 220285 501522 222531
rect 501459 220284 501525 220285
rect 501459 220220 501460 220284
rect 501524 220220 501525 220284
rect 501459 220219 501525 220220
rect 501459 219740 501525 219741
rect 501459 219676 501460 219740
rect 501524 219676 501525 219740
rect 501459 219675 501525 219676
rect 501462 219330 501522 219675
rect 500726 219270 501522 219330
rect 500174 216278 500418 216338
rect 500358 215338 500418 216278
rect 499990 214510 500270 214570
rect 499806 213150 500050 213210
rect 499254 208390 499682 208450
rect 498886 207710 499314 207770
rect 498518 207030 498946 207090
rect 498150 206350 498762 206410
rect 498334 198114 498394 205582
rect 498702 204370 498762 206350
rect 498518 204310 498762 204370
rect 498518 198930 498578 204310
rect 498886 199338 498946 207030
rect 499254 205050 499314 207710
rect 499622 205818 499682 208390
rect 499254 204990 499682 205050
rect 499254 202058 499314 202862
rect 499622 202330 499682 204990
rect 499070 201998 499314 202058
rect 499438 202270 499682 202330
rect 499990 202330 500050 213150
rect 500174 203282 500234 213742
rect 500726 213210 500786 219270
rect 501459 215932 501525 215933
rect 501459 215868 501460 215932
rect 501524 215868 501525 215932
rect 501459 215867 501525 215868
rect 500726 213150 500970 213210
rect 500910 208450 500970 213150
rect 500726 208390 500970 208450
rect 500726 203282 500786 208390
rect 501094 203418 501154 215102
rect 501275 211580 501341 211581
rect 501275 211516 501276 211580
rect 501340 211516 501341 211580
rect 501275 211515 501341 211516
rect 501278 203693 501338 211515
rect 501462 204917 501522 215867
rect 501459 204916 501525 204917
rect 501459 204852 501460 204916
rect 501524 204852 501525 204916
rect 501459 204851 501525 204852
rect 501275 203692 501341 203693
rect 501275 203628 501276 203692
rect 501340 203628 501341 203692
rect 501275 203627 501341 203628
rect 501459 203420 501525 203421
rect 501459 203418 501460 203420
rect 501094 203358 501460 203418
rect 501459 203356 501460 203358
rect 501524 203356 501525 203420
rect 501459 203355 501525 203356
rect 501459 203284 501525 203285
rect 501459 203282 501460 203284
rect 500174 203222 500418 203282
rect 500726 203222 501460 203282
rect 500358 203010 500418 203222
rect 501459 203220 501460 203222
rect 501524 203220 501525 203284
rect 501459 203219 501525 203220
rect 501275 203148 501341 203149
rect 501275 203098 501276 203148
rect 501340 203098 501341 203148
rect 500358 202950 500786 203010
rect 499990 202270 500234 202330
rect 499070 199474 499130 201998
rect 499070 199414 499314 199474
rect 498886 199278 499130 199338
rect 498518 198870 498946 198930
rect 498150 198054 498394 198114
rect 498150 196890 498210 198054
rect 498518 196890 498578 197422
rect 498150 196830 498578 196890
rect 497966 195470 498210 195530
rect 497782 194790 498026 194850
rect 101630 179830 101726 179890
rect 101778 177790 101874 177850
rect 101814 171730 101874 177790
rect 101630 171670 101874 171730
rect 101630 132970 101690 171670
rect 101630 132910 101874 132970
rect 101814 123994 101874 132910
rect 101262 123934 101874 123994
rect 107699 123996 107765 123997
rect 93715 123316 93781 123317
rect 93715 123252 93716 123316
rect 93780 123252 93781 123316
rect 93715 123251 93781 123252
rect 93718 121685 93778 123251
rect 99235 122908 99301 122909
rect 99235 122858 99236 122908
rect 99300 122858 99301 122908
rect 93715 121684 93781 121685
rect 93715 121620 93716 121684
rect 93780 121620 93781 121684
rect 93715 121619 93781 121620
rect 94404 96054 95004 122000
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 92427 3908 92493 3909
rect 92427 3844 92428 3908
rect 92492 3844 92493 3908
rect 92427 3843 92493 3844
rect 93531 3908 93597 3909
rect 93531 3844 93532 3908
rect 93596 3844 93597 3908
rect 93531 3843 93597 3844
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 99654 98604 122000
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 101262 2957 101322 123934
rect 107699 123932 107700 123996
rect 107764 123932 107765 123996
rect 107699 123931 107765 123932
rect 463555 123996 463621 123997
rect 463555 123932 463556 123996
rect 463620 123932 463621 123996
rect 463555 123931 463621 123932
rect 491891 123996 491957 123997
rect 491891 123932 491892 123996
rect 491956 123932 491957 123996
rect 491891 123931 491957 123932
rect 493547 123996 493613 123997
rect 493547 123932 493548 123996
rect 493612 123932 493613 123996
rect 493547 123931 493613 123932
rect 101604 103254 102204 122000
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 101259 2956 101325 2957
rect 101259 2892 101260 2956
rect 101324 2892 101325 2956
rect 101259 2891 101325 2892
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 107702 3093 107762 123931
rect 122787 123860 122853 123861
rect 122787 123796 122788 123860
rect 122852 123796 122853 123860
rect 122787 123795 122853 123796
rect 425467 123860 425533 123861
rect 425467 123796 425468 123860
rect 425532 123796 425533 123860
rect 425467 123795 425533 123796
rect 114326 122710 114754 122770
rect 114326 122637 114386 122710
rect 114694 122637 114754 122710
rect 114323 122636 114389 122637
rect 114323 122572 114324 122636
rect 114388 122572 114389 122636
rect 114323 122571 114389 122572
rect 114691 122636 114757 122637
rect 114691 122572 114692 122636
rect 114756 122572 114757 122636
rect 114691 122571 114757 122572
rect 114691 122228 114757 122229
rect 114691 122164 114692 122228
rect 114756 122164 114757 122228
rect 114691 122163 114757 122164
rect 114694 122090 114754 122163
rect 114326 122030 114754 122090
rect 108804 110454 109404 122000
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 107699 3092 107765 3093
rect 107699 3028 107700 3092
rect 107764 3028 107765 3092
rect 107699 3027 107765 3028
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 114054 113004 122000
rect 114326 121141 114386 122030
rect 114323 121140 114389 121141
rect 114323 121076 114324 121140
rect 114388 121076 114389 121140
rect 114323 121075 114389 121076
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 116004 117654 116604 122000
rect 116715 121412 116781 121413
rect 116715 121348 116716 121412
rect 116780 121348 116781 121412
rect 116715 121347 116781 121348
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 114875 2892 114876 2942
rect 114940 2892 114941 2942
rect 114875 2891 114941 2892
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 -4026 116604 9098
rect 116718 3773 116778 121347
rect 119604 121254 120204 122000
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 116715 3772 116781 3773
rect 116715 3708 116716 3772
rect 116780 3708 116781 3772
rect 116715 3707 116781 3708
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 122790 3501 122850 123795
rect 207059 123724 207125 123725
rect 207059 123660 207060 123724
rect 207124 123660 207125 123724
rect 207059 123659 207125 123660
rect 320035 123724 320101 123725
rect 320035 123660 320036 123724
rect 320100 123660 320101 123724
rect 320035 123659 320101 123660
rect 172467 122636 172533 122637
rect 172467 122572 172468 122636
rect 172532 122572 172533 122636
rect 172467 122571 172533 122572
rect 126804 92454 127404 122000
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 125550 3710 125794 3770
rect 125550 3501 125610 3710
rect 125734 3501 125794 3710
rect 122787 3500 122853 3501
rect 122787 3436 122788 3500
rect 122852 3436 122853 3500
rect 122787 3435 122853 3436
rect 125547 3500 125613 3501
rect 125547 3436 125548 3500
rect 125612 3436 125613 3500
rect 125547 3435 125613 3436
rect 125731 3500 125797 3501
rect 125731 3436 125732 3500
rect 125796 3436 125797 3500
rect 125731 3435 125797 3436
rect 126804 -1266 127404 19898
rect 130404 96054 131004 122000
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 127906 3030 128406 3090
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 -3106 131004 23498
rect 134004 99654 134604 122000
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 133827 3500 133893 3501
rect 133827 3436 133828 3500
rect 133892 3436 133893 3500
rect 133827 3435 133893 3436
rect 133830 2957 133890 3435
rect 133827 2956 133893 2957
rect 133827 2892 133828 2956
rect 133892 2892 133893 2956
rect 133827 2891 133893 2892
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 103254 138204 122000
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 110454 145404 122000
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 143579 3500 143645 3501
rect 143579 3436 143580 3500
rect 143644 3436 143645 3500
rect 143579 3435 143645 3436
rect 143582 2957 143642 3435
rect 143579 2956 143645 2957
rect 143579 2892 143580 2956
rect 143644 2892 143645 2956
rect 143579 2891 143645 2892
rect 144804 2454 145404 37898
rect 148182 3501 148242 121942
rect 148404 114054 149004 122000
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148179 3500 148245 3501
rect 148179 3436 148180 3500
rect 148244 3436 148245 3500
rect 148179 3435 148245 3436
rect 147226 3030 147726 3090
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 117654 152604 122000
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 155604 121254 156204 122000
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 152779 70412 152845 70413
rect 152779 70348 152780 70412
rect 152844 70348 152845 70412
rect 152779 70347 152845 70348
rect 152782 67693 152842 70347
rect 152779 67692 152845 67693
rect 152779 67628 152780 67692
rect 152844 67628 152845 67692
rect 152779 67627 152845 67628
rect 152963 61436 153029 61437
rect 152963 61372 152964 61436
rect 153028 61372 153029 61436
rect 152963 61371 153029 61372
rect 152966 50965 153026 61371
rect 152963 50964 153029 50965
rect 152963 50900 152964 50964
rect 153028 50900 153029 50964
rect 152963 50899 153029 50900
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 153147 3500 153213 3501
rect 153147 3436 153148 3500
rect 153212 3436 153213 3500
rect 153147 3435 153213 3436
rect 153150 2957 153210 3435
rect 153147 2956 153213 2957
rect 153147 2892 153148 2956
rect 153212 2892 153213 2956
rect 153147 2891 153213 2892
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 92454 163404 122000
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 164006 3773 164066 119902
rect 166404 96054 167004 122000
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 164003 3772 164069 3773
rect 164003 3708 164004 3772
rect 164068 3708 164069 3772
rect 164003 3707 164069 3708
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 -3106 167004 23498
rect 170004 99654 170604 122000
rect 172470 121821 172530 122571
rect 172467 121820 172533 121821
rect 172467 121756 172468 121820
rect 172532 121756 172533 121820
rect 172467 121755 172533 121756
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 169155 4452 169221 4453
rect 169155 4388 169156 4452
rect 169220 4388 169221 4452
rect 169155 4387 169221 4388
rect 169158 3858 169218 4387
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 -4946 170604 27098
rect 173604 103254 174204 122000
rect 176150 121410 176210 123302
rect 191790 122710 192034 122770
rect 191790 122365 191850 122710
rect 191974 122637 192034 122710
rect 191971 122636 192037 122637
rect 191971 122572 191972 122636
rect 192036 122572 192037 122636
rect 191971 122571 192037 122572
rect 191787 122364 191853 122365
rect 191787 122300 191788 122364
rect 191852 122300 191853 122364
rect 191787 122299 191853 122300
rect 176150 121350 176578 121410
rect 174494 118693 174554 119902
rect 174491 118692 174557 118693
rect 174491 118628 174492 118692
rect 174556 118628 174557 118692
rect 174491 118627 174557 118628
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 172467 4452 172533 4453
rect 172467 4388 172468 4452
rect 172532 4388 172533 4452
rect 172467 4387 172533 4388
rect 172470 3858 172530 4387
rect 172467 3500 172533 3501
rect 172467 3436 172468 3500
rect 172532 3436 172533 3500
rect 172467 3435 172533 3436
rect 172470 2957 172530 3435
rect 172467 2956 172533 2957
rect 172467 2892 172468 2956
rect 172532 2892 172533 2956
rect 172467 2891 172533 2892
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 176518 3501 176578 121350
rect 180804 110454 181404 122000
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 176515 3500 176581 3501
rect 176515 3436 176516 3500
rect 176580 3436 176581 3500
rect 176515 3435 176581 3436
rect 180804 2454 181404 37898
rect 184404 114054 185004 122000
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 117654 188604 122000
rect 191604 121254 192204 122000
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 85254 192204 120698
rect 193259 120188 193325 120189
rect 193259 120138 193260 120188
rect 193324 120138 193325 120188
rect 196571 120188 196637 120189
rect 196571 120124 196572 120188
rect 196636 120124 196637 120188
rect 196571 120123 196637 120124
rect 196574 119458 196634 120123
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 92454 199404 122000
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 96054 203004 122000
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 206004 99654 206604 122000
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 205186 3030 205686 3090
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 -4946 206604 27098
rect 207062 3773 207122 123659
rect 218099 123588 218165 123589
rect 218099 123524 218100 123588
rect 218164 123524 218165 123588
rect 234107 123588 234173 123589
rect 234107 123538 234108 123588
rect 234172 123538 234173 123588
rect 235211 123588 235277 123589
rect 235211 123538 235212 123588
rect 235276 123538 235277 123588
rect 240179 123588 240245 123589
rect 240179 123538 240180 123588
rect 240244 123538 240245 123588
rect 253059 123588 253125 123589
rect 253059 123538 253060 123588
rect 253124 123538 253125 123588
rect 275875 123588 275941 123589
rect 218099 123523 218165 123524
rect 209819 123252 209820 123302
rect 209884 123252 209885 123302
rect 209819 123251 209885 123252
rect 209604 103254 210204 122000
rect 215155 121892 215156 121942
rect 215220 121892 215221 121942
rect 215155 121891 215221 121892
rect 215523 121892 215524 121942
rect 215588 121892 215589 121942
rect 215523 121891 215589 121892
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 207059 3772 207125 3773
rect 207059 3708 207060 3772
rect 207124 3708 207125 3772
rect 207059 3707 207125 3708
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 110454 217404 122000
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 218102 3773 218162 123523
rect 252507 123452 252573 123453
rect 252507 123388 252508 123452
rect 252572 123388 252573 123452
rect 252507 123387 252573 123388
rect 219203 123252 219204 123302
rect 219268 123252 219269 123302
rect 219203 123251 219269 123252
rect 237235 122772 237301 122773
rect 230430 122710 230674 122770
rect 230430 122229 230490 122710
rect 230427 122228 230493 122229
rect 230427 122164 230428 122228
rect 230492 122164 230493 122228
rect 230427 122163 230493 122164
rect 220404 114054 221004 122000
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 218099 3772 218165 3773
rect 218099 3708 218100 3772
rect 218164 3708 218165 3772
rect 218099 3707 218165 3708
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 117654 224604 122000
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 121254 228204 122000
rect 230614 121685 230674 122710
rect 237235 122708 237236 122772
rect 237300 122708 237301 122772
rect 237235 122707 237301 122708
rect 230611 121684 230677 121685
rect 230611 121620 230612 121684
rect 230676 121620 230677 121684
rect 230611 121619 230677 121620
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 92454 235404 122000
rect 237238 121957 237298 122707
rect 237235 121956 237301 121957
rect 237235 121892 237236 121956
rect 237300 121892 237301 121956
rect 237235 121891 237301 121892
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 96054 239004 122000
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 99654 242604 122000
rect 243494 121821 243554 121942
rect 243491 121820 243557 121821
rect 243491 121756 243492 121820
rect 243556 121756 243557 121820
rect 243491 121755 243557 121756
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 245604 103254 246204 122000
rect 251222 118693 251282 119902
rect 251219 118692 251285 118693
rect 251219 118628 251220 118692
rect 251284 118628 251285 118692
rect 251219 118627 251285 118628
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 243826 3710 244290 3770
rect 244230 3178 244290 3710
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252510 3093 252570 123387
rect 275875 123524 275876 123588
rect 275940 123524 275941 123588
rect 275875 123523 275941 123524
rect 271643 123180 271709 123181
rect 271643 123116 271644 123180
rect 271708 123116 271709 123180
rect 271643 123115 271709 123116
rect 258730 122710 259230 122770
rect 269067 122228 269133 122229
rect 252804 110454 253404 122000
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252507 3092 252573 3093
rect 252507 3028 252508 3092
rect 252572 3028 252573 3092
rect 252507 3027 252573 3028
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 114054 257004 122000
rect 269067 122164 269068 122228
rect 269132 122164 269133 122228
rect 269067 122163 269133 122164
rect 259318 121821 259378 121942
rect 259315 121820 259381 121821
rect 259315 121756 259316 121820
rect 259380 121756 259381 121820
rect 259315 121755 259381 121756
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 117654 260604 122000
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 121254 264204 122000
rect 269070 121821 269130 122163
rect 269067 121820 269133 121821
rect 269067 121756 269068 121820
rect 269132 121756 269133 121820
rect 269067 121755 269133 121756
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 92454 271404 122000
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 268886 2957 268946 3622
rect 268883 2956 268949 2957
rect 264467 2892 264468 2942
rect 264532 2892 264533 2942
rect 264467 2891 264533 2892
rect 268883 2892 268884 2956
rect 268948 2892 268949 2956
rect 268883 2891 268949 2892
rect 270804 -1266 271404 19898
rect 271646 3773 271706 123115
rect 273670 118693 273730 119222
rect 273667 118692 273733 118693
rect 273667 118628 273668 118692
rect 273732 118628 273733 118692
rect 273667 118627 273733 118628
rect 274404 96054 275004 122000
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 271643 3772 271709 3773
rect 271643 3708 271644 3772
rect 271708 3708 271709 3772
rect 271643 3707 271709 3708
rect 273302 3770 273362 4302
rect 272898 3710 273362 3770
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 -3106 275004 23498
rect 275878 4045 275938 123523
rect 277347 123452 277413 123453
rect 277347 123388 277348 123452
rect 277412 123450 277413 123452
rect 295195 123452 295261 123453
rect 277412 123390 277594 123450
rect 277412 123388 277413 123390
rect 277347 123387 277413 123388
rect 277534 123317 277594 123390
rect 295195 123388 295196 123452
rect 295260 123388 295261 123452
rect 295195 123387 295261 123388
rect 296667 123452 296733 123453
rect 296667 123388 296668 123452
rect 296732 123450 296733 123452
rect 314515 123452 314581 123453
rect 296732 123390 296914 123450
rect 296732 123388 296733 123390
rect 296667 123387 296733 123388
rect 277531 123316 277597 123317
rect 277531 123252 277532 123316
rect 277596 123252 277597 123316
rect 277531 123251 277597 123252
rect 285627 123316 285693 123317
rect 285627 123252 285628 123316
rect 285692 123252 285693 123316
rect 285627 123251 285693 123252
rect 285630 123045 285690 123251
rect 295198 123045 295258 123387
rect 296854 123317 296914 123390
rect 314515 123388 314516 123452
rect 314580 123388 314581 123452
rect 314515 123387 314581 123388
rect 315987 123452 316053 123453
rect 315987 123388 315988 123452
rect 316052 123450 316053 123452
rect 316052 123390 316234 123450
rect 316052 123388 316053 123390
rect 315987 123387 316053 123388
rect 296851 123316 296917 123317
rect 296851 123252 296852 123316
rect 296916 123252 296917 123316
rect 296851 123251 296917 123252
rect 304947 123316 305013 123317
rect 304947 123252 304948 123316
rect 305012 123252 305013 123316
rect 304947 123251 305013 123252
rect 304950 123045 305010 123251
rect 314518 123045 314578 123387
rect 316174 123317 316234 123390
rect 316171 123316 316237 123317
rect 316171 123252 316172 123316
rect 316236 123252 316237 123316
rect 316171 123251 316237 123252
rect 285627 123044 285693 123045
rect 285627 122980 285628 123044
rect 285692 122980 285693 123044
rect 285627 122979 285693 122980
rect 295195 123044 295261 123045
rect 295195 122980 295196 123044
rect 295260 122980 295261 123044
rect 295195 122979 295261 122980
rect 304947 123044 305013 123045
rect 304947 122980 304948 123044
rect 305012 122980 305013 123044
rect 304947 122979 305013 122980
rect 314515 123044 314581 123045
rect 314515 122980 314516 123044
rect 314580 122980 314581 123044
rect 314515 122979 314581 122980
rect 299430 122710 299674 122770
rect 299430 122229 299490 122710
rect 299614 122229 299674 122710
rect 288387 122228 288453 122229
rect 278004 99654 278604 122000
rect 288387 122164 288388 122228
rect 288452 122164 288453 122228
rect 299427 122228 299493 122229
rect 288387 122163 288453 122164
rect 281214 121821 281274 121942
rect 281211 121820 281277 121821
rect 281211 121756 281212 121820
rect 281276 121756 281277 121820
rect 281211 121755 281277 121756
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 275875 4044 275941 4045
rect 275875 3980 275876 4044
rect 275940 3980 275941 4044
rect 275875 3979 275941 3980
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 103254 282204 122000
rect 288390 121685 288450 122163
rect 288387 121684 288453 121685
rect 288387 121620 288388 121684
rect 288452 121620 288453 121684
rect 288387 121619 288453 121620
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 110454 289404 122000
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 292404 114054 293004 122000
rect 299427 122164 299428 122228
rect 299492 122164 299493 122228
rect 299427 122163 299493 122164
rect 299611 122228 299677 122229
rect 299611 122164 299612 122228
rect 299676 122164 299677 122228
rect 299611 122163 299677 122164
rect 293174 121821 293234 121942
rect 293171 121820 293237 121821
rect 293171 121756 293172 121820
rect 293236 121756 293237 121820
rect 293171 121755 293237 121756
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 289675 97068 289741 97069
rect 289675 97004 289676 97068
rect 289740 97004 289741 97068
rect 289675 97003 289741 97004
rect 289678 96661 289738 97003
rect 289675 96660 289741 96661
rect 289675 96596 289676 96660
rect 289740 96596 289741 96660
rect 289675 96595 289741 96596
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288387 3636 288453 3637
rect 288387 3572 288388 3636
rect 288452 3572 288453 3636
rect 288387 3571 288453 3572
rect 288390 3093 288450 3571
rect 288387 3092 288453 3093
rect 288387 3028 288388 3092
rect 288452 3028 288453 3092
rect 288387 3027 288453 3028
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 117654 296604 122000
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 121254 300204 122000
rect 318747 122092 318813 122093
rect 318747 122028 318748 122092
rect 318812 122090 318813 122092
rect 319115 122092 319181 122093
rect 319115 122090 319116 122092
rect 318812 122030 319116 122090
rect 318812 122028 318813 122030
rect 318747 122027 318813 122028
rect 319115 122028 319116 122030
rect 319180 122028 319181 122092
rect 319115 122027 319181 122028
rect 301454 121821 301514 121942
rect 301451 121820 301517 121821
rect 301451 121756 301452 121820
rect 301516 121756 301517 121820
rect 301451 121755 301517 121756
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 92454 307404 122000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 310404 96054 311004 122000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 307707 3636 307773 3637
rect 307707 3572 307708 3636
rect 307772 3572 307773 3636
rect 307707 3571 307773 3572
rect 307710 2957 307770 3571
rect 307707 2956 307773 2957
rect 307707 2892 307708 2956
rect 307772 2892 307773 2956
rect 307707 2891 307773 2892
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 99654 314604 122000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 317604 103254 318204 122000
rect 318747 121956 318813 121957
rect 318747 121892 318748 121956
rect 318812 121892 318813 121956
rect 318747 121891 318813 121892
rect 319115 121956 319181 121957
rect 319115 121892 319116 121956
rect 319180 121892 319181 121956
rect 319115 121891 319181 121892
rect 318750 121818 318810 121891
rect 319118 121818 319178 121891
rect 318750 121758 319178 121818
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 317275 3636 317341 3637
rect 317275 3572 317276 3636
rect 317340 3572 317341 3636
rect 317275 3571 317341 3572
rect 317278 2957 317338 3571
rect 317275 2956 317341 2957
rect 317275 2892 317276 2956
rect 317340 2892 317341 2956
rect 317275 2891 317341 2892
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 318750 4390 319178 4450
rect 318750 3909 318810 4390
rect 319118 3909 319178 4390
rect 318747 3908 318813 3909
rect 318747 3844 318748 3908
rect 318812 3844 318813 3908
rect 318747 3843 318813 3844
rect 319115 3908 319181 3909
rect 319115 3844 319116 3908
rect 319180 3844 319181 3908
rect 319115 3843 319181 3844
rect 320038 3773 320098 123659
rect 333835 123452 333901 123453
rect 333835 123388 333836 123452
rect 333900 123388 333901 123452
rect 333835 123387 333901 123388
rect 335307 123452 335373 123453
rect 335307 123388 335308 123452
rect 335372 123450 335373 123452
rect 353155 123452 353221 123453
rect 335372 123390 335554 123450
rect 335372 123388 335373 123390
rect 335307 123387 335373 123388
rect 324267 123316 324333 123317
rect 324267 123252 324268 123316
rect 324332 123252 324333 123316
rect 324267 123251 324333 123252
rect 324270 123045 324330 123251
rect 333838 123045 333898 123387
rect 335494 123317 335554 123390
rect 353155 123388 353156 123452
rect 353220 123388 353221 123452
rect 353155 123387 353221 123388
rect 354627 123452 354693 123453
rect 354627 123388 354628 123452
rect 354692 123450 354693 123452
rect 372475 123452 372541 123453
rect 354692 123390 354874 123450
rect 354692 123388 354693 123390
rect 354627 123387 354693 123388
rect 335491 123316 335557 123317
rect 335491 123252 335492 123316
rect 335556 123252 335557 123316
rect 335491 123251 335557 123252
rect 343587 123316 343653 123317
rect 343587 123252 343588 123316
rect 343652 123252 343653 123316
rect 343587 123251 343653 123252
rect 343590 123045 343650 123251
rect 353158 123045 353218 123387
rect 354814 123317 354874 123390
rect 372475 123388 372476 123452
rect 372540 123388 372541 123452
rect 372475 123387 372541 123388
rect 373947 123452 374013 123453
rect 373947 123388 373948 123452
rect 374012 123450 374013 123452
rect 391795 123452 391861 123453
rect 374012 123390 374194 123450
rect 374012 123388 374013 123390
rect 373947 123387 374013 123388
rect 354811 123316 354877 123317
rect 354811 123252 354812 123316
rect 354876 123252 354877 123316
rect 354811 123251 354877 123252
rect 362907 123316 362973 123317
rect 362907 123252 362908 123316
rect 362972 123252 362973 123316
rect 362907 123251 362973 123252
rect 362910 123045 362970 123251
rect 372478 123045 372538 123387
rect 374134 123317 374194 123390
rect 391795 123388 391796 123452
rect 391860 123388 391861 123452
rect 391795 123387 391861 123388
rect 393267 123452 393333 123453
rect 393267 123388 393268 123452
rect 393332 123450 393333 123452
rect 411115 123452 411181 123453
rect 393332 123390 393514 123450
rect 393332 123388 393333 123390
rect 393267 123387 393333 123388
rect 374131 123316 374197 123317
rect 374131 123252 374132 123316
rect 374196 123252 374197 123316
rect 374131 123251 374197 123252
rect 382227 123316 382293 123317
rect 382227 123252 382228 123316
rect 382292 123252 382293 123316
rect 382227 123251 382293 123252
rect 382230 123045 382290 123251
rect 391798 123045 391858 123387
rect 393454 123317 393514 123390
rect 411115 123388 411116 123452
rect 411180 123388 411181 123452
rect 411115 123387 411181 123388
rect 412587 123452 412653 123453
rect 412587 123388 412588 123452
rect 412652 123450 412653 123452
rect 412652 123390 412834 123450
rect 412652 123388 412653 123390
rect 412587 123387 412653 123388
rect 393451 123316 393517 123317
rect 393451 123252 393452 123316
rect 393516 123252 393517 123316
rect 393451 123251 393517 123252
rect 401547 123316 401613 123317
rect 401547 123252 401548 123316
rect 401612 123252 401613 123316
rect 401547 123251 401613 123252
rect 401550 123045 401610 123251
rect 411118 123045 411178 123387
rect 412774 123317 412834 123390
rect 412771 123316 412837 123317
rect 412771 123252 412772 123316
rect 412836 123252 412837 123316
rect 412771 123251 412837 123252
rect 324267 123044 324333 123045
rect 324267 122980 324268 123044
rect 324332 122980 324333 123044
rect 324267 122979 324333 122980
rect 333835 123044 333901 123045
rect 333835 122980 333836 123044
rect 333900 122980 333901 123044
rect 333835 122979 333901 122980
rect 343587 123044 343653 123045
rect 343587 122980 343588 123044
rect 343652 122980 343653 123044
rect 343587 122979 343653 122980
rect 353155 123044 353221 123045
rect 353155 122980 353156 123044
rect 353220 122980 353221 123044
rect 353155 122979 353221 122980
rect 362907 123044 362973 123045
rect 362907 122980 362908 123044
rect 362972 122980 362973 123044
rect 362907 122979 362973 122980
rect 372475 123044 372541 123045
rect 372475 122980 372476 123044
rect 372540 122980 372541 123044
rect 372475 122979 372541 122980
rect 382227 123044 382293 123045
rect 382227 122980 382228 123044
rect 382292 122980 382293 123044
rect 382227 122979 382293 122980
rect 391795 123044 391861 123045
rect 391795 122980 391796 123044
rect 391860 122980 391861 123044
rect 391795 122979 391861 122980
rect 401547 123044 401613 123045
rect 401547 122980 401548 123044
rect 401612 122980 401613 123044
rect 401547 122979 401613 122980
rect 411115 123044 411181 123045
rect 411115 122980 411116 123044
rect 411180 122980 411181 123044
rect 411115 122979 411181 122980
rect 420134 122909 420194 123302
rect 369899 122908 369965 122909
rect 369899 122844 369900 122908
rect 369964 122844 369965 122908
rect 379283 122908 379349 122909
rect 379283 122858 379284 122908
rect 379348 122858 379349 122908
rect 417555 122908 417621 122909
rect 417555 122858 417556 122908
rect 417620 122858 417621 122908
rect 420131 122908 420197 122909
rect 369899 122843 369965 122844
rect 346350 122710 347146 122770
rect 327027 122228 327093 122229
rect 327027 122164 327028 122228
rect 327092 122164 327093 122228
rect 327027 122163 327093 122164
rect 322614 121821 322674 121942
rect 322611 121820 322677 121821
rect 322611 121756 322612 121820
rect 322676 121756 322677 121820
rect 322611 121755 322677 121756
rect 324804 110454 325404 122000
rect 327030 121685 327090 122163
rect 327027 121684 327093 121685
rect 327027 121620 327028 121684
rect 327092 121620 327093 121684
rect 327027 121619 327093 121620
rect 326846 118693 326906 119902
rect 326843 118692 326909 118693
rect 326843 118628 326844 118692
rect 326908 118628 326909 118692
rect 326843 118627 326909 118628
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 318747 3772 318813 3773
rect 318747 3708 318748 3772
rect 318812 3708 318813 3772
rect 318747 3707 318813 3708
rect 320035 3772 320101 3773
rect 320035 3708 320036 3772
rect 320100 3708 320101 3772
rect 320035 3707 320101 3708
rect 318750 2957 318810 3707
rect 318747 2956 318813 2957
rect 318747 2892 318748 2956
rect 318812 2892 318813 2956
rect 318747 2891 318813 2892
rect 324804 2454 325404 37898
rect 328404 114054 329004 122000
rect 338067 122092 338133 122093
rect 338067 122028 338068 122092
rect 338132 122090 338133 122092
rect 338435 122092 338501 122093
rect 338435 122090 338436 122092
rect 338132 122030 338436 122090
rect 338132 122028 338133 122030
rect 338067 122027 338133 122028
rect 338435 122028 338436 122030
rect 338500 122028 338501 122092
rect 338435 122027 338501 122028
rect 331078 121685 331138 121942
rect 331075 121684 331141 121685
rect 331075 121620 331076 121684
rect 331140 121620 331141 121684
rect 331075 121619 331141 121620
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 327027 3636 327093 3637
rect 327027 3572 327028 3636
rect 327092 3572 327093 3636
rect 327027 3571 327093 3572
rect 327030 2957 327090 3571
rect 327027 2956 327093 2957
rect 327027 2892 327028 2956
rect 327092 2892 327093 2956
rect 327027 2891 327093 2892
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 -2186 329004 5498
rect 332004 117654 332604 122000
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 -4026 332604 9098
rect 335604 121254 336204 122000
rect 338067 121956 338133 121957
rect 338067 121892 338068 121956
rect 338132 121892 338133 121956
rect 338067 121891 338133 121892
rect 338619 121956 338685 121957
rect 338619 121892 338620 121956
rect 338684 121892 338685 121956
rect 338619 121891 338685 121892
rect 338070 121682 338130 121891
rect 338622 121682 338682 121891
rect 338070 121622 338682 121682
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 340643 120052 340709 120053
rect 340643 119988 340644 120052
rect 340708 119988 340709 120052
rect 340643 119987 340709 119988
rect 340646 119458 340706 119987
rect 338067 111484 338133 111485
rect 338067 111420 338068 111484
rect 338132 111420 338133 111484
rect 338067 111419 338133 111420
rect 338070 111213 338130 111419
rect 338067 111212 338133 111213
rect 338067 111148 338068 111212
rect 338132 111148 338133 111212
rect 338067 111147 338133 111148
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 335307 2892 335308 2942
rect 335372 2892 335373 2942
rect 335307 2891 335373 2892
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342302 3773 342362 122622
rect 346350 122229 346410 122710
rect 346347 122228 346413 122229
rect 342804 92454 343404 122000
rect 346347 122164 346348 122228
rect 346412 122164 346413 122228
rect 346347 122163 346413 122164
rect 344878 121685 344938 121942
rect 344875 121684 344941 121685
rect 344875 121620 344876 121684
rect 344940 121620 344941 121684
rect 344875 121619 344941 121620
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342299 3772 342365 3773
rect 342299 3708 342300 3772
rect 342364 3708 342365 3772
rect 342299 3707 342365 3708
rect 340827 2892 340828 2942
rect 340892 2892 340893 2942
rect 340827 2891 340893 2892
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 96054 347004 122000
rect 347086 121685 347146 122710
rect 365667 122228 365733 122229
rect 365667 122164 365668 122228
rect 365732 122164 365733 122228
rect 369902 122178 369962 122843
rect 420131 122844 420132 122908
rect 420196 122844 420197 122908
rect 420131 122843 420197 122844
rect 425099 122908 425165 122909
rect 425099 122844 425100 122908
rect 425164 122844 425165 122908
rect 425099 122843 425165 122844
rect 425102 122178 425162 122843
rect 365667 122163 365733 122164
rect 347083 121684 347149 121685
rect 347083 121620 347084 121684
rect 347148 121620 347149 121684
rect 347083 121619 347149 121620
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 99654 350604 122000
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 103254 354204 122000
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 110454 361404 122000
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 357387 3772 357453 3773
rect 357387 3708 357388 3772
rect 357452 3708 357453 3772
rect 357387 3707 357453 3708
rect 357390 3093 357450 3707
rect 357387 3092 357453 3093
rect 357387 3028 357388 3092
rect 357452 3028 357453 3092
rect 357387 3027 357453 3028
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 114054 365004 122000
rect 365670 121685 365730 122163
rect 365667 121684 365733 121685
rect 365667 121620 365668 121684
rect 365732 121620 365733 121684
rect 365667 121619 365733 121620
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 368004 117654 368604 122000
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 367290 4390 367754 4450
rect 367694 3858 367754 4390
rect 365667 3772 365733 3773
rect 365667 3708 365668 3772
rect 365732 3708 365733 3772
rect 365667 3707 365733 3708
rect 365670 3093 365730 3707
rect 365667 3092 365733 3093
rect 365667 3028 365668 3092
rect 365732 3028 365733 3092
rect 365667 3027 365733 3028
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 121254 372204 122000
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 92454 379404 122000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 382404 96054 383004 122000
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 -3106 383004 23498
rect 386004 99654 386604 122000
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 384987 4180 385053 4181
rect 384987 4116 384988 4180
rect 385052 4116 385053 4180
rect 384987 4115 385053 4116
rect 384990 3637 385050 4115
rect 384987 3636 385053 3637
rect 384987 3572 384988 3636
rect 385052 3572 385053 3636
rect 384987 3571 385053 3572
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 103254 390204 122000
rect 394742 118965 394802 119222
rect 394739 118964 394805 118965
rect 394739 118900 394740 118964
rect 394804 118900 394805 118964
rect 394739 118899 394805 118900
rect 396027 110940 396093 110941
rect 396027 110876 396028 110940
rect 396092 110876 396093 110940
rect 396027 110875 396093 110876
rect 396030 110669 396090 110875
rect 396027 110668 396093 110669
rect 396027 110604 396028 110668
rect 396092 110604 396093 110668
rect 396027 110603 396093 110604
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 110454 397404 122000
rect 398386 122030 399070 122090
rect 399526 118965 399586 119222
rect 399523 118964 399589 118965
rect 399523 118900 399524 118964
rect 399588 118900 399589 118964
rect 399523 118899 399589 118900
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396027 3772 396093 3773
rect 396027 3708 396028 3772
rect 396092 3708 396093 3772
rect 396027 3707 396093 3708
rect 396030 3093 396090 3707
rect 396027 3092 396093 3093
rect 396027 3028 396028 3092
rect 396092 3028 396093 3092
rect 396027 3027 396093 3028
rect 396804 2454 397404 37898
rect 400404 114054 401004 122000
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 398386 3030 398886 3090
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 117654 404604 122000
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 407604 121254 408204 122000
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 408539 120188 408605 120189
rect 408539 120124 408540 120188
rect 408604 120124 408605 120188
rect 408539 120123 408605 120124
rect 408542 119458 408602 120123
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 92454 415404 122000
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 418404 96054 419004 122000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 -3106 419004 23498
rect 422004 99654 422604 122000
rect 422891 120188 422957 120189
rect 422891 120124 422892 120188
rect 422956 120124 422957 120188
rect 422891 120123 422957 120124
rect 422894 119458 422954 120123
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 -4946 422604 27098
rect 425470 3637 425530 123795
rect 434483 122908 434549 122909
rect 434483 122858 434484 122908
rect 434548 122858 434549 122908
rect 444238 122229 444298 122622
rect 434667 122228 434733 122229
rect 434667 122178 434668 122228
rect 434732 122178 434733 122228
rect 444235 122228 444301 122229
rect 425604 103254 426204 122000
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 425467 3636 425533 3637
rect 425467 3572 425468 3636
rect 425532 3572 425533 3636
rect 425467 3571 425533 3572
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 110454 433404 122000
rect 444235 122164 444236 122228
rect 444300 122164 444301 122228
rect 444235 122163 444301 122164
rect 434302 118693 434362 119222
rect 434299 118692 434365 118693
rect 434299 118628 434300 118692
rect 434364 118628 434365 118692
rect 434299 118627 434365 118628
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 436404 114054 437004 122000
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 -2186 437004 5498
rect 440004 117654 440604 122000
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 -4026 440604 9098
rect 443604 121254 444204 122000
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 446627 120188 446693 120189
rect 446627 120138 446628 120188
rect 446692 120138 446693 120188
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 92454 451404 122000
rect 453619 120188 453685 120189
rect 453619 120124 453620 120188
rect 453684 120124 453685 120188
rect 453619 120123 453685 120124
rect 453622 119458 453682 120123
rect 453990 118965 454050 119222
rect 453987 118964 454053 118965
rect 453987 118900 453988 118964
rect 454052 118900 454053 118964
rect 453987 118899 454053 118900
rect 453987 110940 454053 110941
rect 453987 110876 453988 110940
rect 454052 110876 454053 110940
rect 453987 110875 454053 110876
rect 453990 110669 454050 110875
rect 453987 110668 454053 110669
rect 453987 110604 453988 110668
rect 454052 110604 454053 110668
rect 453987 110603 454053 110604
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 444419 4252 444420 4302
rect 444484 4252 444485 4302
rect 444419 4251 444485 4252
rect 450804 -1266 451404 19898
rect 454404 96054 455004 122000
rect 457302 118965 457362 119222
rect 457299 118964 457365 118965
rect 457299 118900 457300 118964
rect 457364 118900 457365 118964
rect 457299 118899 457365 118900
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 451598 2685 451658 2942
rect 451595 2684 451661 2685
rect 451595 2620 451596 2684
rect 451660 2620 451661 2684
rect 451595 2619 451661 2620
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 -3106 455004 23498
rect 458004 99654 458604 122000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 457483 4316 457549 4317
rect 457483 4252 457484 4316
rect 457548 4252 457549 4316
rect 457483 4251 457549 4252
rect 457486 3858 457546 4251
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 -4946 458604 27098
rect 461604 103254 462204 122000
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 461350 2685 461410 2942
rect 461347 2684 461413 2685
rect 461347 2620 461348 2684
rect 461412 2620 461413 2684
rect 461347 2619 461413 2620
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 462454 3773 462514 4302
rect 463558 3773 463618 123931
rect 469259 123452 469325 123453
rect 469259 123388 469260 123452
rect 469324 123450 469325 123452
rect 469324 123390 469506 123450
rect 469324 123388 469325 123390
rect 469259 123387 469325 123388
rect 466315 123252 466316 123302
rect 466380 123252 466381 123302
rect 466315 123251 466381 123252
rect 469446 122909 469506 123390
rect 478643 123452 478709 123453
rect 478643 123388 478644 123452
rect 478708 123388 478709 123452
rect 478643 123387 478709 123388
rect 478275 123316 478341 123317
rect 474043 123252 474044 123302
rect 474108 123252 474109 123302
rect 474043 123251 474109 123252
rect 478275 123252 478276 123316
rect 478340 123252 478341 123316
rect 478275 123251 478341 123252
rect 469443 122908 469509 122909
rect 469443 122844 469444 122908
rect 469508 122844 469509 122908
rect 469443 122843 469509 122844
rect 478278 122229 478338 123251
rect 478646 122909 478706 123387
rect 478643 122908 478709 122909
rect 478643 122844 478644 122908
rect 478708 122844 478709 122908
rect 478643 122843 478709 122844
rect 486555 122908 486621 122909
rect 486555 122844 486556 122908
rect 486620 122844 486621 122908
rect 486555 122843 486621 122844
rect 478275 122228 478341 122229
rect 478275 122164 478276 122228
rect 478340 122164 478341 122228
rect 478275 122163 478341 122164
rect 478643 122228 478709 122229
rect 478643 122164 478644 122228
rect 478708 122164 478709 122228
rect 478643 122163 478709 122164
rect 468804 110454 469404 122000
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 462451 3772 462517 3773
rect 462451 3708 462452 3772
rect 462516 3708 462517 3772
rect 462451 3707 462517 3708
rect 463555 3772 463621 3773
rect 463555 3708 463556 3772
rect 463620 3708 463621 3772
rect 463555 3707 463621 3708
rect 468804 2454 469404 37898
rect 472404 114054 473004 122000
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 476004 117654 476604 122000
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 473307 111484 473373 111485
rect 473307 111420 473308 111484
rect 473372 111420 473373 111484
rect 473307 111419 473373 111420
rect 473310 111213 473370 111419
rect 473307 111212 473373 111213
rect 473307 111148 473308 111212
rect 473372 111148 473373 111212
rect 473307 111147 473373 111148
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 470550 2549 470610 2942
rect 470547 2548 470613 2549
rect 470547 2484 470548 2548
rect 470612 2484 470613 2548
rect 470547 2483 470613 2484
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 478646 3773 478706 122163
rect 479604 121254 480204 122000
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 479379 4180 479445 4181
rect 479379 4116 479380 4180
rect 479444 4116 479445 4180
rect 479379 4115 479445 4116
rect 478643 3772 478709 3773
rect 478643 3708 478644 3772
rect 478708 3708 478709 3772
rect 478643 3707 478709 3708
rect 479382 2549 479442 4115
rect 479379 2548 479445 2549
rect 479379 2484 479380 2548
rect 479444 2484 479445 2548
rect 479379 2483 479445 2484
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 485635 4180 485701 4181
rect 485635 4116 485636 4180
rect 485700 4116 485701 4180
rect 485635 4115 485701 4116
rect 485638 3178 485698 4115
rect 486558 2821 486618 122843
rect 491894 122229 491954 123931
rect 493179 123860 493245 123861
rect 493179 123796 493180 123860
rect 493244 123796 493245 123860
rect 493179 123795 493245 123796
rect 493182 123181 493242 123795
rect 493363 123452 493429 123453
rect 493363 123388 493364 123452
rect 493428 123388 493429 123452
rect 493363 123387 493429 123388
rect 493179 123180 493245 123181
rect 493179 123116 493180 123180
rect 493244 123116 493245 123180
rect 493179 123115 493245 123116
rect 493366 123045 493426 123387
rect 493363 123044 493429 123045
rect 493363 122980 493364 123044
rect 493428 122980 493429 123044
rect 493363 122979 493429 122980
rect 491891 122228 491957 122229
rect 491891 122164 491892 122228
rect 491956 122164 491957 122228
rect 491891 122163 491957 122164
rect 486804 92454 487404 122000
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486555 2820 486621 2821
rect 486555 2756 486556 2820
rect 486620 2756 486621 2820
rect 486555 2755 486621 2756
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 96054 491004 122000
rect 493550 117197 493610 123931
rect 497227 123860 497293 123861
rect 497227 123796 497228 123860
rect 497292 123796 497293 123860
rect 497227 123795 497293 123796
rect 497230 123538 497290 123795
rect 495387 122228 495453 122229
rect 495387 122164 495388 122228
rect 495452 122164 495453 122228
rect 495387 122163 495453 122164
rect 493547 117196 493613 117197
rect 493547 117132 493548 117196
rect 493612 117132 493613 117196
rect 493547 117131 493613 117132
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 99654 494604 122000
rect 495390 121141 495450 122163
rect 495387 121140 495453 121141
rect 495387 121076 495388 121140
rect 495452 121076 495453 121140
rect 495387 121075 495453 121076
rect 495942 121005 496002 122622
rect 496494 121141 496554 123302
rect 497598 122770 497658 194022
rect 497966 190090 498026 194790
rect 498150 194170 498210 195470
rect 498150 194110 498394 194170
rect 496678 122710 497658 122770
rect 497782 190030 498026 190090
rect 496491 121140 496557 121141
rect 496491 121076 496492 121140
rect 496556 121076 496557 121140
rect 496491 121075 496557 121076
rect 495939 121004 496005 121005
rect 495939 120940 495940 121004
rect 496004 120940 496005 121004
rect 495939 120939 496005 120940
rect 495939 118284 496005 118285
rect 495939 118220 495940 118284
rect 496004 118220 496005 118284
rect 495939 118219 496005 118220
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 495206 3773 495266 4302
rect 495387 3908 495453 3909
rect 495387 3844 495388 3908
rect 495452 3844 495453 3908
rect 495387 3843 495453 3844
rect 495203 3772 495269 3773
rect 495203 3708 495204 3772
rect 495268 3708 495269 3772
rect 495390 3770 495450 3843
rect 495942 3770 496002 118219
rect 496678 115290 496738 122710
rect 497782 122362 497842 190030
rect 498334 189410 498394 194110
rect 497966 189350 498394 189410
rect 497966 187370 498026 189350
rect 498518 188050 498578 195382
rect 498886 189410 498946 198870
rect 498334 187990 498578 188050
rect 498702 189350 498946 189410
rect 497966 187310 498210 187370
rect 498150 183970 498210 187310
rect 497966 183910 498210 183970
rect 497966 168330 498026 183910
rect 498334 183378 498394 187990
rect 498702 180570 498762 189350
rect 499070 188730 499130 199278
rect 499254 191178 499314 199414
rect 499438 191314 499498 202270
rect 500174 202058 500234 202270
rect 499622 201998 500234 202058
rect 499622 199338 499682 201998
rect 499622 199278 500234 199338
rect 499806 196346 499866 198782
rect 500174 196978 500234 199278
rect 500726 199018 500786 202950
rect 501646 202197 501706 237491
rect 501830 237285 501890 237627
rect 501827 237284 501893 237285
rect 501827 237220 501828 237284
rect 501892 237220 501893 237284
rect 501827 237219 501893 237220
rect 502014 233205 502074 244155
rect 502011 233204 502077 233205
rect 502011 233140 502012 233204
rect 502076 233140 502077 233204
rect 502011 233139 502077 233140
rect 502198 232250 502258 244699
rect 501830 232190 502258 232250
rect 501830 226810 501890 232190
rect 502382 231845 502442 503643
rect 502379 231844 502445 231845
rect 502379 231780 502380 231844
rect 502444 231780 502445 231844
rect 502379 231779 502445 231780
rect 501830 226750 502074 226810
rect 501827 226676 501893 226677
rect 501827 226612 501828 226676
rect 501892 226612 501893 226676
rect 501827 226611 501893 226612
rect 501830 221509 501890 226611
rect 502014 221509 502074 226750
rect 502198 226677 502258 231422
rect 502379 231300 502445 231301
rect 502379 231236 502380 231300
rect 502444 231236 502445 231300
rect 502379 231235 502445 231236
rect 502195 226676 502261 226677
rect 502195 226612 502196 226676
rect 502260 226612 502261 226676
rect 502195 226611 502261 226612
rect 502195 226540 502261 226541
rect 502195 226476 502196 226540
rect 502260 226476 502261 226540
rect 502195 226475 502261 226476
rect 501827 221508 501893 221509
rect 501827 221444 501828 221508
rect 501892 221444 501893 221508
rect 501827 221443 501893 221444
rect 502011 221508 502077 221509
rect 502011 221444 502012 221508
rect 502076 221444 502077 221508
rect 502011 221443 502077 221444
rect 502198 220013 502258 226475
rect 501827 220012 501893 220013
rect 501827 219948 501828 220012
rect 501892 219948 501893 220012
rect 501827 219947 501893 219948
rect 502195 220012 502261 220013
rect 502195 219948 502196 220012
rect 502260 219948 502261 220012
rect 502195 219947 502261 219948
rect 501643 202196 501709 202197
rect 501094 202058 501154 202182
rect 501643 202132 501644 202196
rect 501708 202132 501709 202196
rect 501643 202131 501709 202132
rect 501094 201998 501522 202058
rect 501462 201245 501522 201998
rect 501459 201244 501525 201245
rect 501459 201180 501460 201244
rect 501524 201180 501525 201244
rect 501459 201179 501525 201180
rect 501275 200428 501341 200429
rect 501275 200364 501276 200428
rect 501340 200364 501341 200428
rect 501275 200363 501341 200364
rect 501278 196618 501338 200363
rect 501830 199610 501890 219947
rect 502195 219876 502261 219877
rect 502195 219812 502196 219876
rect 502260 219812 502261 219876
rect 502195 219811 502261 219812
rect 502011 216340 502077 216341
rect 502011 216276 502012 216340
rect 502076 216276 502077 216340
rect 502011 216275 502077 216276
rect 502014 209269 502074 216275
rect 502198 215797 502258 219811
rect 502195 215796 502261 215797
rect 502195 215732 502196 215796
rect 502260 215732 502261 215796
rect 502195 215731 502261 215732
rect 502195 211852 502261 211853
rect 502195 211850 502196 211852
rect 502152 211788 502196 211850
rect 502260 211788 502261 211852
rect 502152 211787 502261 211788
rect 502011 209268 502077 209269
rect 502011 209204 502012 209268
rect 502076 209204 502077 209268
rect 502011 209203 502077 209204
rect 502152 209130 502212 211787
rect 502014 209070 502212 209130
rect 502014 204098 502074 209070
rect 502149 204100 502215 204101
rect 502149 204098 502150 204100
rect 502014 204038 502150 204098
rect 502149 204036 502150 204038
rect 502214 204036 502215 204100
rect 502149 204035 502215 204036
rect 502011 203284 502077 203285
rect 502011 203220 502012 203284
rect 502076 203220 502077 203284
rect 502011 203219 502077 203220
rect 502014 200429 502074 203219
rect 502195 202196 502261 202197
rect 502195 202132 502196 202196
rect 502260 202132 502261 202196
rect 502195 202131 502261 202132
rect 502011 200428 502077 200429
rect 502011 200364 502012 200428
rect 502076 200364 502077 200428
rect 502011 200363 502077 200364
rect 501462 199550 501890 199610
rect 501462 196757 501522 199550
rect 501643 199476 501709 199477
rect 501643 199412 501644 199476
rect 501708 199412 501709 199476
rect 501643 199411 501709 199412
rect 501459 196756 501525 196757
rect 501459 196692 501460 196756
rect 501524 196692 501525 196756
rect 501459 196691 501525 196692
rect 499622 196286 499866 196346
rect 500174 196558 501338 196618
rect 499622 192130 499682 196286
rect 500174 195618 500234 196558
rect 501459 196348 501525 196349
rect 501459 196284 501460 196348
rect 501524 196284 501525 196348
rect 501459 196283 501525 196284
rect 501275 196212 501341 196213
rect 501275 196210 501276 196212
rect 500726 196150 501276 196210
rect 500726 194850 500786 196150
rect 501275 196148 501276 196150
rect 501340 196148 501341 196212
rect 501275 196147 501341 196148
rect 501462 195805 501522 196283
rect 501459 195804 501525 195805
rect 501459 195740 501460 195804
rect 501524 195740 501525 195804
rect 501459 195739 501525 195740
rect 501646 195666 501706 199411
rect 501827 198116 501893 198117
rect 501827 198052 501828 198116
rect 501892 198052 501893 198116
rect 501827 198051 501893 198052
rect 500174 194790 500786 194850
rect 500910 195606 501706 195666
rect 500174 194258 500234 194790
rect 500910 192946 500970 195606
rect 501459 195532 501525 195533
rect 501459 195530 501460 195532
rect 501094 195470 501460 195530
rect 501094 193082 501154 195470
rect 501459 195468 501460 195470
rect 501524 195468 501525 195532
rect 501459 195467 501525 195468
rect 501462 194445 501522 194702
rect 501459 194444 501525 194445
rect 501459 194380 501460 194444
rect 501524 194380 501525 194444
rect 501459 194379 501525 194380
rect 501462 193221 501522 194022
rect 501459 193220 501525 193221
rect 501459 193156 501460 193220
rect 501524 193156 501525 193220
rect 501459 193155 501525 193156
rect 501094 193022 501706 193082
rect 500910 192886 501522 192946
rect 499622 192070 500602 192130
rect 499438 191302 499902 191314
rect 499438 191254 500050 191302
rect 500542 191178 500602 192070
rect 501275 191452 501341 191453
rect 501275 191450 501276 191452
rect 499254 191118 499498 191178
rect 499438 191042 499498 191118
rect 499990 191118 500602 191178
rect 500910 191390 501276 191450
rect 499438 190982 499866 191042
rect 499438 190090 499498 190622
rect 498334 180510 498762 180570
rect 498886 188670 499130 188730
rect 499254 190030 499498 190090
rect 498334 173090 498394 180510
rect 498886 179978 498946 188670
rect 499254 179890 499314 190030
rect 499806 189410 499866 190982
rect 499438 189350 499866 189410
rect 499438 183562 499498 189350
rect 499990 183698 500050 191118
rect 499990 183638 500602 183698
rect 499438 183502 500418 183562
rect 499254 179830 499498 179890
rect 499438 178938 499498 179830
rect 499070 178878 499498 178938
rect 499070 178618 499130 178878
rect 499806 178258 499866 183142
rect 500358 182610 500418 183502
rect 498518 178198 499866 178258
rect 499990 182550 500418 182610
rect 499990 178258 500050 182550
rect 500542 178618 500602 183638
rect 500910 178394 500970 191390
rect 501275 191388 501276 191390
rect 501340 191388 501341 191452
rect 501275 191387 501341 191388
rect 501275 191316 501341 191317
rect 501275 191252 501276 191316
rect 501340 191252 501341 191316
rect 501275 191251 501341 191252
rect 501278 190090 501338 191251
rect 501462 191181 501522 192886
rect 501646 191317 501706 193022
rect 501643 191316 501709 191317
rect 501643 191252 501644 191316
rect 501708 191252 501709 191316
rect 501643 191251 501709 191252
rect 501459 191180 501525 191181
rect 501459 191116 501460 191180
rect 501524 191116 501525 191180
rect 501459 191115 501525 191116
rect 501643 191180 501709 191181
rect 501643 191116 501644 191180
rect 501708 191116 501709 191180
rect 501643 191115 501709 191116
rect 501459 191044 501525 191045
rect 501459 190980 501460 191044
rect 501524 190980 501525 191044
rect 501459 190979 501525 190980
rect 501094 190030 501338 190090
rect 501094 178530 501154 190030
rect 501275 189820 501341 189821
rect 501275 189756 501276 189820
rect 501340 189756 501341 189820
rect 501275 189755 501341 189756
rect 501278 186285 501338 189755
rect 501275 186284 501341 186285
rect 501275 186220 501276 186284
rect 501340 186220 501341 186284
rect 501275 186219 501341 186220
rect 501462 184789 501522 190979
rect 501646 184789 501706 191115
rect 501830 184789 501890 198051
rect 502011 197436 502077 197437
rect 502011 197372 502012 197436
rect 502076 197372 502077 197436
rect 502011 197371 502077 197372
rect 502014 196893 502074 197371
rect 502011 196892 502077 196893
rect 502011 196828 502012 196892
rect 502076 196828 502077 196892
rect 502011 196827 502077 196828
rect 502011 196756 502077 196757
rect 502011 196692 502012 196756
rect 502076 196692 502077 196756
rect 502011 196691 502077 196692
rect 502014 191045 502074 196691
rect 502198 191181 502258 202131
rect 502195 191180 502261 191181
rect 502195 191116 502196 191180
rect 502260 191116 502261 191180
rect 502195 191115 502261 191116
rect 502011 191044 502077 191045
rect 502011 190980 502012 191044
rect 502076 190980 502077 191044
rect 502011 190979 502077 190980
rect 502011 190908 502077 190909
rect 502011 190844 502012 190908
rect 502076 190844 502077 190908
rect 502011 190843 502077 190844
rect 502014 186965 502074 190843
rect 502195 190772 502261 190773
rect 502195 190708 502196 190772
rect 502260 190708 502261 190772
rect 502195 190707 502261 190708
rect 502011 186964 502077 186965
rect 502011 186900 502012 186964
rect 502076 186900 502077 186964
rect 502011 186899 502077 186900
rect 502198 186690 502258 190707
rect 502014 186630 502258 186690
rect 502014 184789 502074 186630
rect 502195 186420 502261 186421
rect 502195 186356 502196 186420
rect 502260 186356 502261 186420
rect 502195 186355 502261 186356
rect 501459 184788 501525 184789
rect 501459 184724 501460 184788
rect 501524 184724 501525 184788
rect 501459 184723 501525 184724
rect 501643 184788 501709 184789
rect 501643 184724 501644 184788
rect 501708 184724 501709 184788
rect 501643 184723 501709 184724
rect 501827 184788 501893 184789
rect 501827 184724 501828 184788
rect 501892 184724 501893 184788
rect 501827 184723 501893 184724
rect 502011 184788 502077 184789
rect 502011 184724 502012 184788
rect 502076 184724 502077 184788
rect 502011 184723 502077 184724
rect 501827 184516 501893 184517
rect 501827 184452 501828 184516
rect 501892 184452 501893 184516
rect 501827 184451 501893 184452
rect 502011 184516 502077 184517
rect 502011 184452 502012 184516
rect 502076 184452 502077 184516
rect 502011 184451 502077 184452
rect 501275 184380 501341 184381
rect 501275 184316 501276 184380
rect 501340 184316 501341 184380
rect 501275 184315 501341 184316
rect 501459 184380 501525 184381
rect 501459 184316 501460 184380
rect 501524 184316 501525 184380
rect 501459 184315 501525 184316
rect 501643 184380 501709 184381
rect 501643 184316 501644 184380
rect 501708 184316 501709 184380
rect 501643 184315 501709 184316
rect 501278 181930 501338 184315
rect 501462 182341 501522 184315
rect 501459 182340 501525 182341
rect 501459 182276 501460 182340
rect 501524 182276 501525 182340
rect 501459 182275 501525 182276
rect 501459 181932 501525 181933
rect 501459 181930 501460 181932
rect 501278 181870 501460 181930
rect 501459 181868 501460 181870
rect 501524 181868 501525 181932
rect 501459 181867 501525 181868
rect 501459 181796 501525 181797
rect 501459 181732 501460 181796
rect 501524 181732 501525 181796
rect 501459 181731 501525 181732
rect 501462 181250 501522 181731
rect 501278 181190 501522 181250
rect 501278 179213 501338 181190
rect 501459 180028 501525 180029
rect 501459 179964 501460 180028
rect 501524 179964 501525 180028
rect 501459 179963 501525 179964
rect 501275 179212 501341 179213
rect 501275 179148 501276 179212
rect 501340 179148 501341 179212
rect 501275 179147 501341 179148
rect 501275 178532 501341 178533
rect 501275 178530 501276 178532
rect 501094 178470 501276 178530
rect 501275 178468 501276 178470
rect 501340 178468 501341 178532
rect 501275 178467 501341 178468
rect 501462 178397 501522 179963
rect 501459 178396 501525 178397
rect 500910 178334 501154 178394
rect 501094 178258 501154 178334
rect 501459 178332 501460 178396
rect 501524 178332 501525 178396
rect 501459 178331 501525 178332
rect 501459 178260 501525 178261
rect 501459 178258 501460 178260
rect 499990 178198 500418 178258
rect 501094 178198 501460 178258
rect 498518 176490 498578 178198
rect 500358 177850 500418 178198
rect 501459 178196 501460 178198
rect 501524 178196 501525 178260
rect 501459 178195 501525 178196
rect 501459 178124 501525 178125
rect 501459 178060 501460 178124
rect 501524 178060 501525 178124
rect 501459 178059 501525 178060
rect 500358 177790 500786 177850
rect 498518 176430 499498 176490
rect 498702 173226 498762 173622
rect 498702 173166 498946 173226
rect 498334 173030 498762 173090
rect 498334 169098 498394 172262
rect 497966 168270 498578 168330
rect 498150 164250 498210 166822
rect 497966 164190 498210 164250
rect 497966 154050 498026 164190
rect 498518 162346 498578 168270
rect 498150 162286 498578 162346
rect 498150 154730 498210 162286
rect 498702 161802 498762 173030
rect 498886 170234 498946 173166
rect 499070 171050 499130 175662
rect 499438 172498 499498 176430
rect 499070 170990 499498 171050
rect 499438 170594 499498 170990
rect 498886 170174 499682 170234
rect 499254 168330 499314 168862
rect 498886 168270 499314 168330
rect 498886 162346 498946 168270
rect 499622 167650 499682 170174
rect 499070 167590 499682 167650
rect 499070 162482 499130 167590
rect 499806 165698 499866 177702
rect 499990 177258 500418 177306
rect 499990 177246 500270 177258
rect 499990 169010 500050 177246
rect 500726 176898 500786 177790
rect 501462 177173 501522 178059
rect 501459 177172 501525 177173
rect 501459 177108 501460 177172
rect 501524 177108 501525 177172
rect 501459 177107 501525 177108
rect 501459 177036 501525 177037
rect 501459 176972 501460 177036
rect 501524 176972 501525 177036
rect 501459 176971 501525 176972
rect 500358 176838 500786 176898
rect 500358 173858 500418 176838
rect 501275 175812 501341 175813
rect 501275 175810 501276 175812
rect 500726 175750 501276 175810
rect 500726 170370 500786 175750
rect 501275 175748 501276 175750
rect 501340 175748 501341 175812
rect 501275 175747 501341 175748
rect 501275 175676 501341 175677
rect 501275 175612 501276 175676
rect 501340 175612 501341 175676
rect 501275 175611 501341 175612
rect 501278 173090 501338 175611
rect 500542 170310 500786 170370
rect 501094 173030 501338 173090
rect 500542 170234 500602 170310
rect 500358 170174 500602 170234
rect 499990 168950 500234 169010
rect 499438 162482 499498 162742
rect 499070 162422 499498 162482
rect 498886 162286 500050 162346
rect 499990 161802 500050 162286
rect 498334 161742 498762 161802
rect 499070 161742 500050 161802
rect 498334 160850 498394 161742
rect 498334 160790 498946 160850
rect 498150 154670 498578 154730
rect 497966 153990 498210 154050
rect 498150 148698 498210 153990
rect 498518 148018 498578 154670
rect 498886 147522 498946 160790
rect 499070 149970 499130 161742
rect 500174 161394 500234 168950
rect 500358 162210 500418 170174
rect 500726 167058 500786 169542
rect 500726 162346 500786 165462
rect 501094 162890 501154 173030
rect 501275 172412 501341 172413
rect 501275 172348 501276 172412
rect 501340 172348 501341 172412
rect 501275 172347 501341 172348
rect 501278 163706 501338 172347
rect 501462 163845 501522 176971
rect 501646 173365 501706 184315
rect 501643 173364 501709 173365
rect 501643 173300 501644 173364
rect 501708 173300 501709 173364
rect 501643 173299 501709 173300
rect 501643 173228 501709 173229
rect 501643 173164 501644 173228
rect 501708 173164 501709 173228
rect 501643 173163 501709 173164
rect 501646 171050 501706 173163
rect 501830 171189 501890 184451
rect 502014 183565 502074 184451
rect 502198 183837 502258 186355
rect 502195 183836 502261 183837
rect 502195 183772 502196 183836
rect 502260 183772 502261 183836
rect 502195 183771 502261 183772
rect 502195 183700 502261 183701
rect 502195 183636 502196 183700
rect 502260 183636 502261 183700
rect 502195 183635 502261 183636
rect 502011 183564 502077 183565
rect 502011 183500 502012 183564
rect 502076 183500 502077 183564
rect 502011 183499 502077 183500
rect 502011 182340 502077 182341
rect 502011 182276 502012 182340
rect 502076 182276 502077 182340
rect 502011 182275 502077 182276
rect 502014 177309 502074 182275
rect 502198 182069 502258 183635
rect 502195 182068 502261 182069
rect 502195 182004 502196 182068
rect 502260 182004 502261 182068
rect 502195 182003 502261 182004
rect 502195 181932 502261 181933
rect 502195 181868 502196 181932
rect 502260 181868 502261 181932
rect 502195 181867 502261 181868
rect 502198 180165 502258 181867
rect 502195 180164 502261 180165
rect 502195 180100 502196 180164
rect 502260 180100 502261 180164
rect 502195 180099 502261 180100
rect 502195 178940 502261 178941
rect 502195 178876 502196 178940
rect 502260 178876 502261 178940
rect 502195 178875 502261 178876
rect 502011 177308 502077 177309
rect 502011 177244 502012 177308
rect 502076 177244 502077 177308
rect 502011 177243 502077 177244
rect 502011 177172 502077 177173
rect 502011 177108 502012 177172
rect 502076 177108 502077 177172
rect 502011 177107 502077 177108
rect 502014 175677 502074 177107
rect 502011 175676 502077 175677
rect 502011 175612 502012 175676
rect 502076 175612 502077 175676
rect 502011 175611 502077 175612
rect 502198 175541 502258 178875
rect 502011 175540 502077 175541
rect 502011 175476 502012 175540
rect 502076 175476 502077 175540
rect 502011 175475 502077 175476
rect 502195 175540 502261 175541
rect 502195 175476 502196 175540
rect 502260 175476 502261 175540
rect 502195 175475 502261 175476
rect 501827 171188 501893 171189
rect 501827 171124 501828 171188
rect 501892 171124 501893 171188
rect 501827 171123 501893 171124
rect 501646 170990 501890 171050
rect 501643 170508 501709 170509
rect 501643 170444 501644 170508
rect 501708 170444 501709 170508
rect 501643 170443 501709 170444
rect 501459 163844 501525 163845
rect 501459 163780 501460 163844
rect 501524 163780 501525 163844
rect 501459 163779 501525 163780
rect 501459 163708 501525 163709
rect 501459 163706 501460 163708
rect 501278 163646 501460 163706
rect 501459 163644 501460 163646
rect 501524 163644 501525 163708
rect 501459 163643 501525 163644
rect 501459 162892 501525 162893
rect 501459 162890 501460 162892
rect 501094 162830 501460 162890
rect 501459 162828 501460 162830
rect 501524 162828 501525 162892
rect 501459 162827 501525 162828
rect 501459 162484 501525 162485
rect 501459 162420 501460 162484
rect 501524 162420 501525 162484
rect 501459 162419 501525 162420
rect 501462 162346 501522 162419
rect 501646 162349 501706 170443
rect 501830 166429 501890 170990
rect 502014 170509 502074 175475
rect 502195 175404 502261 175405
rect 502195 175340 502196 175404
rect 502260 175340 502261 175404
rect 502195 175339 502261 175340
rect 502198 174045 502258 175339
rect 502195 174044 502261 174045
rect 502195 173980 502196 174044
rect 502260 173980 502261 174044
rect 502195 173979 502261 173980
rect 502195 173092 502261 173093
rect 502195 173028 502196 173092
rect 502260 173028 502261 173092
rect 502195 173027 502261 173028
rect 502011 170508 502077 170509
rect 502011 170444 502012 170508
rect 502076 170444 502077 170508
rect 502011 170443 502077 170444
rect 502198 170370 502258 173027
rect 502014 170310 502258 170370
rect 501827 166428 501893 166429
rect 501827 166364 501828 166428
rect 501892 166364 501893 166428
rect 501827 166363 501893 166364
rect 502014 166021 502074 170310
rect 502195 170236 502261 170237
rect 502195 170172 502196 170236
rect 502260 170172 502261 170236
rect 502195 170171 502261 170172
rect 501827 166020 501893 166021
rect 501827 165956 501828 166020
rect 501892 165956 501893 166020
rect 501827 165955 501893 165956
rect 502011 166020 502077 166021
rect 502011 165956 502012 166020
rect 502076 165956 502077 166020
rect 502011 165955 502077 165956
rect 500726 162286 501522 162346
rect 501643 162348 501709 162349
rect 501643 162284 501644 162348
rect 501708 162284 501709 162348
rect 501643 162283 501709 162284
rect 500358 162150 501522 162210
rect 501275 161804 501341 161805
rect 501275 161740 501276 161804
rect 501340 161740 501341 161804
rect 501275 161739 501341 161740
rect 501278 161397 501338 161739
rect 499438 161334 500234 161394
rect 501275 161396 501341 161397
rect 499438 150738 499498 161334
rect 501275 161332 501276 161396
rect 501340 161332 501341 161396
rect 501275 161331 501341 161332
rect 499806 156178 499866 160702
rect 501275 157996 501341 157997
rect 501275 157932 501276 157996
rect 501340 157932 501341 157996
rect 501275 157931 501341 157932
rect 501278 157450 501338 157931
rect 500174 157390 501338 157450
rect 499070 149910 499314 149970
rect 499254 148970 499314 149910
rect 499806 148610 499866 155262
rect 500174 152690 500234 157390
rect 501462 156770 501522 162150
rect 501643 160852 501709 160853
rect 501643 160788 501644 160852
rect 501708 160788 501709 160852
rect 501643 160787 501709 160788
rect 501646 158810 501706 160787
rect 501830 158949 501890 165955
rect 502011 165884 502077 165885
rect 502011 165820 502012 165884
rect 502076 165820 502077 165884
rect 502011 165819 502077 165820
rect 502014 160853 502074 165819
rect 502011 160852 502077 160853
rect 502011 160788 502012 160852
rect 502076 160788 502077 160852
rect 502011 160787 502077 160788
rect 501827 158948 501893 158949
rect 501827 158884 501828 158948
rect 501892 158884 501893 158948
rect 501827 158883 501893 158884
rect 502011 158812 502077 158813
rect 501646 158750 501890 158810
rect 501643 157452 501709 157453
rect 501643 157388 501644 157452
rect 501708 157388 501709 157452
rect 501643 157387 501709 157388
rect 501278 156710 501522 156770
rect 500174 152630 500418 152690
rect 500358 151330 500418 152630
rect 500358 151270 500970 151330
rect 500358 149970 500418 150502
rect 500358 149910 500786 149970
rect 497966 147462 498946 147522
rect 499070 148550 499866 148610
rect 497966 136642 498026 147462
rect 498334 146842 498394 147102
rect 498334 146782 498762 146842
rect 498334 143850 498394 145062
rect 498702 144618 498762 146782
rect 498334 143790 498578 143850
rect 498518 139906 498578 143790
rect 499070 140538 499130 148550
rect 499438 145298 499498 147782
rect 499990 145298 500050 147102
rect 500358 145890 500418 148462
rect 500726 146026 500786 149910
rect 500910 147930 500970 151270
rect 501278 148610 501338 156710
rect 501459 156636 501525 156637
rect 501459 156572 501460 156636
rect 501524 156572 501525 156636
rect 501459 156571 501525 156572
rect 501462 152149 501522 156571
rect 501459 152148 501525 152149
rect 501459 152084 501460 152148
rect 501524 152084 501525 152148
rect 501459 152083 501525 152084
rect 501459 150924 501525 150925
rect 501459 150860 501460 150924
rect 501524 150860 501525 150924
rect 501459 150859 501525 150860
rect 501462 148885 501522 150859
rect 501459 148884 501525 148885
rect 501459 148820 501460 148884
rect 501524 148820 501525 148884
rect 501459 148819 501525 148820
rect 501459 148612 501525 148613
rect 501459 148610 501460 148612
rect 501278 148550 501460 148610
rect 501459 148548 501460 148550
rect 501524 148548 501525 148612
rect 501459 148547 501525 148548
rect 500910 147870 501338 147930
rect 501278 147525 501338 147870
rect 501275 147524 501341 147525
rect 501275 147460 501276 147524
rect 501340 147460 501341 147524
rect 501275 147459 501341 147460
rect 501459 147252 501525 147253
rect 501459 147250 501460 147252
rect 501242 147190 501460 147250
rect 501459 147188 501460 147190
rect 501524 147188 501525 147252
rect 501459 147187 501525 147188
rect 501459 146028 501525 146029
rect 501459 146026 501460 146028
rect 500726 145966 501460 146026
rect 501459 145964 501460 145966
rect 501524 145964 501525 146028
rect 501459 145963 501525 145964
rect 501459 145892 501525 145893
rect 500358 145830 501338 145890
rect 499448 145150 499498 145298
rect 498518 139846 499130 139906
rect 499070 137322 499130 139846
rect 498886 137262 499130 137322
rect 497966 136582 498578 136642
rect 498518 133738 498578 136582
rect 498150 130250 498210 132822
rect 497966 130190 498210 130250
rect 497966 123997 498026 130190
rect 497963 123996 498029 123997
rect 497963 123932 497964 123996
rect 498028 123932 498029 123996
rect 497963 123931 498029 123932
rect 498331 123996 498397 123997
rect 498331 123932 498332 123996
rect 498396 123932 498397 123996
rect 498331 123931 498397 123932
rect 497230 122302 497842 122362
rect 496678 115230 496922 115290
rect 496862 102237 496922 115230
rect 496859 102236 496925 102237
rect 496859 102172 496860 102236
rect 496924 102172 496925 102236
rect 496859 102171 496925 102172
rect 497043 102236 497109 102237
rect 497043 102172 497044 102236
rect 497108 102172 497109 102236
rect 497043 102171 497109 102172
rect 497046 26349 497106 102171
rect 497230 101690 497290 122302
rect 497411 122228 497477 122229
rect 497411 122164 497412 122228
rect 497476 122164 497477 122228
rect 497411 122163 497477 122164
rect 497414 118965 497474 122163
rect 497411 118964 497477 118965
rect 497411 118900 497412 118964
rect 497476 118900 497477 118964
rect 497411 118899 497477 118900
rect 497604 103254 498204 122000
rect 498334 121005 498394 123931
rect 498518 123589 498578 130782
rect 498886 123994 498946 137262
rect 499438 137050 499498 140302
rect 499990 140178 500050 144382
rect 500726 143986 500786 145062
rect 500174 143926 500786 143986
rect 500174 140450 500234 143926
rect 501278 140589 501338 145830
rect 501459 145828 501460 145892
rect 501524 145828 501525 145892
rect 501459 145827 501525 145828
rect 501275 140588 501341 140589
rect 501275 140524 501276 140588
rect 501340 140524 501341 140588
rect 501275 140523 501341 140524
rect 501275 140452 501341 140453
rect 501275 140450 501276 140452
rect 500174 140390 501276 140450
rect 501275 140388 501276 140390
rect 501340 140388 501341 140452
rect 501275 140387 501341 140388
rect 501275 140316 501341 140317
rect 501275 140252 501276 140316
rect 501340 140252 501341 140316
rect 501275 140251 501341 140252
rect 501278 140178 501338 140251
rect 501462 140181 501522 145827
rect 499990 140118 501338 140178
rect 501459 140180 501525 140181
rect 501459 140116 501460 140180
rect 501524 140116 501525 140180
rect 501459 140115 501525 140116
rect 501459 138684 501525 138685
rect 501459 138682 501460 138684
rect 499070 136990 499498 137050
rect 499622 138622 501460 138682
rect 499070 123997 499130 136990
rect 499254 134418 499314 136222
rect 499254 131018 499314 133502
rect 499622 129978 499682 138622
rect 501459 138620 501460 138622
rect 501524 138620 501525 138684
rect 501459 138619 501525 138620
rect 501459 138548 501525 138549
rect 501459 138546 501460 138548
rect 500542 138486 501460 138546
rect 499990 131018 500050 136902
rect 500542 132290 500602 138486
rect 501459 138484 501460 138486
rect 501524 138484 501525 138548
rect 501459 138483 501525 138484
rect 501459 138412 501525 138413
rect 501459 138410 501460 138412
rect 500910 138350 501460 138410
rect 500910 136458 500970 138350
rect 501459 138348 501460 138350
rect 501524 138348 501525 138412
rect 501459 138347 501525 138348
rect 501646 137869 501706 157387
rect 501830 140045 501890 158750
rect 502011 158748 502012 158812
rect 502076 158748 502077 158812
rect 502011 158747 502077 158748
rect 501827 140044 501893 140045
rect 501827 139980 501828 140044
rect 501892 139980 501893 140044
rect 501827 139979 501893 139980
rect 501827 139908 501893 139909
rect 501827 139844 501828 139908
rect 501892 139844 501893 139908
rect 501827 139843 501893 139844
rect 501830 138685 501890 139843
rect 501827 138684 501893 138685
rect 501827 138620 501828 138684
rect 501892 138620 501893 138684
rect 501827 138619 501893 138620
rect 502014 138005 502074 158747
rect 502198 155685 502258 170171
rect 502195 155684 502261 155685
rect 502195 155620 502196 155684
rect 502260 155620 502261 155684
rect 502195 155619 502261 155620
rect 502195 155276 502261 155277
rect 502195 155212 502196 155276
rect 502260 155212 502261 155276
rect 502195 155211 502261 155212
rect 502011 138004 502077 138005
rect 502011 137940 502012 138004
rect 502076 137940 502077 138004
rect 502011 137939 502077 137940
rect 501643 137868 501709 137869
rect 501643 137804 501644 137868
rect 501708 137804 501709 137868
rect 501643 137803 501709 137804
rect 502011 137732 502077 137733
rect 502011 137668 502012 137732
rect 502076 137668 502077 137732
rect 502011 137667 502077 137668
rect 501275 136780 501341 136781
rect 501275 136716 501276 136780
rect 501340 136716 501341 136780
rect 501275 136715 501341 136716
rect 501278 135690 501338 136715
rect 501827 136644 501893 136645
rect 501827 136580 501828 136644
rect 501892 136580 501893 136644
rect 501827 136579 501893 136580
rect 501459 136372 501525 136373
rect 501459 136308 501460 136372
rect 501524 136308 501525 136372
rect 501459 136307 501525 136308
rect 501094 135630 501338 135690
rect 500542 132230 500786 132290
rect 500726 131610 500786 132230
rect 500542 131550 500786 131610
rect 499622 129918 500418 129978
rect 498702 123934 498946 123994
rect 499067 123996 499133 123997
rect 498515 123588 498581 123589
rect 498515 123524 498516 123588
rect 498580 123524 498581 123588
rect 498515 123523 498581 123524
rect 498702 123450 498762 123934
rect 499067 123932 499068 123996
rect 499132 123932 499133 123996
rect 499067 123931 499133 123932
rect 499438 123861 499498 129422
rect 499619 123996 499685 123997
rect 499619 123932 499620 123996
rect 499684 123932 499685 123996
rect 499619 123931 499685 123932
rect 499435 123860 499501 123861
rect 499435 123796 499436 123860
rect 499500 123796 499501 123860
rect 499435 123795 499501 123796
rect 499435 123724 499501 123725
rect 499435 123722 499436 123724
rect 498518 123390 498762 123450
rect 499254 123662 499436 123722
rect 498518 121005 498578 123390
rect 499254 121682 499314 123662
rect 499435 123660 499436 123662
rect 499500 123660 499501 123724
rect 499435 123659 499501 123660
rect 499435 123180 499501 123181
rect 499435 123116 499436 123180
rect 499500 123116 499501 123180
rect 499435 123115 499501 123116
rect 499116 121622 499314 121682
rect 498331 121004 498397 121005
rect 498331 120940 498332 121004
rect 498396 120940 498397 121004
rect 498331 120939 498397 120940
rect 498515 121004 498581 121005
rect 498515 120940 498516 121004
rect 498580 120940 498581 121004
rect 499116 121002 499176 121622
rect 499438 121413 499498 123115
rect 499435 121412 499501 121413
rect 499435 121348 499436 121412
rect 499500 121348 499501 121412
rect 499435 121347 499501 121348
rect 499116 120942 499314 121002
rect 498515 120939 498581 120940
rect 498515 120596 498581 120597
rect 498515 120532 498516 120596
rect 498580 120532 498581 120596
rect 498515 120531 498581 120532
rect 498331 116788 498397 116789
rect 498331 116724 498332 116788
rect 498396 116724 498397 116788
rect 498331 116723 498397 116724
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497230 101630 497474 101690
rect 497043 26348 497109 26349
rect 497043 26284 497044 26348
rect 497108 26284 497109 26348
rect 497043 26283 497109 26284
rect 496859 26076 496925 26077
rect 496859 26012 496860 26076
rect 496924 26012 496925 26076
rect 496859 26011 496925 26012
rect 496862 6765 496922 26011
rect 496859 6764 496925 6765
rect 496859 6700 496860 6764
rect 496924 6700 496925 6764
rect 496859 6699 496925 6700
rect 497414 6493 497474 101630
rect 497604 67254 498204 102698
rect 498334 73130 498394 116723
rect 498518 106997 498578 120531
rect 498699 120324 498765 120325
rect 498699 120260 498700 120324
rect 498764 120260 498765 120324
rect 498699 120259 498765 120260
rect 498515 106996 498581 106997
rect 498515 106932 498516 106996
rect 498580 106932 498581 106996
rect 498515 106931 498581 106932
rect 498334 73070 498578 73130
rect 498518 67557 498578 73070
rect 498515 67556 498581 67557
rect 498515 67492 498516 67556
rect 498580 67492 498581 67556
rect 498515 67491 498581 67492
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 498331 62796 498397 62797
rect 498331 62732 498332 62796
rect 498396 62732 498397 62796
rect 498331 62731 498397 62732
rect 498334 57901 498394 62731
rect 498331 57900 498397 57901
rect 498331 57836 498332 57900
rect 498396 57836 498397 57900
rect 498331 57835 498397 57836
rect 498515 48380 498581 48381
rect 498515 48316 498516 48380
rect 498580 48316 498581 48380
rect 498515 48315 498581 48316
rect 498518 44437 498578 48315
rect 498515 44436 498581 44437
rect 498515 44372 498516 44436
rect 498580 44372 498581 44436
rect 498515 44371 498581 44372
rect 498331 44300 498397 44301
rect 498331 44236 498332 44300
rect 498396 44236 498397 44300
rect 498331 44235 498397 44236
rect 498334 34373 498394 44235
rect 498331 34372 498397 34373
rect 498331 34308 498332 34372
rect 498396 34308 498397 34372
rect 498331 34307 498397 34308
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 497411 6492 497477 6493
rect 497411 6428 497412 6492
rect 497476 6428 497477 6492
rect 497411 6427 497477 6428
rect 495390 3710 495634 3770
rect 495203 3707 495269 3708
rect 495574 3637 495634 3710
rect 495758 3710 496002 3770
rect 495387 3636 495453 3637
rect 495387 3572 495388 3636
rect 495452 3572 495453 3636
rect 495387 3571 495453 3572
rect 495571 3636 495637 3637
rect 495571 3572 495572 3636
rect 495636 3572 495637 3636
rect 495571 3571 495637 3572
rect 495390 3090 495450 3571
rect 495758 3229 495818 3710
rect 495755 3228 495821 3229
rect 495755 3164 495756 3228
rect 495820 3164 495821 3228
rect 495755 3163 495821 3164
rect 496123 3092 496189 3093
rect 496123 3090 496124 3092
rect 495390 3030 496124 3090
rect 496123 3028 496124 3030
rect 496188 3028 496189 3092
rect 496123 3027 496189 3028
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 498331 24988 498397 24989
rect 498331 24924 498332 24988
rect 498396 24924 498397 24988
rect 498331 24923 498397 24924
rect 498334 15333 498394 24923
rect 498331 15332 498397 15333
rect 498331 15268 498332 15332
rect 498396 15268 498397 15332
rect 498331 15267 498397 15268
rect 498515 9756 498581 9757
rect 498515 9692 498516 9756
rect 498580 9692 498581 9756
rect 498515 9691 498581 9692
rect 498518 5813 498578 9691
rect 498515 5812 498581 5813
rect 498515 5748 498516 5812
rect 498580 5748 498581 5812
rect 498515 5747 498581 5748
rect 498331 5676 498397 5677
rect 498331 5612 498332 5676
rect 498396 5612 498397 5676
rect 498331 5611 498397 5612
rect 498334 3365 498394 5611
rect 498331 3364 498397 3365
rect 498331 3300 498332 3364
rect 498396 3300 498397 3364
rect 498331 3299 498397 3300
rect 498702 3178 498762 120259
rect 499067 116108 499133 116109
rect 499067 116044 499068 116108
rect 499132 116044 499133 116108
rect 499067 116043 499133 116044
rect 498883 104548 498949 104549
rect 498883 104484 498884 104548
rect 498948 104484 498949 104548
rect 498883 104483 498949 104484
rect 498886 19005 498946 104483
rect 498883 19004 498949 19005
rect 498883 18940 498884 19004
rect 498948 18940 498949 19004
rect 498883 18939 498949 18940
rect 499070 3229 499130 116043
rect 499254 104549 499314 120942
rect 499622 120325 499682 123931
rect 499803 123588 499869 123589
rect 499803 123524 499804 123588
rect 499868 123524 499869 123588
rect 499803 123523 499869 123524
rect 499806 123181 499866 123523
rect 499803 123180 499869 123181
rect 499803 123116 499804 123180
rect 499868 123116 499869 123180
rect 499803 123115 499869 123116
rect 500358 122637 500418 129918
rect 500542 123586 500602 131550
rect 501094 130930 501154 135630
rect 501462 135149 501522 136307
rect 501459 135148 501525 135149
rect 501459 135084 501460 135148
rect 501524 135084 501525 135148
rect 501459 135083 501525 135084
rect 501459 134876 501525 134877
rect 501459 134812 501460 134876
rect 501524 134812 501525 134876
rect 501459 134811 501525 134812
rect 501643 134876 501709 134877
rect 501643 134812 501644 134876
rect 501708 134812 501709 134876
rect 501643 134811 501709 134812
rect 501275 133516 501341 133517
rect 501275 133452 501276 133516
rect 501340 133452 501341 133516
rect 501275 133451 501341 133452
rect 501278 130933 501338 133451
rect 500726 130870 501154 130930
rect 501275 130932 501341 130933
rect 500726 123997 500786 130870
rect 501275 130868 501276 130932
rect 501340 130868 501341 130932
rect 501275 130867 501341 130868
rect 501275 126172 501341 126173
rect 501275 126170 501276 126172
rect 501094 126110 501276 126170
rect 500723 123996 500789 123997
rect 500723 123932 500724 123996
rect 500788 123932 500789 123996
rect 500723 123931 500789 123932
rect 500907 123724 500973 123725
rect 500907 123660 500908 123724
rect 500972 123660 500973 123724
rect 500907 123659 500973 123660
rect 500542 123526 500786 123586
rect 500539 123452 500605 123453
rect 500539 123388 500540 123452
rect 500604 123388 500605 123452
rect 500539 123387 500605 123388
rect 500355 122636 500421 122637
rect 500355 122572 500356 122636
rect 500420 122572 500421 122636
rect 500355 122571 500421 122572
rect 499619 120324 499685 120325
rect 499619 120260 499620 120324
rect 499684 120260 499685 120324
rect 499619 120259 499685 120260
rect 499987 120324 500053 120325
rect 499987 120260 499988 120324
rect 500052 120260 500053 120324
rect 499987 120259 500053 120260
rect 499803 118012 499869 118013
rect 499803 117948 499804 118012
rect 499868 117948 499869 118012
rect 499803 117947 499869 117948
rect 499435 106996 499501 106997
rect 499435 106932 499436 106996
rect 499500 106932 499501 106996
rect 499435 106931 499501 106932
rect 499251 104548 499317 104549
rect 499251 104484 499252 104548
rect 499316 104484 499317 104548
rect 499251 104483 499317 104484
rect 499438 92445 499498 106931
rect 499435 92444 499501 92445
rect 499435 92380 499436 92444
rect 499500 92380 499501 92444
rect 499435 92379 499501 92380
rect 499251 92308 499317 92309
rect 499251 92244 499252 92308
rect 499316 92244 499317 92308
rect 499251 92243 499317 92244
rect 499254 72997 499314 92243
rect 499251 72996 499317 72997
rect 499251 72932 499252 72996
rect 499316 72932 499317 72996
rect 499251 72931 499317 72932
rect 499435 55316 499501 55317
rect 499435 55252 499436 55316
rect 499500 55252 499501 55316
rect 499435 55251 499501 55252
rect 499438 37365 499498 55251
rect 499435 37364 499501 37365
rect 499435 37300 499436 37364
rect 499500 37300 499501 37364
rect 499435 37299 499501 37300
rect 499619 37092 499685 37093
rect 499619 37028 499620 37092
rect 499684 37028 499685 37092
rect 499619 37027 499685 37028
rect 499622 18733 499682 37027
rect 499619 18732 499685 18733
rect 499619 18668 499620 18732
rect 499684 18668 499685 18732
rect 499619 18667 499685 18668
rect 499806 3501 499866 117947
rect 499990 95165 500050 120259
rect 500355 114612 500421 114613
rect 500355 114548 500356 114612
rect 500420 114548 500421 114612
rect 500355 114547 500421 114548
rect 500171 113252 500237 113253
rect 500171 113188 500172 113252
rect 500236 113188 500237 113252
rect 500171 113187 500237 113188
rect 500174 109717 500234 113187
rect 500171 109716 500237 109717
rect 500171 109652 500172 109716
rect 500236 109652 500237 109716
rect 500171 109651 500237 109652
rect 500358 104821 500418 114547
rect 500355 104820 500421 104821
rect 500355 104756 500356 104820
rect 500420 104756 500421 104820
rect 500355 104755 500421 104756
rect 500171 96796 500237 96797
rect 500171 96732 500172 96796
rect 500236 96732 500237 96796
rect 500171 96731 500237 96732
rect 499987 95164 500053 95165
rect 499987 95100 499988 95164
rect 500052 95100 500053 95164
rect 499987 95099 500053 95100
rect 499987 56676 500053 56677
rect 499987 56612 499988 56676
rect 500052 56612 500053 56676
rect 499987 56611 500053 56612
rect 499990 49061 500050 56611
rect 499987 49060 500053 49061
rect 499987 48996 499988 49060
rect 500052 48996 500053 49060
rect 499987 48995 500053 48996
rect 499987 38724 500053 38725
rect 499987 38660 499988 38724
rect 500052 38660 500053 38724
rect 499987 38659 500053 38660
rect 499990 29749 500050 38659
rect 499987 29748 500053 29749
rect 499987 29684 499988 29748
rect 500052 29684 500053 29748
rect 499987 29683 500053 29684
rect 500174 4045 500234 96731
rect 500542 92853 500602 123387
rect 500726 123317 500786 123526
rect 500723 123316 500789 123317
rect 500723 123252 500724 123316
rect 500788 123252 500789 123316
rect 500723 123251 500789 123252
rect 500910 123178 500970 123659
rect 500726 123118 500970 123178
rect 500726 123045 500786 123118
rect 500723 123044 500789 123045
rect 500723 122980 500724 123044
rect 500788 122980 500789 123044
rect 500723 122979 500789 122980
rect 501094 121005 501154 126110
rect 501275 126108 501276 126110
rect 501340 126108 501341 126172
rect 501275 126107 501341 126108
rect 501275 123860 501341 123861
rect 501275 123796 501276 123860
rect 501340 123796 501341 123860
rect 501275 123795 501341 123796
rect 501091 121004 501157 121005
rect 501091 120940 501092 121004
rect 501156 120940 501157 121004
rect 501091 120939 501157 120940
rect 501091 120732 501157 120733
rect 501091 120668 501092 120732
rect 501156 120668 501157 120732
rect 501091 120667 501157 120668
rect 500723 116244 500789 116245
rect 500723 116180 500724 116244
rect 500788 116180 500789 116244
rect 500723 116179 500789 116180
rect 500539 92852 500605 92853
rect 500539 92788 500540 92852
rect 500604 92788 500605 92852
rect 500539 92787 500605 92788
rect 500726 92717 500786 116179
rect 501094 111349 501154 120667
rect 501278 115429 501338 123795
rect 501462 121141 501522 134811
rect 501459 121140 501525 121141
rect 501459 121076 501460 121140
rect 501524 121076 501525 121140
rect 501459 121075 501525 121076
rect 501646 120869 501706 134811
rect 501643 120868 501709 120869
rect 501643 120804 501644 120868
rect 501708 120804 501709 120868
rect 501643 120803 501709 120804
rect 501830 116650 501890 136579
rect 501646 116590 501890 116650
rect 501275 115428 501341 115429
rect 501275 115364 501276 115428
rect 501340 115364 501341 115428
rect 501275 115363 501341 115364
rect 501091 111348 501157 111349
rect 501091 111284 501092 111348
rect 501156 111284 501157 111348
rect 501091 111283 501157 111284
rect 500723 92716 500789 92717
rect 500723 92652 500724 92716
rect 500788 92652 500789 92716
rect 500723 92651 500789 92652
rect 500539 91764 500605 91765
rect 500539 91700 500540 91764
rect 500604 91700 500605 91764
rect 500539 91699 500605 91700
rect 500355 82924 500421 82925
rect 500355 82860 500356 82924
rect 500420 82860 500421 82924
rect 500355 82859 500421 82860
rect 500358 77213 500418 82859
rect 500355 77212 500421 77213
rect 500355 77148 500356 77212
rect 500420 77148 500421 77212
rect 500355 77147 500421 77148
rect 500355 68372 500421 68373
rect 500355 68308 500356 68372
rect 500420 68308 500421 68372
rect 500355 68307 500421 68308
rect 500358 49061 500418 68307
rect 500542 56541 500602 91699
rect 501091 87004 501157 87005
rect 501091 86940 501092 87004
rect 501156 86940 501157 87004
rect 501091 86939 501157 86940
rect 501094 83061 501154 86939
rect 501091 83060 501157 83061
rect 501091 82996 501092 83060
rect 501156 82996 501157 83060
rect 501091 82995 501157 82996
rect 501646 60757 501706 116590
rect 501643 60756 501709 60757
rect 501643 60692 501644 60756
rect 501708 60692 501709 60756
rect 501643 60691 501709 60692
rect 501827 60756 501893 60757
rect 501827 60692 501828 60756
rect 501892 60692 501893 60756
rect 501827 60691 501893 60692
rect 500539 56540 500605 56541
rect 500539 56476 500540 56540
rect 500604 56476 500605 56540
rect 500539 56475 500605 56476
rect 500355 49060 500421 49061
rect 500355 48996 500356 49060
rect 500420 48996 500421 49060
rect 500355 48995 500421 48996
rect 500539 48924 500605 48925
rect 500539 48860 500540 48924
rect 500604 48860 500605 48924
rect 500539 48859 500605 48860
rect 500542 37229 500602 48859
rect 500539 37228 500605 37229
rect 500539 37164 500540 37228
rect 500604 37164 500605 37228
rect 500539 37163 500605 37164
rect 500355 29748 500421 29749
rect 500355 29684 500356 29748
rect 500420 29684 500421 29748
rect 500355 29683 500421 29684
rect 500539 29748 500605 29749
rect 500539 29684 500540 29748
rect 500604 29684 500605 29748
rect 500539 29683 500605 29684
rect 500358 8941 500418 29683
rect 500542 16013 500602 29683
rect 501830 29610 501890 60691
rect 501462 29550 501890 29610
rect 501462 21994 501522 29550
rect 501462 21934 501706 21994
rect 500539 16012 500605 16013
rect 500539 15948 500540 16012
rect 500604 15948 500605 16012
rect 500539 15947 500605 15948
rect 500355 8940 500421 8941
rect 500355 8876 500356 8940
rect 500420 8876 500421 8940
rect 500355 8875 500421 8876
rect 500171 4044 500237 4045
rect 500171 3980 500172 4044
rect 500236 3980 500237 4044
rect 500171 3979 500237 3980
rect 499803 3500 499869 3501
rect 499803 3436 499804 3500
rect 499868 3436 499869 3500
rect 499803 3435 499869 3436
rect 499067 3228 499133 3229
rect 499067 3164 499068 3228
rect 499132 3164 499133 3228
rect 499067 3163 499133 3164
rect 501646 3093 501706 21934
rect 502014 3909 502074 137667
rect 502198 125085 502258 155211
rect 502195 125084 502261 125085
rect 502195 125020 502196 125084
rect 502260 125020 502261 125084
rect 502195 125019 502261 125020
rect 502195 124948 502261 124949
rect 502195 124884 502196 124948
rect 502260 124884 502261 124948
rect 502195 124883 502261 124884
rect 502198 4997 502258 124883
rect 502382 16285 502442 231235
rect 502566 84829 502626 542267
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 502931 531452 502997 531453
rect 502931 531388 502932 531452
rect 502996 531388 502997 531452
rect 502931 531387 502997 531388
rect 502747 461276 502813 461277
rect 502747 461212 502748 461276
rect 502812 461212 502813 461276
rect 502747 461211 502813 461212
rect 502563 84828 502629 84829
rect 502563 84764 502564 84828
rect 502628 84764 502629 84828
rect 502563 84763 502629 84764
rect 502379 16284 502445 16285
rect 502379 16220 502380 16284
rect 502444 16220 502445 16284
rect 502379 16219 502445 16220
rect 502750 14653 502810 461211
rect 502934 121685 502994 531387
rect 504219 507244 504285 507245
rect 504219 507180 504220 507244
rect 504284 507180 504285 507244
rect 504219 507179 504285 507180
rect 503667 475420 503733 475421
rect 503667 475356 503668 475420
rect 503732 475356 503733 475420
rect 503667 475355 503733 475356
rect 503670 454018 503730 475355
rect 503667 450668 503733 450669
rect 503667 450604 503668 450668
rect 503732 450604 503733 450668
rect 503667 450603 503733 450604
rect 503299 394364 503365 394365
rect 503299 394300 503300 394364
rect 503364 394300 503365 394364
rect 503299 394299 503365 394300
rect 503302 388738 503362 394299
rect 503299 388380 503365 388381
rect 503299 388316 503300 388380
rect 503364 388316 503365 388380
rect 503299 388315 503365 388316
rect 503302 385338 503362 388315
rect 503115 355740 503181 355741
rect 503115 355676 503116 355740
rect 503180 355676 503181 355740
rect 503115 355675 503181 355676
rect 502931 121684 502997 121685
rect 502931 121620 502932 121684
rect 502996 121620 502997 121684
rect 502931 121619 502997 121620
rect 503118 16421 503178 355675
rect 503299 313308 503365 313309
rect 503299 313244 503300 313308
rect 503364 313244 503365 313308
rect 503299 313243 503365 313244
rect 503115 16420 503181 16421
rect 503115 16356 503116 16420
rect 503180 16356 503181 16420
rect 503115 16355 503181 16356
rect 502747 14652 502813 14653
rect 502747 14588 502748 14652
rect 502812 14588 502813 14652
rect 502747 14587 502813 14588
rect 502195 4996 502261 4997
rect 502195 4932 502196 4996
rect 502260 4932 502261 4996
rect 502195 4931 502261 4932
rect 503302 4861 503362 313243
rect 503483 249796 503549 249797
rect 503483 249732 503484 249796
rect 503548 249732 503549 249796
rect 503483 249731 503549 249732
rect 503486 242181 503546 249731
rect 503483 242180 503549 242181
rect 503483 242116 503484 242180
rect 503548 242116 503549 242180
rect 503483 242115 503549 242116
rect 503483 242044 503549 242045
rect 503483 241980 503484 242044
rect 503548 241980 503549 242044
rect 503483 241979 503549 241980
rect 503486 235653 503546 241979
rect 503483 235652 503549 235653
rect 503483 235588 503484 235652
rect 503548 235588 503549 235652
rect 503483 235587 503549 235588
rect 503483 229124 503549 229125
rect 503483 229060 503484 229124
rect 503548 229060 503549 229124
rect 503483 229059 503549 229060
rect 503486 193085 503546 229059
rect 503483 193084 503549 193085
rect 503483 193020 503484 193084
rect 503548 193020 503549 193084
rect 503483 193019 503549 193020
rect 503483 192948 503549 192949
rect 503483 192884 503484 192948
rect 503548 192884 503549 192948
rect 503483 192883 503549 192884
rect 503486 190909 503546 192883
rect 503483 190908 503549 190909
rect 503483 190844 503484 190908
rect 503548 190844 503549 190908
rect 503483 190843 503549 190844
rect 503483 186964 503549 186965
rect 503483 186900 503484 186964
rect 503548 186900 503549 186964
rect 503483 186899 503549 186900
rect 503486 183701 503546 186899
rect 503483 183700 503549 183701
rect 503483 183636 503484 183700
rect 503548 183636 503549 183700
rect 503483 183635 503549 183636
rect 503483 180164 503549 180165
rect 503483 180100 503484 180164
rect 503548 180100 503549 180164
rect 503483 180099 503549 180100
rect 503486 165069 503546 180099
rect 503483 165068 503549 165069
rect 503483 165004 503484 165068
rect 503548 165004 503549 165068
rect 503483 165003 503549 165004
rect 503483 164932 503549 164933
rect 503483 164868 503484 164932
rect 503548 164868 503549 164932
rect 503483 164867 503549 164868
rect 503486 155821 503546 164867
rect 503483 155820 503549 155821
rect 503483 155756 503484 155820
rect 503548 155756 503549 155820
rect 503483 155755 503549 155756
rect 503483 155684 503549 155685
rect 503483 155620 503484 155684
rect 503548 155620 503549 155684
rect 503483 155619 503549 155620
rect 503486 146981 503546 155619
rect 503483 146980 503549 146981
rect 503483 146916 503484 146980
rect 503548 146916 503549 146980
rect 503483 146915 503549 146916
rect 503483 143988 503549 143989
rect 503483 143924 503484 143988
rect 503548 143924 503549 143988
rect 503483 143923 503549 143924
rect 503486 138821 503546 143923
rect 503483 138820 503549 138821
rect 503483 138756 503484 138820
rect 503548 138756 503549 138820
rect 503483 138755 503549 138756
rect 503483 138684 503549 138685
rect 503483 138620 503484 138684
rect 503548 138620 503549 138684
rect 503483 138619 503549 138620
rect 503486 125221 503546 138619
rect 503483 125220 503549 125221
rect 503483 125156 503484 125220
rect 503548 125156 503549 125220
rect 503483 125155 503549 125156
rect 503483 124948 503549 124949
rect 503483 124884 503484 124948
rect 503548 124884 503549 124948
rect 503483 124883 503549 124884
rect 503486 116245 503546 124883
rect 503483 116244 503549 116245
rect 503483 116180 503484 116244
rect 503548 116180 503549 116244
rect 503483 116179 503549 116180
rect 503670 17509 503730 450603
rect 504222 427957 504282 507179
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504587 447132 504653 447133
rect 504587 447068 504588 447132
rect 504652 447068 504653 447132
rect 504587 447067 504653 447068
rect 504219 427956 504285 427957
rect 504219 427892 504220 427956
rect 504284 427892 504285 427956
rect 504219 427891 504285 427892
rect 504219 427684 504285 427685
rect 504219 427620 504220 427684
rect 504284 427620 504285 427684
rect 504219 427619 504285 427620
rect 504035 408644 504101 408645
rect 504035 408580 504036 408644
rect 504100 408580 504101 408644
rect 504035 408579 504101 408580
rect 503851 408508 503917 408509
rect 503851 408444 503852 408508
rect 503916 408444 503917 408508
rect 503851 408443 503917 408444
rect 503667 17508 503733 17509
rect 503667 17444 503668 17508
rect 503732 17444 503733 17508
rect 503667 17443 503733 17444
rect 503854 17373 503914 408443
rect 504038 398853 504098 408579
rect 504035 398852 504101 398853
rect 504035 398788 504036 398852
rect 504100 398788 504101 398852
rect 504035 398787 504101 398788
rect 504035 387292 504101 387293
rect 504035 387228 504036 387292
rect 504100 387228 504101 387292
rect 504035 387227 504101 387228
rect 504038 349621 504098 387227
rect 504035 349620 504101 349621
rect 504035 349556 504036 349620
rect 504100 349556 504101 349620
rect 504035 349555 504101 349556
rect 504035 339012 504101 339013
rect 504035 338948 504036 339012
rect 504100 338948 504101 339012
rect 504035 338947 504101 338948
rect 504038 326365 504098 338947
rect 504035 326364 504101 326365
rect 504035 326300 504036 326364
rect 504100 326300 504101 326364
rect 504035 326299 504101 326300
rect 504035 326228 504101 326229
rect 504035 326164 504036 326228
rect 504100 326164 504101 326228
rect 504035 326163 504101 326164
rect 504038 316709 504098 326163
rect 504035 316708 504101 316709
rect 504035 316644 504036 316708
rect 504100 316644 504101 316708
rect 504035 316643 504101 316644
rect 504035 316572 504101 316573
rect 504035 316508 504036 316572
rect 504100 316508 504101 316572
rect 504035 316507 504101 316508
rect 504038 307053 504098 316507
rect 504035 307052 504101 307053
rect 504035 306988 504036 307052
rect 504100 306988 504101 307052
rect 504035 306987 504101 306988
rect 504035 297532 504101 297533
rect 504035 297468 504036 297532
rect 504100 297468 504101 297532
rect 504035 297467 504101 297468
rect 504038 287061 504098 297467
rect 504222 290189 504282 427619
rect 504403 425100 504469 425101
rect 504403 425036 504404 425100
rect 504468 425036 504469 425100
rect 504403 425035 504469 425036
rect 504406 408645 504466 425035
rect 504403 408644 504469 408645
rect 504403 408580 504404 408644
rect 504468 408580 504469 408644
rect 504403 408579 504469 408580
rect 504403 398716 504469 398717
rect 504403 398652 504404 398716
rect 504468 398652 504469 398716
rect 504403 398651 504469 398652
rect 504406 347717 504466 398651
rect 504590 349893 504650 447067
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504587 349892 504653 349893
rect 504587 349828 504588 349892
rect 504652 349828 504653 349892
rect 504587 349827 504653 349828
rect 504587 349620 504653 349621
rect 504587 349556 504588 349620
rect 504652 349556 504653 349620
rect 504587 349555 504653 349556
rect 504403 347716 504469 347717
rect 504403 347652 504404 347716
rect 504468 347652 504469 347716
rect 504403 347651 504469 347652
rect 504590 339013 504650 349555
rect 504587 339012 504653 339013
rect 504587 338948 504588 339012
rect 504652 338948 504653 339012
rect 504587 338947 504653 338948
rect 504587 338876 504653 338877
rect 504587 338812 504588 338876
rect 504652 338812 504653 338876
rect 504587 338811 504653 338812
rect 504590 326501 504650 338811
rect 504587 326500 504653 326501
rect 504587 326436 504588 326500
rect 504652 326436 504653 326500
rect 504587 326435 504653 326436
rect 504804 326454 505404 361898
rect 504587 326364 504653 326365
rect 504587 326300 504588 326364
rect 504652 326300 504653 326364
rect 504587 326299 504653 326300
rect 504590 316845 504650 326299
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504587 316844 504653 316845
rect 504587 316780 504588 316844
rect 504652 316780 504653 316844
rect 504587 316779 504653 316780
rect 504587 316708 504653 316709
rect 504587 316644 504588 316708
rect 504652 316644 504653 316708
rect 504587 316643 504653 316644
rect 504590 307189 504650 316643
rect 504587 307188 504653 307189
rect 504587 307124 504588 307188
rect 504652 307124 504653 307188
rect 504587 307123 504653 307124
rect 504587 307052 504653 307053
rect 504587 306988 504588 307052
rect 504652 306988 504653 307052
rect 504587 306987 504653 306988
rect 504590 297533 504650 306987
rect 504587 297532 504653 297533
rect 504587 297468 504588 297532
rect 504652 297468 504653 297532
rect 504587 297467 504653 297468
rect 504403 297396 504469 297397
rect 504403 297332 504404 297396
rect 504468 297332 504469 297396
rect 504403 297331 504469 297332
rect 504406 290730 504466 297331
rect 504406 290670 504650 290730
rect 504219 290188 504285 290189
rect 504219 290124 504220 290188
rect 504284 290124 504285 290188
rect 504219 290123 504285 290124
rect 504035 287060 504101 287061
rect 504035 286996 504036 287060
rect 504100 286996 504101 287060
rect 504035 286995 504101 286996
rect 504219 287060 504285 287061
rect 504219 286996 504220 287060
rect 504284 286996 504285 287060
rect 504219 286995 504285 286996
rect 504035 251972 504101 251973
rect 504035 251908 504036 251972
rect 504100 251908 504101 251972
rect 504035 251907 504101 251908
rect 504038 246125 504098 251907
rect 504222 249797 504282 286995
rect 504590 271829 504650 290670
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504587 271828 504653 271829
rect 504587 271764 504588 271828
rect 504652 271764 504653 271828
rect 504587 271763 504653 271764
rect 504587 267068 504653 267069
rect 504587 267004 504588 267068
rect 504652 267004 504653 267068
rect 504587 267003 504653 267004
rect 504219 249796 504285 249797
rect 504219 249732 504220 249796
rect 504284 249732 504285 249796
rect 504219 249731 504285 249732
rect 504403 249660 504469 249661
rect 504403 249596 504404 249660
rect 504468 249596 504469 249660
rect 504403 249595 504469 249596
rect 504219 246532 504285 246533
rect 504219 246468 504220 246532
rect 504284 246468 504285 246532
rect 504219 246467 504285 246468
rect 504035 246124 504101 246125
rect 504035 246060 504036 246124
rect 504100 246060 504101 246124
rect 504035 246059 504101 246060
rect 504035 242180 504101 242181
rect 504035 242116 504036 242180
rect 504100 242116 504101 242180
rect 504035 242115 504101 242116
rect 504038 235381 504098 242115
rect 504035 235380 504101 235381
rect 504035 235316 504036 235380
rect 504100 235316 504101 235380
rect 504035 235315 504101 235316
rect 504035 222052 504101 222053
rect 504035 221988 504036 222052
rect 504100 221988 504101 222052
rect 504035 221987 504101 221988
rect 504038 214573 504098 221987
rect 504035 214572 504101 214573
rect 504035 214508 504036 214572
rect 504100 214508 504101 214572
rect 504035 214507 504101 214508
rect 504035 210764 504101 210765
rect 504035 210700 504036 210764
rect 504100 210700 504101 210764
rect 504035 210699 504101 210700
rect 504038 199477 504098 210699
rect 504035 199476 504101 199477
rect 504035 199412 504036 199476
rect 504100 199412 504101 199476
rect 504035 199411 504101 199412
rect 504035 199340 504101 199341
rect 504035 199276 504036 199340
rect 504100 199276 504101 199340
rect 504035 199275 504101 199276
rect 504038 192949 504098 199275
rect 504035 192948 504101 192949
rect 504035 192884 504036 192948
rect 504100 192884 504101 192948
rect 504035 192883 504101 192884
rect 504222 186829 504282 246467
rect 504406 239053 504466 249595
rect 504403 239052 504469 239053
rect 504403 238988 504404 239052
rect 504468 238988 504469 239052
rect 504403 238987 504469 238988
rect 504590 235517 504650 267003
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504587 235516 504653 235517
rect 504587 235452 504588 235516
rect 504652 235452 504653 235516
rect 504587 235451 504653 235452
rect 504587 235380 504653 235381
rect 504587 235316 504588 235380
rect 504652 235316 504653 235380
rect 504587 235315 504653 235316
rect 504403 222052 504469 222053
rect 504403 221988 504404 222052
rect 504468 222050 504469 222052
rect 504590 222050 504650 235315
rect 504468 221990 504650 222050
rect 504468 221988 504469 221990
rect 504403 221987 504469 221988
rect 504587 221916 504653 221917
rect 504587 221852 504588 221916
rect 504652 221852 504653 221916
rect 504587 221851 504653 221852
rect 504590 219418 504650 221851
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504403 214572 504469 214573
rect 504403 214508 504404 214572
rect 504468 214508 504469 214572
rect 504403 214507 504469 214508
rect 504219 186828 504285 186829
rect 504219 186764 504220 186828
rect 504284 186764 504285 186828
rect 504219 186763 504285 186764
rect 504406 186010 504466 214507
rect 504590 211581 504650 215102
rect 504587 211580 504653 211581
rect 504587 211516 504588 211580
rect 504652 211516 504653 211580
rect 504587 211515 504653 211516
rect 504587 203420 504653 203421
rect 504587 203356 504588 203420
rect 504652 203356 504653 203420
rect 504587 203355 504653 203356
rect 504590 196349 504650 203355
rect 504587 196348 504653 196349
rect 504587 196284 504588 196348
rect 504652 196284 504653 196348
rect 504587 196283 504653 196284
rect 504587 193220 504653 193221
rect 504587 193156 504588 193220
rect 504652 193156 504653 193220
rect 504587 193155 504653 193156
rect 504590 191453 504650 193155
rect 504587 191452 504653 191453
rect 504587 191388 504588 191452
rect 504652 191388 504653 191452
rect 504587 191387 504653 191388
rect 504038 185950 504466 186010
rect 504038 164250 504098 185950
rect 504403 185876 504469 185877
rect 504403 185812 504404 185876
rect 504468 185812 504469 185876
rect 504403 185811 504469 185812
rect 504219 183836 504285 183837
rect 504219 183772 504220 183836
rect 504284 183772 504285 183836
rect 504219 183771 504285 183772
rect 504222 175813 504282 183771
rect 504219 175812 504285 175813
rect 504219 175748 504220 175812
rect 504284 175748 504285 175812
rect 504219 175747 504285 175748
rect 504219 173228 504285 173229
rect 504219 173164 504220 173228
rect 504284 173164 504285 173228
rect 504219 173163 504285 173164
rect 504222 164933 504282 173163
rect 504219 164932 504285 164933
rect 504219 164868 504220 164932
rect 504284 164868 504285 164932
rect 504219 164867 504285 164868
rect 504038 164190 504282 164250
rect 504035 161396 504101 161397
rect 504035 161332 504036 161396
rect 504100 161332 504101 161396
rect 504035 161331 504101 161332
rect 504038 157997 504098 161331
rect 504035 157996 504101 157997
rect 504035 157932 504036 157996
rect 504100 157932 504101 157996
rect 504035 157931 504101 157932
rect 504222 156090 504282 164190
rect 504038 156030 504282 156090
rect 504038 138685 504098 156030
rect 504219 155820 504285 155821
rect 504219 155756 504220 155820
rect 504284 155756 504285 155820
rect 504219 155755 504285 155756
rect 504035 138684 504101 138685
rect 504035 138620 504036 138684
rect 504100 138620 504101 138684
rect 504035 138619 504101 138620
rect 504035 137324 504101 137325
rect 504035 137260 504036 137324
rect 504100 137260 504101 137324
rect 504035 137259 504101 137260
rect 504038 135149 504098 137259
rect 504035 135148 504101 135149
rect 504035 135084 504036 135148
rect 504100 135084 504101 135148
rect 504035 135083 504101 135084
rect 504035 135012 504101 135013
rect 504035 134948 504036 135012
rect 504100 134948 504101 135012
rect 504035 134947 504101 134948
rect 504038 130661 504098 134947
rect 504035 130660 504101 130661
rect 504035 130596 504036 130660
rect 504100 130596 504101 130660
rect 504035 130595 504101 130596
rect 504035 130524 504101 130525
rect 504035 130460 504036 130524
rect 504100 130460 504101 130524
rect 504035 130459 504101 130460
rect 504038 126037 504098 130459
rect 504035 126036 504101 126037
rect 504035 125972 504036 126036
rect 504100 125972 504101 126036
rect 504035 125971 504101 125972
rect 504035 125220 504101 125221
rect 504035 125156 504036 125220
rect 504100 125156 504101 125220
rect 504035 125155 504101 125156
rect 504038 118285 504098 125155
rect 504035 118284 504101 118285
rect 504035 118220 504036 118284
rect 504100 118220 504101 118284
rect 504035 118219 504101 118220
rect 504035 98700 504101 98701
rect 504035 98636 504036 98700
rect 504100 98636 504101 98700
rect 504035 98635 504101 98636
rect 504038 87685 504098 98635
rect 504222 96797 504282 155755
rect 504406 115293 504466 185811
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504587 178532 504653 178533
rect 504587 178468 504588 178532
rect 504652 178468 504653 178532
rect 504587 178467 504653 178468
rect 504590 172413 504650 178467
rect 504587 172412 504653 172413
rect 504587 172348 504588 172412
rect 504652 172348 504653 172412
rect 504587 172347 504653 172348
rect 504587 165476 504653 165477
rect 504587 165412 504588 165476
rect 504652 165412 504653 165476
rect 504587 165411 504653 165412
rect 504590 158133 504650 165411
rect 504587 158132 504653 158133
rect 504587 158068 504588 158132
rect 504652 158068 504653 158132
rect 504587 158067 504653 158068
rect 504587 157452 504653 157453
rect 504587 157388 504588 157452
rect 504652 157388 504653 157452
rect 504587 157387 504653 157388
rect 504590 122093 504650 157387
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504587 122092 504653 122093
rect 504587 122028 504588 122092
rect 504652 122028 504653 122092
rect 504587 122027 504653 122028
rect 504403 115292 504469 115293
rect 504403 115228 504404 115292
rect 504468 115228 504469 115292
rect 504403 115227 504469 115228
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504403 106044 504469 106045
rect 504403 105980 504404 106044
rect 504468 105980 504469 106044
rect 504403 105979 504469 105980
rect 504406 98701 504466 105979
rect 504403 98700 504469 98701
rect 504403 98636 504404 98700
rect 504468 98636 504469 98700
rect 504403 98635 504469 98636
rect 504219 96796 504285 96797
rect 504219 96732 504220 96796
rect 504284 96732 504285 96796
rect 504219 96731 504285 96732
rect 504219 96524 504285 96525
rect 504219 96460 504220 96524
rect 504284 96460 504285 96524
rect 504219 96459 504285 96460
rect 504035 87684 504101 87685
rect 504035 87620 504036 87684
rect 504100 87620 504101 87684
rect 504035 87619 504101 87620
rect 504222 80205 504282 96459
rect 504219 80204 504285 80205
rect 504219 80140 504220 80204
rect 504284 80140 504285 80204
rect 504219 80139 504285 80140
rect 504035 77348 504101 77349
rect 504035 77284 504036 77348
rect 504100 77284 504101 77348
rect 504035 77283 504101 77284
rect 504219 77348 504285 77349
rect 504219 77284 504220 77348
rect 504284 77284 504285 77348
rect 504219 77283 504285 77284
rect 504038 57629 504098 77283
rect 504035 57628 504101 57629
rect 504035 57564 504036 57628
rect 504100 57564 504101 57628
rect 504035 57563 504101 57564
rect 504222 49061 504282 77283
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504587 57628 504653 57629
rect 504587 57564 504588 57628
rect 504652 57564 504653 57628
rect 504587 57563 504653 57564
rect 504590 49061 504650 57563
rect 504219 49060 504285 49061
rect 504219 48996 504220 49060
rect 504284 48996 504285 49060
rect 504219 48995 504285 48996
rect 504587 49060 504653 49061
rect 504587 48996 504588 49060
rect 504652 48996 504653 49060
rect 504587 48995 504653 48996
rect 504219 38724 504285 38725
rect 504219 38660 504220 38724
rect 504284 38660 504285 38724
rect 504219 38659 504285 38660
rect 504403 38724 504469 38725
rect 504403 38660 504404 38724
rect 504468 38660 504469 38724
rect 504403 38659 504469 38660
rect 503851 17372 503917 17373
rect 503851 17308 503852 17372
rect 503916 17308 503917 17372
rect 503851 17307 503917 17308
rect 504222 16149 504282 38659
rect 504219 16148 504285 16149
rect 504219 16084 504220 16148
rect 504284 16084 504285 16148
rect 504219 16083 504285 16084
rect 504406 10301 504466 38659
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504403 10300 504469 10301
rect 504403 10236 504404 10300
rect 504468 10236 504469 10300
rect 504403 10235 504469 10236
rect 503299 4860 503365 4861
rect 503299 4796 503300 4860
rect 503364 4796 503365 4860
rect 503299 4795 503365 4796
rect 502011 3908 502077 3909
rect 502011 3844 502012 3908
rect 502076 3844 502077 3908
rect 502011 3843 502077 3844
rect 501643 3092 501709 3093
rect 501643 3028 501644 3092
rect 501708 3028 501709 3092
rect 501643 3027 501709 3028
rect 504804 2454 505404 37898
rect 505510 18597 505570 570011
rect 505694 121277 505754 696899
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 506243 584764 506309 584765
rect 506243 584700 506244 584764
rect 506308 584700 506309 584764
rect 506243 584699 506309 584700
rect 506059 582588 506125 582589
rect 506059 582524 506060 582588
rect 506124 582524 506125 582588
rect 506059 582523 506125 582524
rect 505875 582452 505941 582453
rect 505875 582388 505876 582452
rect 505940 582388 505941 582452
rect 505875 582387 505941 582388
rect 505691 121276 505757 121277
rect 505691 121212 505692 121276
rect 505756 121212 505757 121276
rect 505691 121211 505757 121212
rect 505691 116788 505757 116789
rect 505691 116724 505692 116788
rect 505756 116724 505757 116788
rect 505691 116723 505757 116724
rect 505694 101421 505754 116723
rect 505691 101420 505757 101421
rect 505691 101356 505692 101420
rect 505756 101356 505757 101420
rect 505691 101355 505757 101356
rect 505878 29069 505938 582387
rect 506062 87005 506122 582523
rect 506246 139365 506306 584699
rect 508404 582054 509004 617498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 509371 583812 509437 583813
rect 509371 583748 509372 583812
rect 509436 583748 509437 583812
rect 509371 583747 509437 583748
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 506427 581500 506493 581501
rect 506427 581436 506428 581500
rect 506492 581436 506493 581500
rect 506427 581435 506493 581436
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 506243 139364 506309 139365
rect 506243 139300 506244 139364
rect 506308 139300 506309 139364
rect 506243 139299 506309 139300
rect 506243 132020 506309 132021
rect 506243 131956 506244 132020
rect 506308 131956 506309 132020
rect 506243 131955 506309 131956
rect 506246 116789 506306 131955
rect 506243 116788 506309 116789
rect 506243 116724 506244 116788
rect 506308 116724 506309 116788
rect 506243 116723 506309 116724
rect 506059 87004 506125 87005
rect 506059 86940 506060 87004
rect 506124 86940 506125 87004
rect 506059 86939 506125 86940
rect 505875 29068 505941 29069
rect 505875 29004 505876 29068
rect 505940 29004 505941 29068
rect 505875 29003 505941 29004
rect 505507 18596 505573 18597
rect 505507 18532 505508 18596
rect 505572 18532 505573 18596
rect 505507 18531 505573 18532
rect 506430 2957 506490 581435
rect 508083 577692 508149 577693
rect 508083 577628 508084 577692
rect 508148 577628 508149 577692
rect 508083 577627 508149 577628
rect 506979 575516 507045 575517
rect 506979 575452 506980 575516
rect 507044 575452 507045 575516
rect 506979 575451 507045 575452
rect 506982 553890 507042 575451
rect 506982 553830 507226 553890
rect 507166 552530 507226 553830
rect 506798 552470 507226 552530
rect 506798 543965 506858 552470
rect 507899 545868 507965 545869
rect 507899 545804 507900 545868
rect 507964 545804 507965 545868
rect 507899 545803 507965 545804
rect 507163 545460 507229 545461
rect 507163 545396 507164 545460
rect 507228 545396 507229 545460
rect 507163 545395 507229 545396
rect 506795 543964 506861 543965
rect 506795 543900 506796 543964
rect 506860 543900 506861 543964
rect 506795 543899 506861 543900
rect 506795 543692 506861 543693
rect 506795 543628 506796 543692
rect 506860 543628 506861 543692
rect 506795 543627 506861 543628
rect 506611 538796 506677 538797
rect 506611 538732 506612 538796
rect 506676 538732 506677 538796
rect 506611 538731 506677 538732
rect 506614 122501 506674 538731
rect 506798 531450 506858 543627
rect 506798 531390 507042 531450
rect 506982 502210 507042 531390
rect 506798 502150 507042 502210
rect 506798 492693 506858 502150
rect 506795 492692 506861 492693
rect 506795 492628 506796 492692
rect 506860 492628 506861 492692
rect 506795 492627 506861 492628
rect 506979 492692 507045 492693
rect 506979 492628 506980 492692
rect 507044 492628 507045 492692
rect 506979 492627 507045 492628
rect 506795 464812 506861 464813
rect 506795 464748 506796 464812
rect 506860 464748 506861 464812
rect 506795 464747 506861 464748
rect 506798 425509 506858 464747
rect 506982 434621 507042 492627
rect 507166 444549 507226 545395
rect 507163 444548 507229 444549
rect 507163 444484 507164 444548
rect 507228 444484 507229 444548
rect 507163 444483 507229 444484
rect 507163 444412 507229 444413
rect 507163 444348 507164 444412
rect 507228 444348 507229 444412
rect 507163 444347 507229 444348
rect 506979 434620 507045 434621
rect 506979 434556 506980 434620
rect 507044 434556 507045 434620
rect 506979 434555 507045 434556
rect 506795 425508 506861 425509
rect 506795 425444 506796 425508
rect 506860 425444 506861 425508
rect 506795 425443 506861 425444
rect 507166 425237 507226 444347
rect 506979 425236 507045 425237
rect 506979 425172 506980 425236
rect 507044 425172 507045 425236
rect 506979 425171 507045 425172
rect 507163 425236 507229 425237
rect 507163 425172 507164 425236
rect 507228 425172 507229 425236
rect 507163 425171 507229 425172
rect 506795 425100 506861 425101
rect 506795 425036 506796 425100
rect 506860 425036 506861 425100
rect 506795 425035 506861 425036
rect 506798 328405 506858 425035
rect 506982 405653 507042 425171
rect 507163 425100 507229 425101
rect 507163 425036 507164 425100
rect 507228 425036 507229 425100
rect 507163 425035 507229 425036
rect 506979 405652 507045 405653
rect 506979 405588 506980 405652
rect 507044 405588 507045 405652
rect 506979 405587 507045 405588
rect 506979 396132 507045 396133
rect 506979 396068 506980 396132
rect 507044 396068 507045 396132
rect 506979 396067 507045 396068
rect 506982 394637 507042 396067
rect 506979 394636 507045 394637
rect 506979 394572 506980 394636
rect 507044 394572 507045 394636
rect 506979 394571 507045 394572
rect 506979 387156 507045 387157
rect 506979 387092 506980 387156
rect 507044 387092 507045 387156
rect 506979 387091 507045 387092
rect 506982 345133 507042 387091
rect 506979 345132 507045 345133
rect 506979 345068 506980 345132
rect 507044 345068 507045 345132
rect 506979 345067 507045 345068
rect 506795 328404 506861 328405
rect 506795 328340 506796 328404
rect 506860 328340 506861 328404
rect 506795 328339 506861 328340
rect 506795 323644 506861 323645
rect 506795 323580 506796 323644
rect 506860 323580 506861 323644
rect 506795 323579 506861 323580
rect 506611 122500 506677 122501
rect 506611 122436 506612 122500
rect 506676 122436 506677 122500
rect 506611 122435 506677 122436
rect 506798 121957 506858 323579
rect 506979 297396 507045 297397
rect 506979 297332 506980 297396
rect 507044 297332 507045 297396
rect 506979 297331 507045 297332
rect 506982 290461 507042 297331
rect 506979 290460 507045 290461
rect 506979 290396 506980 290460
rect 507044 290396 507045 290460
rect 506979 290395 507045 290396
rect 506979 270604 507045 270605
rect 506979 270540 506980 270604
rect 507044 270540 507045 270604
rect 506979 270539 507045 270540
rect 506982 261493 507042 270539
rect 506979 261492 507045 261493
rect 506979 261428 506980 261492
rect 507044 261428 507045 261492
rect 506979 261427 507045 261428
rect 506979 235380 507045 235381
rect 506979 235316 506980 235380
rect 507044 235316 507045 235380
rect 506979 235315 507045 235316
rect 506982 193901 507042 235315
rect 506979 193900 507045 193901
rect 506979 193836 506980 193900
rect 507044 193836 507045 193900
rect 506979 193835 507045 193836
rect 506979 173228 507045 173229
rect 506979 173164 506980 173228
rect 507044 173164 507045 173228
rect 506979 173163 507045 173164
rect 506982 164933 507042 173163
rect 506979 164932 507045 164933
rect 506979 164868 506980 164932
rect 507044 164868 507045 164932
rect 506979 164867 507045 164868
rect 506979 155276 507045 155277
rect 506979 155212 506980 155276
rect 507044 155212 507045 155276
rect 506979 155211 507045 155212
rect 506982 145621 507042 155211
rect 506979 145620 507045 145621
rect 506979 145556 506980 145620
rect 507044 145556 507045 145620
rect 506979 145555 507045 145556
rect 506979 139364 507045 139365
rect 506979 139300 506980 139364
rect 507044 139300 507045 139364
rect 506979 139299 507045 139300
rect 506795 121956 506861 121957
rect 506795 121892 506796 121956
rect 506860 121892 506861 121956
rect 506795 121891 506861 121892
rect 506982 119458 507042 139299
rect 507166 120461 507226 425035
rect 507715 422652 507781 422653
rect 507715 422588 507716 422652
rect 507780 422588 507781 422652
rect 507715 422587 507781 422588
rect 507531 382532 507597 382533
rect 507531 382468 507532 382532
rect 507596 382468 507597 382532
rect 507531 382467 507597 382468
rect 507347 345132 507413 345133
rect 507347 345068 507348 345132
rect 507412 345068 507413 345132
rect 507347 345067 507413 345068
rect 507350 316029 507410 345067
rect 507534 319565 507594 382467
rect 507531 319564 507597 319565
rect 507531 319500 507532 319564
rect 507596 319500 507597 319564
rect 507531 319499 507597 319500
rect 507531 318884 507597 318885
rect 507531 318820 507532 318884
rect 507596 318820 507597 318884
rect 507531 318819 507597 318820
rect 507347 316028 507413 316029
rect 507347 315964 507348 316028
rect 507412 315964 507413 316028
rect 507347 315963 507413 315964
rect 507347 290460 507413 290461
rect 507347 290396 507348 290460
rect 507412 290396 507413 290460
rect 507347 290395 507413 290396
rect 507350 280805 507410 290395
rect 507347 280804 507413 280805
rect 507347 280740 507348 280804
rect 507412 280740 507413 280804
rect 507347 280739 507413 280740
rect 507534 263669 507594 318819
rect 507531 263668 507597 263669
rect 507531 263604 507532 263668
rect 507596 263604 507597 263668
rect 507531 263603 507597 263604
rect 507347 261492 507413 261493
rect 507347 261428 507348 261492
rect 507412 261428 507413 261492
rect 507347 261427 507413 261428
rect 507350 242181 507410 261427
rect 507347 242180 507413 242181
rect 507347 242116 507348 242180
rect 507412 242116 507413 242180
rect 507347 242115 507413 242116
rect 507531 241772 507597 241773
rect 507531 241708 507532 241772
rect 507596 241708 507597 241772
rect 507531 241707 507597 241708
rect 507347 193900 507413 193901
rect 507347 193836 507348 193900
rect 507412 193836 507413 193900
rect 507347 193835 507413 193836
rect 507350 173229 507410 193835
rect 507534 181117 507594 241707
rect 507531 181116 507597 181117
rect 507531 181052 507532 181116
rect 507596 181052 507597 181116
rect 507531 181051 507597 181052
rect 507347 173228 507413 173229
rect 507347 173164 507348 173228
rect 507412 173164 507413 173228
rect 507347 173163 507413 173164
rect 507347 164932 507413 164933
rect 507347 164868 507348 164932
rect 507412 164868 507413 164932
rect 507347 164867 507413 164868
rect 507350 155277 507410 164867
rect 507347 155276 507413 155277
rect 507347 155212 507348 155276
rect 507412 155212 507413 155276
rect 507347 155211 507413 155212
rect 507347 148612 507413 148613
rect 507347 148548 507348 148612
rect 507412 148548 507413 148612
rect 507347 148547 507413 148548
rect 507350 145893 507410 148547
rect 507531 147388 507597 147389
rect 507531 147324 507532 147388
rect 507596 147324 507597 147388
rect 507531 147323 507597 147324
rect 507347 145892 507413 145893
rect 507347 145828 507348 145892
rect 507412 145828 507413 145892
rect 507347 145827 507413 145828
rect 507347 145620 507413 145621
rect 507347 145556 507348 145620
rect 507412 145556 507413 145620
rect 507347 145555 507413 145556
rect 507350 133925 507410 145555
rect 507347 133924 507413 133925
rect 507347 133860 507348 133924
rect 507412 133860 507413 133924
rect 507347 133859 507413 133860
rect 507163 120460 507229 120461
rect 507163 120396 507164 120460
rect 507228 120396 507229 120460
rect 507163 120395 507229 120396
rect 507534 6629 507594 147323
rect 507718 122637 507778 422587
rect 507715 122636 507781 122637
rect 507715 122572 507716 122636
rect 507780 122572 507781 122636
rect 507715 122571 507781 122572
rect 507902 21997 507962 545803
rect 508086 122365 508146 577627
rect 508404 546054 509004 581498
rect 509187 581228 509253 581229
rect 509187 581164 509188 581228
rect 509252 581164 509253 581228
rect 509187 581163 509253 581164
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508267 486028 508333 486029
rect 508267 485964 508268 486028
rect 508332 485964 508333 486028
rect 508267 485963 508333 485964
rect 508083 122364 508149 122365
rect 508083 122300 508084 122364
rect 508148 122300 508149 122364
rect 508083 122299 508149 122300
rect 508270 80069 508330 485963
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508267 80068 508333 80069
rect 508267 80004 508268 80068
rect 508332 80004 508333 80068
rect 508267 80003 508333 80004
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 507899 21996 507965 21997
rect 507899 21932 507900 21996
rect 507964 21932 507965 21996
rect 507899 21931 507965 21932
rect 507531 6628 507597 6629
rect 507531 6564 507532 6628
rect 507596 6564 507597 6628
rect 507531 6563 507597 6564
rect 508404 6054 509004 41498
rect 509190 6085 509250 581163
rect 509374 119237 509434 583747
rect 510659 582316 510725 582317
rect 510659 582252 510660 582316
rect 510724 582252 510725 582316
rect 510659 582251 510725 582252
rect 510107 560012 510173 560013
rect 510107 559948 510108 560012
rect 510172 559948 510173 560012
rect 510107 559947 510173 559948
rect 509739 467940 509805 467941
rect 509739 467876 509740 467940
rect 509804 467876 509805 467940
rect 509739 467875 509805 467876
rect 509742 119645 509802 467875
rect 510110 122858 510170 559947
rect 509739 119644 509805 119645
rect 509739 119580 509740 119644
rect 509804 119580 509805 119644
rect 509739 119579 509805 119580
rect 509371 119236 509437 119237
rect 509371 119172 509372 119236
rect 509436 119172 509437 119236
rect 509371 119171 509437 119172
rect 510662 6901 510722 582251
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 510659 6900 510725 6901
rect 510659 6836 510660 6900
rect 510724 6836 510725 6900
rect 510659 6835 510725 6836
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 509187 6084 509253 6085
rect 509187 6020 509188 6084
rect 509252 6020 509253 6084
rect 509187 6019 509253 6020
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 507715 3772 507781 3773
rect 507715 3708 507716 3772
rect 507780 3708 507781 3772
rect 507715 3707 507781 3708
rect 507718 3178 507778 3707
rect 506427 2956 506493 2957
rect 506427 2892 506428 2956
rect 506492 2892 506493 2956
rect 506427 2891 506493 2892
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 -4026 512604 9098
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 520046 3093 520106 3622
rect 520043 3092 520109 3093
rect 520043 3028 520044 3092
rect 520108 3028 520109 3092
rect 520043 3027 520109 3028
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 531083 3772 531149 3773
rect 531083 3708 531084 3772
rect 531148 3708 531149 3772
rect 531083 3707 531149 3708
rect 531086 3178 531146 3707
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 550587 581364 550653 581365
rect 550587 581300 550588 581364
rect 550652 581300 550653 581364
rect 550587 581299 550653 581300
rect 550590 581093 550650 581299
rect 550587 581092 550653 581093
rect 550587 581028 550588 581092
rect 550652 581028 550653 581092
rect 550587 581027 550653 581028
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 3838 453102 4074 453338
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 75966 216462 76202 216698
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 78542 403462 78778 403698
rect 78542 395982 78778 396218
rect 78174 382382 78410 382618
rect 78174 375582 78410 375818
rect 78174 330702 78410 330938
rect 78174 302822 78410 303058
rect 78174 298742 78410 298978
rect 78174 295492 78410 295578
rect 78174 295428 78260 295492
rect 78260 295428 78324 295492
rect 78324 295428 78410 295492
rect 78174 295342 78410 295428
rect 77806 294662 78042 294898
rect 77806 292622 78042 292858
rect 77438 283782 77674 284018
rect 78174 277662 78410 277898
rect 78174 274262 78410 274498
rect 77438 272902 77674 273138
rect 78174 270862 78410 271098
rect 78174 269652 78410 269738
rect 78174 269588 78260 269652
rect 78260 269588 78324 269652
rect 78324 269588 78410 269652
rect 78174 269502 78410 269588
rect 77806 266102 78042 266338
rect 77806 264062 78042 264298
rect 77806 259982 78042 260218
rect 77806 258622 78042 258858
rect 77438 247892 77674 247978
rect 77438 247828 77524 247892
rect 77524 247828 77588 247892
rect 77588 247828 77674 247892
rect 77438 247742 77674 247828
rect 78174 252502 78410 252738
rect 78174 245022 78410 245258
rect 77806 242302 78042 242538
rect 78174 240942 78410 241178
rect 77990 237692 78226 237778
rect 77990 237628 78076 237692
rect 78076 237628 78140 237692
rect 78140 237628 78226 237692
rect 77990 237542 78226 237628
rect 78174 233462 78410 233698
rect 77806 230742 78042 230978
rect 77806 222582 78042 222818
rect 77806 219862 78042 220098
rect 77806 215782 78042 216018
rect 77806 212382 78042 212618
rect 77438 208302 77674 208538
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 78174 205582 78410 205818
rect 78174 202862 78410 203098
rect 77990 195382 78226 195618
rect 77438 194022 77674 194258
rect 77806 191302 78042 191538
rect 77438 184652 77674 184738
rect 77438 184588 77524 184652
rect 77524 184588 77588 184652
rect 77588 184588 77674 184652
rect 77438 184502 77674 184588
rect 77806 183822 78042 184058
rect 77806 177022 78042 177258
rect 78174 176342 78410 176578
rect 78174 168862 78410 169098
rect 78174 166822 78410 167058
rect 78174 165612 78410 165698
rect 78174 165548 78260 165612
rect 78260 165548 78324 165612
rect 78324 165548 78410 165612
rect 78174 165462 78410 165548
rect 77806 162742 78042 162978
rect 78174 158662 78410 158898
rect 77806 155262 78042 155498
rect 78174 151862 78410 152098
rect 77806 150502 78042 150738
rect 77438 130782 77674 131018
rect 77438 130102 77674 130338
rect 78174 141662 78410 141898
rect 78174 129422 78410 129658
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 82590 574822 82826 575058
rect 82222 570062 82458 570298
rect 83694 574822 83930 575058
rect 84062 573462 84298 573698
rect 84798 573462 85034 573698
rect 82590 569382 82826 569618
rect 83326 565302 83562 565538
rect 84246 569382 84482 569618
rect 83510 559182 83746 559418
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80750 504782 80986 505018
rect 80750 487102 80986 487338
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80750 420462 80986 420698
rect 80750 418422 80986 418658
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80750 394092 80986 394178
rect 80750 394028 80836 394092
rect 80836 394028 80900 394092
rect 80900 394028 80986 394092
rect 80750 393942 80986 394028
rect 80750 393262 80986 393498
rect 80750 385782 80986 386018
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80750 356542 80986 356778
rect 80750 353822 80986 354058
rect 80750 349742 80986 349978
rect 80750 349062 80986 349298
rect 80750 346342 80986 346578
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80750 328662 80986 328898
rect 80750 328132 80986 328218
rect 80750 328068 80836 328132
rect 80836 328068 80900 328132
rect 80900 328068 80986 328132
rect 80750 327982 80986 328068
rect 80750 313022 80986 313258
rect 80750 299422 80986 299658
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 82038 539612 82274 539698
rect 82038 539548 82124 539612
rect 82124 539548 82188 539612
rect 82188 539548 82274 539612
rect 82038 539462 82274 539548
rect 80198 237012 80434 237098
rect 80198 236948 80284 237012
rect 80284 236948 80348 237012
rect 80348 236948 80434 237012
rect 80198 236862 80434 236948
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 77070 3622 77306 3858
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 83510 543542 83746 543778
rect 84430 543542 84666 543778
rect 84062 539462 84298 539698
rect 83326 537422 83562 537658
rect 84062 537422 84298 537658
rect 83694 536062 83930 536298
rect 84430 536062 84666 536298
rect 82774 529942 83010 530178
rect 83142 519062 83378 519298
rect 82406 515662 82642 515898
rect 84062 515662 84298 515898
rect 83694 504782 83930 505018
rect 82590 504102 82826 504338
rect 83142 504102 83378 504338
rect 82222 500852 82458 500938
rect 82222 500788 82308 500852
rect 82308 500788 82372 500852
rect 82372 500788 82458 500852
rect 82222 500702 82458 500788
rect 82222 498132 82458 498218
rect 82222 498068 82308 498132
rect 82308 498068 82372 498132
rect 82372 498068 82458 498132
rect 82222 497982 82458 498068
rect 82222 496622 82458 496858
rect 83510 501382 83746 501618
rect 83694 500702 83930 500938
rect 83142 487102 83378 487338
rect 83142 481662 83378 481898
rect 83142 472822 83378 473058
rect 84246 497982 84482 498218
rect 84246 492542 84482 492778
rect 84430 486422 84666 486658
rect 84430 479622 84666 479858
rect 84430 478942 84666 479178
rect 83326 468742 83562 468978
rect 83326 467382 83562 467618
rect 83878 420462 84114 420698
rect 84062 418422 84298 418658
rect 83326 403462 83562 403698
rect 82590 396662 82826 396898
rect 83326 396662 83562 396898
rect 82958 393942 83194 394178
rect 82958 392582 83194 392818
rect 83510 392582 83746 392818
rect 82774 377622 83010 377858
rect 84062 382382 84298 382618
rect 83694 377622 83930 377858
rect 82774 367422 83010 367658
rect 84062 376942 84298 377178
rect 84062 376262 84298 376498
rect 84430 375582 84666 375818
rect 83694 367422 83930 367658
rect 82958 359262 83194 359498
rect 82774 357222 83010 357458
rect 83510 356270 83746 356506
rect 82774 353142 83010 353378
rect 83510 353822 83746 354058
rect 83510 353142 83746 353378
rect 83142 349742 83378 349978
rect 82590 340902 82826 341138
rect 82406 332212 82642 332298
rect 82406 332148 82492 332212
rect 82492 332148 82556 332212
rect 82556 332148 82642 332212
rect 82406 332062 82642 332148
rect 83510 340902 83746 341138
rect 83142 331382 83378 331618
rect 84614 349062 84850 349298
rect 84430 345662 84666 345898
rect 84430 342942 84666 343178
rect 83878 332062 84114 332298
rect 83326 328662 83562 328898
rect 82958 321182 83194 321418
rect 83694 327982 83930 328218
rect 84614 339542 84850 339778
rect 84246 327302 84482 327538
rect 84246 322542 84482 322778
rect 83694 321862 83930 322098
rect 83694 321182 83930 321418
rect 83142 313022 83378 313258
rect 83510 299422 83746 299658
rect 83510 298742 83746 298978
rect 83142 295342 83378 295578
rect 84430 321182 84666 321418
rect 84430 302822 84666 303058
rect 84430 302142 84666 302378
rect 84430 296022 84666 296258
rect 83878 294662 84114 294898
rect 82958 292622 83194 292858
rect 84246 283782 84482 284018
rect 84246 281062 84482 281298
rect 84430 280382 84666 280618
rect 84062 279702 84298 279938
rect 82958 276982 83194 277218
rect 84062 277262 84298 277498
rect 83878 272902 84114 273138
rect 84614 273582 84850 273818
rect 84430 270862 84666 271098
rect 83326 269502 83562 269738
rect 83326 266102 83562 266338
rect 83326 264062 83562 264298
rect 82958 259982 83194 260218
rect 84062 258622 84298 258858
rect 82958 255222 83194 255458
rect 83694 255222 83930 255458
rect 83510 252502 83746 252738
rect 83878 247742 84114 247978
rect 83878 245022 84114 245258
rect 83142 242302 83378 242538
rect 82774 237542 83010 237778
rect 83510 241622 83746 241858
rect 83510 238222 83746 238458
rect 82452 235638 82688 235874
rect 83878 236862 84114 237098
rect 82590 234142 82826 234378
rect 82958 233462 83194 233698
rect 82406 232102 82642 232338
rect 82774 231422 83010 231658
rect 82452 229532 82688 229618
rect 82452 229468 82492 229532
rect 82492 229468 82556 229532
rect 82556 229468 82688 229532
rect 82452 229382 82688 229468
rect 82406 228022 82642 228258
rect 82590 223942 82826 224178
rect 83878 227342 84114 227578
rect 84246 226390 84482 226626
rect 82958 219182 83194 219418
rect 83326 219182 83562 219418
rect 82406 209132 82642 209218
rect 82406 209068 82492 209132
rect 82492 209068 82556 209132
rect 82556 209068 82642 209132
rect 84246 219182 84482 219418
rect 84430 218502 84666 218738
rect 84062 217142 84298 217378
rect 83694 216462 83930 216698
rect 83878 215782 84114 216018
rect 83510 215102 83746 215338
rect 83326 213742 83562 213978
rect 82406 208982 82642 209068
rect 84798 216462 85034 216698
rect 84798 215782 85034 216018
rect 84430 214422 84666 214658
rect 82958 206262 83194 206498
rect 83694 206262 83930 206498
rect 84614 211702 84850 211938
rect 84614 210342 84850 210578
rect 84798 209662 85034 209898
rect 84246 204902 84482 205138
rect 82590 196742 82826 196978
rect 83142 196062 83378 196298
rect 82774 195382 83010 195618
rect 86270 569822 86506 570058
rect 86638 565302 86874 565538
rect 87006 557822 87242 558058
rect 86638 529942 86874 530178
rect 86638 520422 86874 520658
rect 86638 519742 86874 519978
rect 86638 519062 86874 519298
rect 86822 502062 87058 502298
rect 86638 496622 86874 496858
rect 86638 492542 86874 492778
rect 86638 483022 86874 483258
rect 86638 481662 86874 481898
rect 86638 472142 86874 472378
rect 86638 349742 86874 349978
rect 86638 349062 86874 349298
rect 86638 328662 86874 328898
rect 86638 327982 86874 328218
rect 86638 327302 86874 327538
rect 86270 320042 86506 320278
rect 86270 318462 86506 318698
rect 87190 325262 87426 325498
rect 87190 324582 87426 324818
rect 87558 323902 87794 324138
rect 87926 322542 88162 322778
rect 87006 315902 87242 316138
rect 86638 302142 86874 302378
rect 86822 300102 87058 300338
rect 86638 296022 86874 296258
rect 87374 298062 87610 298298
rect 86270 288302 86506 288538
rect 86270 279702 86506 279938
rect 86270 278342 86506 278578
rect 87558 286502 87794 286738
rect 86270 232782 86506 233018
rect 86454 232102 86690 232338
rect 87006 241622 87242 241858
rect 87558 238902 87794 239138
rect 86638 231422 86874 231658
rect 87558 238222 87794 238458
rect 87558 236862 87794 237098
rect 87144 234142 87380 234378
rect 87374 232782 87610 233018
rect 86454 230062 86690 230298
rect 88294 231422 88530 231658
rect 86270 229382 86506 229618
rect 86270 227342 86506 227578
rect 86638 223262 86874 223498
rect 86638 222582 86874 222818
rect 87374 219182 87610 219418
rect 86270 214422 86506 214658
rect 87742 215782 87978 216018
rect 87558 214422 87794 214658
rect 88294 214422 88530 214658
rect 87926 213062 88162 213298
rect 86638 210342 86874 210578
rect 85902 208302 86138 208538
rect 85902 206262 86138 206498
rect 85166 205582 85402 205818
rect 84798 202182 85034 202418
rect 85534 204902 85770 205138
rect 85166 201502 85402 201738
rect 86270 205582 86506 205818
rect 86638 205582 86874 205818
rect 87374 206126 87610 206362
rect 86822 204902 87058 205138
rect 85902 202182 86138 202418
rect 85902 201502 86138 201738
rect 84798 198782 85034 199018
rect 82774 194702 83010 194938
rect 84614 196062 84850 196298
rect 85902 198782 86138 199018
rect 82774 194022 83010 194258
rect 84246 194702 84482 194938
rect 83510 194022 83746 194258
rect 83878 191982 84114 192218
rect 82406 190844 82492 190858
rect 82492 190844 82556 190858
rect 82556 190844 82642 190858
rect 82406 190622 82642 190844
rect 83510 191302 83746 191538
rect 84246 191302 84482 191538
rect 82590 187902 82826 188138
rect 82590 179062 82826 179298
rect 83694 187222 83930 187458
rect 83878 186542 84114 186778
rect 84798 190622 85034 190858
rect 84798 187902 85034 188138
rect 84614 186542 84850 186778
rect 83326 183142 83562 183378
rect 84430 183142 84666 183378
rect 83326 179742 83562 179978
rect 84062 179742 84298 179978
rect 83326 178382 83562 178618
rect 84246 179062 84482 179298
rect 83510 177022 83746 177258
rect 83326 172262 83562 172498
rect 83878 170222 84114 170458
rect 84062 169542 84298 169778
rect 84246 166822 84482 167058
rect 83878 165462 84114 165698
rect 83694 162742 83930 162978
rect 84246 160702 84482 160938
rect 83694 158662 83930 158898
rect 83878 157982 84114 158218
rect 83694 155262 83930 155498
rect 83510 151862 83746 152098
rect 83510 150502 83746 150738
rect 84062 144382 84298 144618
rect 83694 141662 83930 141898
rect 83878 140982 84114 141218
rect 83510 140302 83746 140538
rect 84246 140302 84482 140538
rect 84246 132822 84482 133058
rect 83878 130782 84114 131018
rect 83510 130102 83746 130338
rect 84062 129422 84298 129658
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 88248 212382 88484 212618
rect 87742 204902 87978 205138
rect 87190 202182 87426 202418
rect 86638 196742 86874 196978
rect 86270 195382 86506 195618
rect 86638 194022 86874 194258
rect 86638 191982 86874 192218
rect 87742 201502 87978 201738
rect 87742 196062 87978 196298
rect 88110 191982 88346 192218
rect 88294 190622 88530 190858
rect 88110 189942 88346 190178
rect 87926 187222 88162 187458
rect 86638 181102 86874 181338
rect 86638 180422 86874 180658
rect 87006 180422 87242 180658
rect 87190 176342 87426 176578
rect 87926 177022 88162 177258
rect 87190 175662 87426 175898
rect 87236 174302 87472 174538
rect 87006 172942 87242 173178
rect 87236 172262 87472 172498
rect 88984 173622 89220 173858
rect 88662 172262 88898 172498
rect 86638 168862 86874 169098
rect 86270 163422 86506 163658
rect 88294 170222 88530 170458
rect 88662 169542 88898 169778
rect 87420 168182 87656 168418
rect 87420 166142 87656 166378
rect 87144 164782 87380 165018
rect 87558 163422 87794 163658
rect 88616 168862 88852 169098
rect 88478 166142 88714 166378
rect 88478 165462 88714 165698
rect 88616 163422 88852 163658
rect 87190 161382 87426 161618
rect 87374 160022 87610 160258
rect 88616 162062 88852 162298
rect 87006 143702 87242 143938
rect 87006 142342 87242 142578
rect 86638 137582 86874 137818
rect 87006 136902 87242 137138
rect 86638 132822 86874 133058
rect 88294 106302 88530 106538
rect 88294 105622 88530 105858
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90502 215102 90738 215338
rect 90686 213742 90922 213978
rect 90502 181102 90738 181338
rect 90686 178382 90922 178618
rect 90502 170222 90738 170458
rect 90686 169542 90922 169778
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 92894 583662 93130 583898
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 93630 584342 93866 584578
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 93998 580262 94234 580498
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 233102 583812 233338 583898
rect 233102 583748 233188 583812
rect 233188 583748 233252 583812
rect 233252 583748 233338 583812
rect 233102 583662 233338 583748
rect 233838 583662 234074 583898
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 99886 580484 99972 580498
rect 99972 580484 100036 580498
rect 100036 580484 100122 580498
rect 99886 580262 100122 580484
rect 105958 580262 106194 580498
rect 113686 580484 113772 580498
rect 113772 580484 113836 580498
rect 113836 580484 113922 580498
rect 113686 580262 113922 580484
rect 114422 580484 114508 580498
rect 114508 580484 114572 580498
rect 114572 580484 114658 580498
rect 114422 580262 114658 580484
rect 123622 580484 123708 580498
rect 123708 580484 123772 580498
rect 123772 580484 123858 580498
rect 123622 580262 123858 580484
rect 124174 580484 124260 580498
rect 124260 580484 124324 580498
rect 124324 580484 124410 580498
rect 124174 580262 124410 580484
rect 137054 580484 137140 580498
rect 137140 580484 137204 580498
rect 137204 580484 137290 580498
rect 137054 580262 137290 580484
rect 142022 580484 142108 580498
rect 142108 580484 142172 580498
rect 142172 580484 142258 580498
rect 142022 580262 142258 580484
rect 151406 580484 151492 580498
rect 151492 580484 151556 580498
rect 151556 580484 151642 580498
rect 151406 580262 151642 580484
rect 151774 580484 151860 580498
rect 151860 580484 151924 580498
rect 151924 580484 152010 580498
rect 151774 580262 152010 580484
rect 161158 580484 161244 580498
rect 161244 580484 161308 580498
rect 161308 580484 161394 580498
rect 161158 580262 161394 580484
rect 166126 580484 166212 580498
rect 166212 580484 166276 580498
rect 166276 580484 166362 580498
rect 166126 580262 166362 580484
rect 167598 580484 167684 580498
rect 167684 580484 167748 580498
rect 167748 580484 167834 580498
rect 167598 580262 167834 580484
rect 197222 580484 197308 580498
rect 197308 580484 197372 580498
rect 197372 580484 197458 580498
rect 197222 580262 197458 580484
rect 206790 580484 206876 580498
rect 206876 580484 206940 580498
rect 206940 580484 207026 580498
rect 206790 580262 207026 580484
rect 215070 580262 215306 580498
rect 215806 580262 216042 580498
rect 216542 580484 216628 580498
rect 216628 580484 216692 580498
rect 216692 580484 216778 580498
rect 216542 580262 216778 580484
rect 226110 580484 226196 580498
rect 226196 580484 226260 580498
rect 226260 580484 226346 580498
rect 226110 580262 226346 580484
rect 226846 580262 227082 580498
rect 227582 580262 227818 580498
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 298054 584342 298290 584578
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 245614 580412 245850 580498
rect 245614 580348 245700 580412
rect 245700 580348 245764 580412
rect 245764 580348 245850 580412
rect 245614 580262 245850 580348
rect 254814 580412 255050 580498
rect 254814 580348 254900 580412
rect 254900 580348 254964 580412
rect 254964 580348 255050 580412
rect 254814 580262 255050 580348
rect 260886 580412 261122 580498
rect 260886 580348 260972 580412
rect 260972 580348 261036 580412
rect 261036 580348 261122 580412
rect 260886 580262 261122 580348
rect 270270 580412 270506 580498
rect 270270 580348 270356 580412
rect 270356 580348 270420 580412
rect 270420 580348 270506 580412
rect 270270 580262 270506 580348
rect 272478 580412 272714 580498
rect 272478 580348 272564 580412
rect 272564 580348 272628 580412
rect 272628 580348 272714 580412
rect 272478 580262 272714 580348
rect 273766 580412 274002 580498
rect 273766 580348 273852 580412
rect 273852 580348 273916 580412
rect 273916 580348 274002 580412
rect 273766 580262 274002 580348
rect 282230 580412 282466 580498
rect 282230 580348 282316 580412
rect 282316 580348 282380 580412
rect 282380 580348 282466 580412
rect 282230 580262 282466 580348
rect 283334 580412 283570 580498
rect 283334 580348 283420 580412
rect 283420 580348 283484 580412
rect 283484 580348 283570 580412
rect 283334 580262 283570 580348
rect 291798 580412 292034 580498
rect 291798 580348 291884 580412
rect 291884 580348 291948 580412
rect 291948 580348 292034 580412
rect 291798 580262 292034 580348
rect 293086 580412 293322 580498
rect 293086 580348 293172 580412
rect 293172 580348 293236 580412
rect 293236 580348 293322 580412
rect 293086 580262 293322 580348
rect 311670 580262 311906 580498
rect 312406 580262 312642 580498
rect 318662 580140 318898 580362
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 328230 580262 328466 580498
rect 330622 580412 330858 580498
rect 330622 580348 330708 580412
rect 330708 580348 330772 580412
rect 330772 580348 330858 580412
rect 330622 580262 330858 580348
rect 331726 580412 331962 580498
rect 331726 580348 331812 580412
rect 331812 580348 331876 580412
rect 331876 580348 331962 580412
rect 331726 580262 331962 580348
rect 337982 580412 338218 580498
rect 337982 580348 338068 580412
rect 338068 580348 338132 580412
rect 338132 580348 338218 580412
rect 337982 580262 338218 580348
rect 341294 580412 341530 580498
rect 341294 580348 341380 580412
rect 341380 580348 341444 580412
rect 341444 580348 341530 580412
rect 341294 580262 341530 580348
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 365030 580262 365266 580498
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 318662 580126 318748 580140
rect 318748 580126 318812 580140
rect 318812 580126 318898 580140
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 499350 583884 499436 583898
rect 499436 583884 499500 583898
rect 499500 583884 499586 583898
rect 101726 578902 101962 579138
rect 101726 576182 101962 576418
rect 101726 573462 101962 573698
rect 101542 540822 101778 541058
rect 101726 535382 101962 535618
rect 101542 521102 101778 521338
rect 101542 519742 101778 519978
rect 101726 487062 101962 487298
rect 101726 458542 101962 458778
rect 101542 456516 101778 456738
rect 101542 456502 101628 456516
rect 101628 456502 101692 456516
rect 101692 456502 101778 456516
rect 101358 451892 101594 451978
rect 101358 451828 101444 451892
rect 101444 451828 101508 451892
rect 101508 451828 101594 451892
rect 101358 451742 101594 451828
rect 101542 446982 101778 447218
rect 101726 394622 101962 394858
rect 101542 392582 101778 392818
rect 101542 378302 101778 378538
rect 101542 376262 101778 376498
rect 101542 324582 101778 324818
rect 101726 322542 101962 322778
rect 101542 305542 101778 305778
rect 101726 303502 101962 303738
rect 499350 583662 499586 583884
rect 498614 568702 498850 568938
rect 499534 568702 499770 568938
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 500638 507502 500874 507738
rect 501374 507502 501610 507738
rect 500822 500022 501058 500258
rect 500086 472822 500322 473058
rect 501006 472822 501242 473058
rect 501926 500022 502162 500258
rect 498614 417062 498850 417298
rect 498614 411622 498850 411858
rect 499718 417062 499954 417298
rect 500454 413662 500690 413898
rect 500270 412302 500506 412538
rect 499902 411622 500138 411858
rect 498430 388502 498666 388738
rect 498614 381022 498850 381258
rect 498062 366742 498298 366978
rect 499350 386462 499586 386698
rect 499902 385102 500138 385338
rect 499350 382382 499586 382618
rect 499350 381022 499586 381258
rect 498430 364702 498666 364938
rect 498062 360622 498298 360858
rect 498614 358582 498850 358818
rect 499902 366742 500138 366978
rect 499166 356542 499402 356778
rect 498982 353822 499218 354058
rect 499902 364702 500138 364938
rect 499534 352462 499770 352698
rect 499534 349742 499770 349978
rect 500638 357222 500874 357458
rect 500270 350422 500506 350658
rect 499166 349062 499402 349298
rect 498614 345662 498850 345898
rect 498246 304862 498482 305098
rect 498982 323902 499218 324138
rect 500270 345662 500506 345898
rect 499902 341582 500138 341818
rect 501190 349062 501426 349298
rect 500270 340222 500506 340458
rect 499350 321862 499586 322098
rect 498798 303502 499034 303738
rect 498062 294662 498298 294898
rect 498430 287182 498666 287418
rect 499166 302142 499402 302378
rect 499166 289222 499402 289458
rect 499718 287862 499954 288098
rect 499166 287182 499402 287418
rect 498062 285142 498298 285378
rect 497510 269502 497746 269738
rect 497510 266102 497746 266338
rect 499166 285822 499402 286058
rect 498430 283782 498666 284018
rect 498798 283782 499034 284018
rect 499166 281742 499402 281978
rect 498430 280382 498666 280618
rect 499166 281062 499402 281298
rect 501742 304862 501978 305098
rect 501742 294662 501978 294898
rect 500086 285142 500322 285378
rect 500638 283782 500874 284018
rect 500270 280382 500506 280618
rect 499166 278342 499402 278578
rect 499166 274262 499402 274498
rect 500638 278342 500874 278578
rect 500638 274806 500874 275042
rect 499166 270182 499402 270418
rect 500086 272902 500322 273138
rect 501006 273582 501242 273818
rect 500454 270862 500690 271098
rect 499902 269502 500138 269738
rect 499534 268822 499770 269058
rect 499166 268142 499402 268378
rect 498798 267462 499034 267698
rect 497878 264062 498114 264298
rect 497878 263382 498114 263618
rect 497510 259982 497746 260218
rect 498062 258622 498298 258858
rect 498062 253182 498298 253418
rect 497694 252502 497930 252738
rect 498062 252502 498298 252738
rect 500454 266102 500690 266338
rect 500086 264062 500322 264298
rect 500822 264062 501058 264298
rect 101542 234142 101778 234378
rect 101542 230062 101778 230298
rect 101358 199462 101594 199698
rect 497878 245022 498114 245258
rect 498614 245974 498850 246210
rect 499350 262702 499586 262938
rect 499350 259302 499586 259538
rect 499350 258622 499586 258858
rect 500454 262702 500690 262938
rect 500086 258622 500322 258858
rect 498246 240942 498482 241178
rect 499534 255494 499770 255730
rect 501006 259302 501242 259538
rect 501006 255902 501242 256138
rect 501006 252502 501242 252738
rect 501006 245022 501242 245258
rect 500270 244342 500506 244578
rect 499166 240942 499402 241178
rect 498798 238222 499034 238458
rect 498798 234822 499034 235058
rect 498062 232782 498298 233018
rect 498430 232782 498666 233018
rect 497878 232102 498114 232338
rect 498430 227342 498666 227578
rect 501374 241772 501610 241858
rect 501374 241708 501460 241772
rect 501460 241708 501524 241772
rect 501524 241708 501610 241772
rect 501374 241622 501610 241708
rect 500270 238222 500506 238458
rect 501006 238222 501242 238458
rect 501006 236862 501242 237098
rect 500454 234142 500690 234378
rect 500086 232782 500322 233018
rect 500822 232782 501058 233018
rect 499902 226662 500138 226898
rect 497878 219182 498114 219418
rect 497510 217142 497746 217378
rect 101542 196062 101778 196298
rect 498982 222582 499218 222818
rect 499902 223942 500138 224178
rect 499902 223262 500138 223498
rect 499534 220542 499770 220778
rect 499350 219862 499586 220098
rect 499534 219182 499770 219418
rect 499534 216462 499770 216698
rect 498798 212382 499034 212618
rect 498798 209662 499034 209898
rect 499166 209662 499402 209898
rect 498798 208982 499034 209218
rect 500822 223262 501058 223498
rect 501190 219862 501426 220098
rect 500270 215102 500506 215338
rect 500270 214422 500506 214658
rect 500086 213742 500322 213978
rect 499534 208982 499770 209218
rect 498246 205582 498482 205818
rect 499534 205582 499770 205818
rect 499166 202862 499402 203098
rect 501006 215102 501242 215338
rect 501190 203084 501276 203098
rect 501276 203084 501340 203098
rect 501340 203084 501426 203098
rect 498430 197422 498666 197658
rect 497510 194022 497746 194258
rect 101726 179742 101962 179978
rect 101542 177702 101778 177938
rect 99150 122844 99236 122858
rect 99236 122844 99300 122858
rect 99300 122844 99386 122858
rect 99150 122622 99386 122844
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 114790 2956 115026 3178
rect 114790 2942 114876 2956
rect 114876 2942 114940 2956
rect 114940 2942 115026 2956
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 176062 123302 176298 123538
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 127670 2942 127906 3178
rect 128406 2942 128642 3178
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 148094 121942 148330 122178
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 146990 2942 147226 3178
rect 147726 2942 147962 3178
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 163918 119902 164154 120138
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 164286 4452 164522 4538
rect 164286 4388 164372 4452
rect 164372 4388 164436 4452
rect 164436 4388 164522 4452
rect 164286 4302 164522 4388
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 169070 3622 169306 3858
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 174406 119902 174642 120138
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 172382 3622 172618 3858
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 183238 118692 183474 118778
rect 183238 118628 183324 118692
rect 183324 118628 183388 118692
rect 183388 118628 183474 118692
rect 183238 118542 183474 118628
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 186182 118692 186418 118778
rect 186182 118628 186268 118692
rect 186268 118628 186332 118692
rect 186332 118628 186418 118692
rect 186182 118542 186418 118628
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 181950 4452 182186 4538
rect 181950 4388 182036 4452
rect 182036 4388 182100 4452
rect 182100 4388 182186 4452
rect 181950 4302 182186 4388
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 190414 118692 190650 118778
rect 190414 118628 190500 118692
rect 190500 118628 190564 118692
rect 190564 118628 190650 118692
rect 190414 118542 190650 118628
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 193174 120124 193260 120138
rect 193260 120124 193324 120138
rect 193324 120124 193410 120138
rect 193174 119902 193410 120124
rect 196486 119222 196722 119458
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 204950 2942 205186 3178
rect 205686 2942 205922 3178
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 209734 123316 209970 123538
rect 209734 123302 209820 123316
rect 209820 123302 209884 123316
rect 209884 123302 209970 123316
rect 215070 121956 215306 122178
rect 215070 121942 215156 121956
rect 215156 121942 215220 121956
rect 215220 121942 215306 121956
rect 215438 121956 215674 122178
rect 215438 121942 215524 121956
rect 215524 121942 215588 121956
rect 215588 121942 215674 121956
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 219118 123316 219354 123538
rect 219118 123302 219204 123316
rect 219204 123302 219268 123316
rect 219268 123302 219354 123316
rect 234022 123524 234108 123538
rect 234108 123524 234172 123538
rect 234172 123524 234258 123538
rect 234022 123302 234258 123524
rect 235126 123524 235212 123538
rect 235212 123524 235276 123538
rect 235276 123524 235362 123538
rect 235126 123302 235362 123524
rect 240094 123524 240180 123538
rect 240180 123524 240244 123538
rect 240244 123524 240330 123538
rect 240094 123302 240330 123524
rect 252974 123524 253060 123538
rect 253060 123524 253124 123538
rect 253124 123524 253210 123538
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 243406 121942 243642 122178
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 251134 119902 251370 120138
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 243590 3622 243826 3858
rect 243406 3092 243642 3178
rect 243406 3028 243492 3092
rect 243492 3028 243556 3092
rect 243556 3028 243642 3092
rect 243406 2942 243642 3028
rect 244142 2942 244378 3178
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252974 123302 253210 123524
rect 257942 123452 258178 123538
rect 257942 123388 258028 123452
rect 258028 123388 258092 123452
rect 258092 123388 258178 123452
rect 257942 123302 258178 123388
rect 259966 123452 260202 123538
rect 259966 123388 260052 123452
rect 260052 123388 260116 123452
rect 260116 123388 260202 123452
rect 259966 123302 260202 123388
rect 258494 122622 258730 122858
rect 259230 122622 259466 122858
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 259230 121942 259466 122178
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 265486 118692 265722 118778
rect 265486 118628 265572 118692
rect 265572 118628 265636 118692
rect 265636 118628 265722 118692
rect 265486 118542 265722 118628
rect 269718 118692 269954 118778
rect 269718 118628 269804 118692
rect 269804 118628 269868 118692
rect 269868 118628 269954 118692
rect 269718 118542 269954 118628
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 268798 3622 269034 3858
rect 264382 2956 264618 3178
rect 264382 2942 264468 2956
rect 264468 2942 264532 2956
rect 264532 2942 264618 2956
rect 267510 3092 267746 3178
rect 267510 3028 267596 3092
rect 267596 3028 267660 3092
rect 267660 3028 267746 3092
rect 267510 2942 267746 3028
rect 273582 119222 273818 119458
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 273214 4302 273450 4538
rect 272662 3622 272898 3858
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 281126 121942 281362 122178
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 293086 121942 293322 122178
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 301366 121942 301602 122178
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 301918 3092 302154 3178
rect 301918 3028 302004 3092
rect 302004 3028 302068 3092
rect 302068 3028 302154 3092
rect 301918 2942 302154 3028
rect 306150 3092 306386 3178
rect 306150 3028 306236 3092
rect 306236 3028 306300 3092
rect 306300 3028 306386 3092
rect 306150 2942 306386 3028
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 315902 118692 316138 118778
rect 315902 118628 315988 118692
rect 315988 118628 316052 118692
rect 316052 118628 316138 118692
rect 315902 118542 316138 118628
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 315902 3092 316138 3178
rect 315902 3028 315988 3092
rect 315988 3028 316052 3092
rect 316052 3028 316138 3092
rect 315902 2942 316138 3028
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 420046 123302 420282 123538
rect 342214 122622 342450 122858
rect 379198 122844 379284 122858
rect 379284 122844 379348 122858
rect 379348 122844 379434 122858
rect 322526 121942 322762 122178
rect 326758 119902 326994 120138
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 330990 121942 331226 122178
rect 331174 120052 331410 120138
rect 331174 119988 331260 120052
rect 331260 119988 331324 120052
rect 331324 119988 331410 120052
rect 331174 119902 331410 119988
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 325470 3092 325706 3178
rect 325470 3028 325556 3092
rect 325556 3028 325620 3092
rect 325620 3028 325706 3092
rect 325470 2942 325706 3028
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 329150 4452 329386 4538
rect 329150 4388 329236 4452
rect 329236 4388 329300 4452
rect 329300 4388 329386 4452
rect 329150 4302 329386 4388
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 340558 119222 340794 119458
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 335222 2956 335458 3178
rect 335222 2942 335308 2956
rect 335308 2942 335372 2956
rect 335372 2942 335458 2956
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 337798 4452 338034 4538
rect 337798 4388 337884 4452
rect 337884 4388 337948 4452
rect 337948 4388 338034 4452
rect 337798 4302 338034 4388
rect 344790 121942 345026 122178
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 340742 2956 340978 3178
rect 340742 2942 340828 2956
rect 340828 2942 340892 2956
rect 340892 2942 340978 2956
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 379198 122622 379434 122844
rect 417470 122844 417556 122858
rect 417556 122844 417620 122858
rect 417620 122844 417706 122858
rect 417470 122622 417706 122844
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 369814 121942 370050 122178
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 367054 4302 367290 4538
rect 367606 3622 367842 3858
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 376622 120052 376858 120138
rect 376622 119988 376708 120052
rect 376708 119988 376772 120052
rect 376772 119988 376858 120052
rect 376622 119902 376858 119988
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378462 3092 378698 3178
rect 378462 3028 378548 3092
rect 378548 3028 378612 3092
rect 378612 3028 378698 3092
rect 378462 2942 378698 3028
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 379566 3092 379802 3178
rect 379566 3028 379652 3092
rect 379652 3028 379716 3092
rect 379716 3028 379802 3092
rect 379566 2942 379802 3028
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 394654 119222 394890 119458
rect 394470 118692 394706 118778
rect 394470 118628 394556 118692
rect 394556 118628 394620 118692
rect 394620 118628 394706 118692
rect 394470 118542 394706 118628
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 398150 121942 398386 122178
rect 399070 121942 399306 122178
rect 399438 119222 399674 119458
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 395942 4452 396178 4538
rect 395942 4388 396028 4452
rect 396028 4388 396092 4452
rect 396092 4388 396178 4452
rect 395942 4302 396178 4388
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 398150 2942 398386 3178
rect 398886 2942 399122 3178
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 408454 119222 408690 119458
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 405510 4452 405746 4538
rect 405510 4388 405596 4452
rect 405596 4388 405660 4452
rect 405660 4388 405746 4452
rect 405510 4302 405746 4388
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 415630 4452 415866 4538
rect 415630 4388 415716 4452
rect 415716 4388 415780 4452
rect 415780 4388 415866 4452
rect 415630 4302 415866 4388
rect 417470 3092 417706 3178
rect 417470 3028 417556 3092
rect 417556 3028 417620 3092
rect 417620 3028 417706 3092
rect 417470 2942 417706 3028
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 425014 121942 425250 122178
rect 422806 119222 423042 119458
rect 425014 118692 425250 118778
rect 425014 118628 425100 118692
rect 425100 118628 425164 118692
rect 425164 118628 425250 118692
rect 425014 118542 425250 118628
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 419126 3092 419362 3178
rect 419126 3028 419212 3092
rect 419212 3028 419276 3092
rect 419276 3028 419362 3092
rect 419126 2942 419362 3028
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 424830 4452 425066 4538
rect 424830 4388 424916 4452
rect 424916 4388 424980 4452
rect 424980 4388 425066 4452
rect 424830 4302 425066 4388
rect 434398 122844 434484 122858
rect 434484 122844 434548 122858
rect 434548 122844 434634 122858
rect 434398 122622 434634 122844
rect 444150 122622 444386 122858
rect 434582 122164 434668 122178
rect 434668 122164 434732 122178
rect 434732 122164 434818 122178
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 434582 121942 434818 122164
rect 434214 119222 434450 119458
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 434582 4452 434818 4538
rect 434582 4388 434668 4452
rect 434668 4388 434732 4452
rect 434732 4388 434818 4452
rect 434582 4302 434818 4388
rect 436054 3092 436290 3178
rect 436054 3028 436140 3092
rect 436140 3028 436204 3092
rect 436204 3028 436290 3092
rect 436054 2942 436290 3028
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 437342 3092 437578 3178
rect 437342 3028 437428 3092
rect 437428 3028 437492 3092
rect 437492 3028 437578 3092
rect 437342 2942 437578 3028
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 446542 120124 446628 120138
rect 446628 120124 446692 120138
rect 446692 120124 446778 120138
rect 446542 119902 446778 120124
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 443230 4452 443466 4538
rect 443230 4388 443316 4452
rect 443316 4388 443380 4452
rect 443380 4388 443466 4452
rect 443230 4302 443466 4388
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 453534 119222 453770 119458
rect 453902 119222 454138 119458
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 444334 4316 444570 4538
rect 444334 4302 444420 4316
rect 444420 4302 444484 4316
rect 444484 4302 444570 4316
rect 457214 119222 457450 119458
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 451510 2942 451746 3178
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 457398 3622 457634 3858
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 460894 3772 461130 3858
rect 460894 3708 460980 3772
rect 460980 3708 461044 3772
rect 461044 3708 461130 3772
rect 460894 3622 461130 3708
rect 461262 2942 461498 3178
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 462366 4302 462602 4538
rect 466230 123316 466466 123538
rect 466230 123302 466316 123316
rect 466316 123302 466380 123316
rect 466380 123302 466466 123316
rect 473958 123316 474194 123538
rect 473958 123302 474044 123316
rect 474044 123302 474108 123316
rect 474108 123302 474194 123316
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 470462 2942 470698 3178
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 485550 2942 485786 3178
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 496406 123302 496642 123538
rect 497142 123302 497378 123538
rect 495854 122622 496090 122858
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 498430 195382 498666 195618
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 495118 4302 495354 4538
rect 498246 183142 498482 183378
rect 499718 198782 499954 199018
rect 501190 202862 501426 203084
rect 501006 202182 501242 202418
rect 502110 231422 502346 231658
rect 500638 198782 500874 199018
rect 500086 196742 500322 196978
rect 500086 195382 500322 195618
rect 500086 194022 500322 194258
rect 501374 194702 501610 194938
rect 501374 194022 501610 194258
rect 499902 191302 500138 191538
rect 499350 190622 499586 190858
rect 498798 179742 499034 179978
rect 499718 183142 499954 183378
rect 498982 178382 499218 178618
rect 500454 178382 500690 178618
rect 499718 177702 499954 177938
rect 498982 175662 499218 175898
rect 498614 173622 498850 173858
rect 498246 172262 498482 172498
rect 498246 168862 498482 169098
rect 498062 166822 498298 167058
rect 499350 172262 499586 172498
rect 499350 170358 499586 170594
rect 499166 168862 499402 169098
rect 500270 177022 500506 177258
rect 500270 173622 500506 173858
rect 499718 165462 499954 165698
rect 499350 162742 499586 162978
rect 498062 148462 498298 148698
rect 498430 147782 498666 148018
rect 500638 169542 500874 169778
rect 500638 166822 500874 167058
rect 500638 165462 500874 165698
rect 499718 160702 499954 160938
rect 499718 155942 499954 156178
rect 499718 155262 499954 155498
rect 499350 150502 499586 150738
rect 499166 148734 499402 148970
rect 500270 150502 500506 150738
rect 498246 147102 498482 147338
rect 498246 145062 498482 145298
rect 498614 144382 498850 144618
rect 500270 148462 500506 148698
rect 499350 147782 499586 148018
rect 499902 147102 500138 147338
rect 501006 147102 501242 147338
rect 499212 145062 499448 145298
rect 499902 145062 500138 145298
rect 500638 145062 500874 145298
rect 499902 144382 500138 144618
rect 498982 140302 499218 140538
rect 499350 140302 499586 140538
rect 498430 133502 498666 133738
rect 498062 132822 498298 133058
rect 498430 130782 498666 131018
rect 499212 136222 499448 136458
rect 499212 134182 499448 134418
rect 499212 133502 499448 133738
rect 499212 130782 499448 131018
rect 499902 136902 500138 137138
rect 501190 137052 501426 137138
rect 501190 136988 501276 137052
rect 501276 136988 501340 137052
rect 501340 136988 501426 137052
rect 501190 136902 501426 136988
rect 500822 136222 501058 136458
rect 499902 130782 500138 131018
rect 499350 129422 499586 129658
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 498614 2942 498850 3178
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 503582 453782 503818 454018
rect 503214 388502 503450 388738
rect 503214 385102 503450 385338
rect 503214 382532 503450 382618
rect 503214 382468 503300 382532
rect 503300 382468 503364 382532
rect 503364 382468 503450 382532
rect 503214 382382 503450 382468
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504502 270332 504738 270418
rect 504502 270268 504588 270332
rect 504588 270268 504652 270332
rect 504652 270268 504738 270332
rect 504502 270182 504738 270268
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504502 219182 504738 219418
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504502 215102 504738 215338
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 506894 119222 507130 119458
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 510022 122622 510258 122858
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 507630 2942 507866 3178
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 513886 3092 514122 3178
rect 513886 3028 513972 3092
rect 513972 3028 514036 3092
rect 514036 3028 514122 3092
rect 513886 2942 514122 3028
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 519958 3622 520194 3858
rect 521614 3772 521850 3858
rect 521614 3708 521700 3772
rect 521700 3708 521764 3772
rect 521764 3708 521850 3772
rect 521614 3622 521850 3708
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 530998 2942 531234 3178
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 557862 3772 558098 3858
rect 557862 3708 557948 3772
rect 557948 3708 558012 3772
rect 558012 3708 558098 3772
rect 557862 3622 558098 3708
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect 93588 584578 298332 584620
rect 93588 584342 93630 584578
rect 93866 584342 298054 584578
rect 298290 584342 298332 584578
rect 93588 584300 298332 584342
rect 92852 583898 233380 583940
rect 92852 583662 92894 583898
rect 93130 583662 233102 583898
rect 233338 583662 233380 583898
rect 92852 583620 233380 583662
rect 233796 583898 499628 583940
rect 233796 583662 233838 583898
rect 234074 583662 499350 583898
rect 499586 583662 499628 583898
rect 233796 583620 499628 583662
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect 151364 580540 151868 580676
rect 93956 580498 100164 580540
rect 93956 580262 93998 580498
rect 94234 580262 99886 580498
rect 100122 580262 100164 580498
rect 93956 580220 100164 580262
rect 105916 580498 106236 580540
rect 105916 580262 105958 580498
rect 106194 580262 106236 580498
rect 105916 579180 106236 580262
rect 113644 580498 113964 580540
rect 113644 580262 113686 580498
rect 113922 580262 113964 580498
rect 113644 579860 113964 580262
rect 114380 580498 114700 580540
rect 114380 580262 114422 580498
rect 114658 580262 114700 580498
rect 114380 579860 114700 580262
rect 123580 580498 124452 580540
rect 123580 580262 123622 580498
rect 123858 580262 124174 580498
rect 124410 580262 124452 580498
rect 123580 580220 124452 580262
rect 137012 580498 137332 580540
rect 137012 580262 137054 580498
rect 137290 580262 137332 580498
rect 113644 579540 114700 579860
rect 137012 579860 137332 580262
rect 141980 580498 142300 580540
rect 141980 580262 142022 580498
rect 142258 580262 142300 580498
rect 137012 579540 138988 579860
rect 101684 579138 106236 579180
rect 101684 578902 101726 579138
rect 101962 578902 106236 579138
rect 101684 578860 106236 578902
rect 138668 579180 138988 579540
rect 141980 579180 142300 580262
rect 151364 580498 152052 580540
rect 151364 580262 151406 580498
rect 151642 580262 151774 580498
rect 152010 580262 152052 580498
rect 151364 580220 152052 580262
rect 151548 579540 152052 580220
rect 161116 580498 161436 580540
rect 161116 580262 161158 580498
rect 161394 580262 161436 580498
rect 138668 578860 142300 579180
rect 161116 579180 161436 580262
rect 166084 580498 166404 580540
rect 166084 580262 166126 580498
rect 166362 580262 166404 580498
rect 166084 579180 166404 580262
rect 167556 580498 167876 580540
rect 167556 580262 167598 580498
rect 167834 580262 167876 580498
rect 167556 579860 167876 580262
rect 197180 580498 197500 580540
rect 197180 580262 197222 580498
rect 197458 580262 197500 580498
rect 197180 579860 197500 580262
rect 167556 579540 172660 579860
rect 161116 578860 166404 579180
rect 172340 579180 172660 579540
rect 187612 579540 197500 579860
rect 206748 580498 207068 580540
rect 206748 580262 206790 580498
rect 207026 580262 207068 580498
rect 206748 579860 207068 580262
rect 215028 580498 215348 580540
rect 215028 580262 215070 580498
rect 215306 580262 215348 580498
rect 215028 579860 215348 580262
rect 206748 579540 215348 579860
rect 215764 580498 216084 580540
rect 215764 580262 215806 580498
rect 216042 580262 216084 580498
rect 215764 579860 216084 580262
rect 216500 580498 216820 580540
rect 216500 580262 216542 580498
rect 216778 580262 216820 580498
rect 216500 579860 216820 580262
rect 226068 580498 227124 580540
rect 226068 580262 226110 580498
rect 226346 580262 226846 580498
rect 227082 580262 227124 580498
rect 226068 580220 227124 580262
rect 227540 580498 237612 580540
rect 227540 580262 227582 580498
rect 227818 580262 237612 580498
rect 227540 580220 237612 580262
rect 215764 579540 216820 579860
rect 187612 579180 187932 579540
rect 172340 578860 187932 579180
rect 206748 578860 207252 579540
rect 237292 579180 237612 580220
rect 245572 580498 245892 580540
rect 245572 580262 245614 580498
rect 245850 580262 245892 580498
rect 245572 579860 245892 580262
rect 238580 579540 245892 579860
rect 254772 580498 255092 580540
rect 254772 580262 254814 580498
rect 255050 580262 255092 580498
rect 238580 579180 238900 579540
rect 237292 578860 238900 579180
rect 254772 579180 255092 580262
rect 260844 580498 261164 580540
rect 260844 580262 260886 580498
rect 261122 580262 261164 580498
rect 260844 579180 261164 580262
rect 270228 580498 270548 580540
rect 270228 580262 270270 580498
rect 270506 580262 270548 580498
rect 270228 579860 270548 580262
rect 272436 580498 272756 580540
rect 272436 580262 272478 580498
rect 272714 580262 272756 580498
rect 272436 579860 272756 580262
rect 273724 580498 282508 580540
rect 273724 580262 273766 580498
rect 274002 580262 282230 580498
rect 282466 580262 282508 580498
rect 273724 580220 282508 580262
rect 283292 580498 283612 580540
rect 283292 580262 283334 580498
rect 283570 580262 283612 580498
rect 270228 579540 272756 579860
rect 283292 579860 283612 580262
rect 291756 580498 292076 580540
rect 291756 580262 291798 580498
rect 292034 580262 292076 580498
rect 291756 579860 292076 580262
rect 283292 579540 292076 579860
rect 293044 580498 293364 580540
rect 293044 580262 293086 580498
rect 293322 580262 293364 580498
rect 254772 578860 261164 579180
rect 293044 579180 293364 580262
rect 298012 580220 307716 580540
rect 298012 579180 298332 580220
rect 293044 578860 298332 579180
rect 307396 579180 307716 580220
rect 311076 580498 311948 580540
rect 311076 580262 311670 580498
rect 311906 580262 311948 580498
rect 311076 580220 311948 580262
rect 312364 580498 318940 580540
rect 312364 580262 312406 580498
rect 312642 580362 318940 580498
rect 312642 580262 318662 580362
rect 312364 580220 318662 580262
rect 311076 579180 311396 580220
rect 318620 580126 318662 580220
rect 318898 580126 318940 580362
rect 328188 580498 330900 580540
rect 328188 580262 328230 580498
rect 328466 580262 330622 580498
rect 330858 580262 330900 580498
rect 328188 580220 330900 580262
rect 331684 580498 332004 580540
rect 331684 580262 331726 580498
rect 331962 580262 332004 580498
rect 318620 580084 318940 580126
rect 331684 579860 332004 580262
rect 337940 580498 338260 580540
rect 337940 580262 337982 580498
rect 338218 580262 338260 580498
rect 337940 579860 338260 580262
rect 341252 580498 365308 580540
rect 341252 580262 341294 580498
rect 341530 580262 365030 580498
rect 365266 580262 365308 580498
rect 341252 580220 365308 580262
rect 331684 579540 338260 579860
rect 307396 578860 311396 579180
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect 101500 576418 102004 576460
rect 101500 576182 101726 576418
rect 101962 576182 102004 576418
rect 101500 576140 102004 576182
rect 82548 575058 83972 575100
rect 82548 574822 82590 575058
rect 82826 574822 83694 575058
rect 83930 574822 83972 575058
rect 82548 574780 83972 574822
rect 101500 573740 101820 576140
rect 84020 573698 85076 573740
rect 84020 573462 84062 573698
rect 84298 573462 84798 573698
rect 85034 573462 85076 573698
rect 84020 573420 85076 573462
rect 101500 573698 102004 573740
rect 101500 573462 101726 573698
rect 101962 573462 102004 573698
rect 101500 573420 102004 573462
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect 82180 570298 85076 570340
rect 82180 570062 82222 570298
rect 82458 570204 85076 570298
rect 82458 570062 86548 570204
rect 82180 570058 86548 570062
rect 82180 570020 86270 570058
rect 84756 569884 86270 570020
rect 86228 569822 86270 569884
rect 86506 569822 86548 570058
rect 86228 569780 86548 569822
rect 82548 569618 84524 569660
rect 82548 569382 82590 569618
rect 82826 569382 84246 569618
rect 84482 569382 84524 569618
rect 82548 569340 84524 569382
rect 498572 568938 499812 568980
rect 498572 568702 498614 568938
rect 498850 568702 499534 568938
rect 499770 568702 499812 568938
rect 498572 568660 499812 568702
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect 83284 565538 86916 565580
rect 83284 565302 83326 565538
rect 83562 565302 86638 565538
rect 86874 565302 86916 565538
rect 83284 565260 86916 565302
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect 83468 559418 83788 559460
rect 83468 559182 83510 559418
rect 83746 559182 83788 559418
rect 83468 558100 83788 559182
rect 83468 558058 87284 558100
rect 83468 557822 87006 558058
rect 87242 557822 87284 558058
rect 83468 557780 87284 557822
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect 83468 543778 84708 543820
rect 83468 543542 83510 543778
rect 83746 543542 84430 543778
rect 84666 543542 84708 543778
rect 83468 543500 84708 543542
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect 101316 541058 101820 541100
rect 101316 540822 101542 541058
rect 101778 540822 101820 541058
rect 101316 540780 101820 540822
rect 81996 539698 84340 539740
rect 81996 539462 82038 539698
rect 82274 539462 84062 539698
rect 84298 539462 84340 539698
rect 81996 539420 84340 539462
rect 83284 537658 84340 537700
rect 83284 537422 83326 537658
rect 83562 537422 84062 537658
rect 84298 537422 84340 537658
rect 83284 537380 84340 537422
rect 83652 536298 84708 536340
rect 83652 536062 83694 536298
rect 83930 536062 84430 536298
rect 84666 536062 84708 536298
rect 83652 536020 84708 536062
rect 101316 535660 101636 540780
rect 101316 535618 102004 535660
rect 101316 535382 101726 535618
rect 101962 535382 102004 535618
rect 101316 535340 102004 535382
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect 82732 530178 86916 530220
rect 82732 529942 82774 530178
rect 83010 529942 86638 530178
rect 86874 529942 86916 530178
rect 82732 529900 86916 529942
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect 101500 521338 102004 521380
rect 101500 521102 101542 521338
rect 101778 521102 102004 521338
rect 101500 521060 102004 521102
rect 86596 520658 86916 520700
rect 86596 520422 86638 520658
rect 86874 520422 86916 520658
rect 86596 519978 86916 520422
rect 101684 520020 102004 521060
rect 86596 519742 86638 519978
rect 86874 519742 86916 519978
rect 86596 519700 86916 519742
rect 101500 519978 102004 520020
rect 101500 519742 101542 519978
rect 101778 519742 102004 519978
rect 101500 519700 102004 519742
rect 83100 519298 86916 519340
rect 83100 519062 83142 519298
rect 83378 519062 86638 519298
rect 86874 519062 86916 519298
rect 83100 519020 86916 519062
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect 82364 515898 84340 515940
rect 82364 515662 82406 515898
rect 82642 515662 84062 515898
rect 84298 515662 84340 515898
rect 82364 515620 84340 515662
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect 500596 507738 501652 507780
rect 500596 507502 500638 507738
rect 500874 507502 501374 507738
rect 501610 507502 501652 507738
rect 500596 507460 501652 507502
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect 80708 505018 83972 505060
rect 80708 504782 80750 505018
rect 80986 504782 83694 505018
rect 83930 504782 83972 505018
rect 80708 504740 83972 504782
rect 82548 504338 83420 504380
rect 82548 504102 82590 504338
rect 82826 504102 83142 504338
rect 83378 504102 83420 504338
rect 82548 504060 83420 504102
rect 82180 502298 87100 502340
rect 82180 502062 86822 502298
rect 87058 502062 87100 502298
rect 82180 502020 87100 502062
rect 82180 500938 82500 502020
rect 83468 501618 84892 501660
rect 83468 501382 83510 501618
rect 83746 501382 84892 501618
rect 83468 501340 84892 501382
rect 84572 500980 84892 501340
rect 82180 500702 82222 500938
rect 82458 500702 82500 500938
rect 82180 500660 82500 500702
rect 83652 500938 84892 500980
rect 83652 500702 83694 500938
rect 83930 500702 84892 500938
rect 83652 500660 84892 500702
rect 500780 500258 502204 500300
rect 500780 500022 500822 500258
rect 501058 500022 501926 500258
rect 502162 500022 502204 500258
rect 500780 499980 502204 500022
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect 82180 498218 84524 498260
rect 82180 497982 82222 498218
rect 82458 497982 84246 498218
rect 84482 497982 84524 498218
rect 82180 497940 84524 497982
rect 82180 496858 86916 496900
rect 82180 496622 82222 496858
rect 82458 496622 86638 496858
rect 86874 496622 86916 496858
rect 82180 496580 86916 496622
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect 84204 492778 86916 492820
rect 84204 492542 84246 492778
rect 84482 492542 86638 492778
rect 86874 492542 86916 492778
rect 84204 492500 86916 492542
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect 80708 487338 83420 487380
rect 80708 487102 80750 487338
rect 80986 487102 83142 487338
rect 83378 487102 83420 487338
rect 101684 487300 102004 487380
rect 80708 487060 83420 487102
rect 101550 487298 102004 487300
rect 101550 487062 101726 487298
rect 101962 487062 102004 487298
rect 101550 486980 102004 487062
rect 84388 486658 84708 486700
rect 84388 486422 84430 486658
rect 84666 486422 84708 486658
rect 84388 483300 84708 486422
rect 84388 483258 86916 483300
rect 84388 483022 86638 483258
rect 86874 483022 86916 483258
rect 84388 482980 86916 483022
rect 83100 481898 86916 481940
rect 83100 481662 83142 481898
rect 83378 481662 86638 481898
rect 86874 481662 86916 481898
rect 83100 481620 86916 481662
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect 84388 479858 84708 479900
rect 84388 479622 84430 479858
rect 84666 479622 84708 479858
rect 84388 479178 84708 479622
rect 84388 478942 84430 479178
rect 84666 478942 84708 479178
rect 84388 478900 84708 478942
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect 83100 473058 86916 473100
rect 83100 472822 83142 473058
rect 83378 472822 86916 473058
rect 83100 472780 86916 472822
rect 500044 473058 501284 473100
rect 500044 472822 500086 473058
rect 500322 472822 501006 473058
rect 501242 472822 501284 473058
rect 500044 472780 501284 472822
rect 86596 472378 86916 472780
rect 86596 472142 86638 472378
rect 86874 472142 86916 472378
rect 86596 472100 86916 472142
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect 83284 468978 83604 469020
rect 83284 468742 83326 468978
rect 83562 468742 83604 468978
rect 83284 467618 83604 468742
rect 83284 467382 83326 467618
rect 83562 467382 83604 467618
rect 83284 467340 83604 467382
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect 101684 458778 102004 458820
rect 101684 458542 101726 458778
rect 101962 458542 102004 458778
rect 101684 456780 102004 458542
rect 101500 456738 102004 456780
rect 101500 456502 101542 456738
rect 101778 456502 102004 456738
rect 101500 456460 102004 456502
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect 16492 454420 26196 454740
rect 16492 453380 16812 454420
rect 3796 453338 16812 453380
rect 3796 453102 3838 453338
rect 4074 453102 16812 453338
rect 3796 453060 16812 453102
rect 25876 453380 26196 454420
rect 35812 454420 45516 454740
rect 35812 453380 36132 454420
rect 25876 453060 36132 453380
rect 45196 453380 45516 454420
rect 55132 454420 60972 454740
rect 55132 453380 55452 454420
rect 45196 453060 55452 453380
rect 60652 453380 60972 454420
rect 99844 454420 101084 454740
rect 66172 453740 92804 454060
rect 66172 453380 66492 453740
rect 60652 453060 66492 453380
rect 92484 453380 92804 453740
rect 99844 453380 100164 454420
rect 100764 454060 101084 454420
rect 113092 454420 122796 454740
rect 100764 453740 101820 454060
rect 92484 453060 100164 453380
rect 101500 453380 101820 453740
rect 113092 453380 113412 454420
rect 101500 453060 113412 453380
rect 122476 453380 122796 454420
rect 132412 454420 142116 454740
rect 132412 453380 132732 454420
rect 122476 453060 132732 453380
rect 141796 453380 142116 454420
rect 151732 454420 161436 454740
rect 151732 453380 152052 454420
rect 141796 453060 152052 453380
rect 161116 453380 161436 454420
rect 171052 454420 180756 454740
rect 171052 453380 171372 454420
rect 161116 453060 171372 453380
rect 180436 453380 180756 454420
rect 190372 454420 200076 454740
rect 190372 453380 190692 454420
rect 180436 453060 190692 453380
rect 199756 453380 200076 454420
rect 209692 454420 219396 454740
rect 209692 453380 210012 454420
rect 199756 453060 210012 453380
rect 219076 453380 219396 454420
rect 229012 454420 238716 454740
rect 229012 453380 229332 454420
rect 219076 453060 229332 453380
rect 238396 453380 238716 454420
rect 248332 454420 258036 454740
rect 248332 453380 248652 454420
rect 238396 453060 248652 453380
rect 257716 453380 258036 454420
rect 267652 454420 277356 454740
rect 267652 453380 267972 454420
rect 257716 453060 267972 453380
rect 277036 453380 277356 454420
rect 286972 454420 296676 454740
rect 286972 453380 287292 454420
rect 277036 453060 287292 453380
rect 296356 453380 296676 454420
rect 306292 454420 315996 454740
rect 306292 453380 306612 454420
rect 296356 453060 306612 453380
rect 315676 453380 315996 454420
rect 325612 454420 335316 454740
rect 325612 453380 325932 454420
rect 315676 453060 325932 453380
rect 334996 453380 335316 454420
rect 344932 454420 354636 454740
rect 344932 453380 345252 454420
rect 334996 453060 345252 453380
rect 354316 453380 354636 454420
rect 364252 454420 373956 454740
rect 364252 453380 364572 454420
rect 354316 453060 364572 453380
rect 373636 453380 373956 454420
rect 383572 454420 393276 454740
rect 383572 453380 383892 454420
rect 373636 453060 383892 453380
rect 392956 453380 393276 454420
rect 402892 454420 412596 454740
rect 402892 453380 403212 454420
rect 392956 453060 403212 453380
rect 412276 453380 412596 454420
rect 422212 454420 431916 454740
rect 422212 453380 422532 454420
rect 412276 453060 422532 453380
rect 431596 453380 431916 454420
rect 441532 454420 451236 454740
rect 441532 453380 441852 454420
rect 431596 453060 441852 453380
rect 450916 453380 451236 454420
rect 460852 454420 470556 454740
rect 460852 453380 461172 454420
rect 450916 453060 461172 453380
rect 470236 453380 470556 454420
rect 480172 454420 486012 454740
rect 480172 453380 480492 454420
rect 470236 453060 480492 453380
rect 485692 453380 486012 454420
rect 497284 454018 503860 454060
rect 497284 453782 503582 454018
rect 503818 453782 503860 454018
rect 497284 453740 503860 453782
rect 497284 453380 497604 453740
rect 485692 453060 497604 453380
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451978 522986 452134
rect 55222 451898 101358 451978
rect -2916 451876 101358 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 101316 451742 101358 451876
rect 101594 451898 522986 451978
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect 101594 451876 586840 451898
rect 101594 451742 101636 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect 101316 451340 101636 451742
rect 100948 451020 101636 451340
rect 100948 447260 101268 451020
rect 100948 447218 101820 447260
rect 100948 446982 101542 447218
rect 101778 446982 101820 447218
rect 100948 446940 101820 446982
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect 80708 420698 84156 420740
rect 80708 420462 80750 420698
rect 80986 420462 83878 420698
rect 84114 420462 84156 420698
rect 80708 420420 84156 420462
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect 80708 418658 84340 418700
rect 80708 418422 80750 418658
rect 80986 418422 84062 418658
rect 84298 418422 84340 418658
rect 80708 418380 84340 418422
rect 498572 417298 499996 417340
rect 498572 417062 498614 417298
rect 498850 417062 499718 417298
rect 499954 417062 499996 417298
rect 498572 417020 499996 417062
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect 500044 413898 500732 413940
rect 500044 413662 500454 413898
rect 500690 413662 500732 413898
rect 500044 413620 500732 413662
rect 500044 412580 500364 413620
rect 500044 412538 500548 412580
rect 500044 412302 500270 412538
rect 500506 412302 500548 412538
rect 500044 412260 500548 412302
rect 498572 411858 500180 411900
rect 498572 411622 498614 411858
rect 498850 411622 499902 411858
rect 500138 411622 500180 411858
rect 498572 411580 500180 411622
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect 78500 403698 83604 403740
rect 78500 403462 78542 403698
rect 78778 403462 83326 403698
rect 83562 403462 83604 403698
rect 78500 403420 83604 403462
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 82548 396898 83604 396940
rect 82548 396662 82590 396898
rect 82826 396662 83326 396898
rect 83562 396662 83604 396898
rect 82548 396620 83604 396662
rect 78500 396218 85076 396260
rect 78500 395982 78542 396218
rect 78778 395982 85076 396218
rect 78500 395940 85076 395982
rect 80708 394178 83236 394220
rect 80708 393942 80750 394178
rect 80986 393942 82958 394178
rect 83194 393942 83236 394178
rect 80708 393900 83236 393942
rect 84756 393540 85076 395940
rect 80708 393498 85076 393540
rect 80708 393262 80750 393498
rect 80986 393262 85076 393498
rect 80708 393220 85076 393262
rect 101684 394858 102004 394900
rect 101684 394622 101726 394858
rect 101962 394622 102004 394858
rect 101684 392860 102004 394622
rect 82916 392818 83788 392860
rect 82916 392582 82958 392818
rect 83194 392582 83510 392818
rect 83746 392582 83788 392818
rect 82916 392540 83788 392582
rect 101500 392818 102004 392860
rect 101500 392582 101542 392818
rect 101778 392582 102004 392818
rect 101500 392540 102004 392582
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect 498388 388738 503492 388780
rect 498388 388502 498430 388738
rect 498666 388502 503214 388738
rect 503450 388502 503492 388738
rect 498388 388460 503492 388502
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect 122476 386060 122980 386740
rect 141796 386060 142300 386740
rect 161116 386060 161620 386740
rect 180436 386060 180940 386740
rect 80708 386018 99796 386060
rect 80708 385782 80750 386018
rect 80986 385782 99796 386018
rect 80708 385740 99796 385782
rect 99476 385380 99796 385740
rect 103708 385740 107156 386060
rect 103708 385380 104028 385740
rect 99476 385060 104028 385380
rect 106836 385380 107156 385740
rect 122476 385740 128500 386060
rect 122476 385380 122796 385740
rect 106836 385060 122796 385380
rect 128180 385380 128500 385740
rect 141796 385740 147820 386060
rect 141796 385380 142116 385740
rect 128180 385060 142116 385380
rect 147500 385380 147820 385740
rect 161116 385740 167140 386060
rect 161116 385380 161436 385740
rect 147500 385060 161436 385380
rect 166820 385380 167140 385740
rect 180436 385740 186460 386060
rect 180436 385380 180756 385740
rect 166820 385060 180756 385380
rect 186140 385380 186460 385740
rect 199756 385380 200260 386740
rect 215028 386420 219580 386740
rect 215028 386060 215348 386420
rect 205460 385740 215348 386060
rect 205460 385380 205780 385740
rect 186140 385060 205780 385380
rect 219260 385380 219580 386420
rect 228828 386420 238900 386740
rect 228828 385380 229148 386420
rect 219260 385060 229148 385380
rect 238580 385380 238900 386420
rect 248148 386420 258220 386740
rect 248148 385380 248468 386420
rect 238580 385060 248468 385380
rect 257900 385380 258220 386420
rect 267468 386420 277540 386740
rect 267468 385380 267788 386420
rect 257900 385060 267788 385380
rect 277220 385380 277540 386420
rect 286788 386420 296860 386740
rect 286788 385380 287108 386420
rect 277220 385060 287108 385380
rect 296540 385380 296860 386420
rect 306108 386420 316180 386740
rect 306108 385380 306428 386420
rect 296540 385060 306428 385380
rect 315860 385380 316180 386420
rect 325428 386420 335500 386740
rect 325428 385380 325748 386420
rect 315860 385060 325748 385380
rect 335180 385380 335500 386420
rect 344748 386420 354820 386740
rect 344748 385380 345068 386420
rect 335180 385060 345068 385380
rect 354500 385380 354820 386420
rect 364068 386420 374140 386740
rect 364068 385380 364388 386420
rect 354500 385060 364388 385380
rect 373820 385380 374140 386420
rect 383388 386420 393460 386740
rect 383388 385380 383708 386420
rect 373820 385060 383708 385380
rect 393140 385380 393460 386420
rect 402708 386420 412780 386740
rect 402708 385380 403028 386420
rect 393140 385060 403028 385380
rect 412460 385380 412780 386420
rect 422028 386420 432100 386740
rect 422028 385380 422348 386420
rect 412460 385060 422348 385380
rect 431780 385380 432100 386420
rect 441348 386420 451420 386740
rect 441348 385380 441668 386420
rect 431780 385060 441668 385380
rect 451100 385380 451420 386420
rect 460668 386420 470740 386740
rect 460668 385380 460988 386420
rect 451100 385060 460988 385380
rect 470420 385380 470740 386420
rect 485508 386698 499628 386740
rect 485508 386462 499350 386698
rect 499586 386462 499628 386698
rect 485508 386420 499628 386462
rect 485508 386060 485828 386420
rect 475940 385740 485828 386060
rect 475940 385380 476260 385740
rect 470420 385060 476260 385380
rect 499860 385338 503492 385380
rect 499860 385102 499902 385338
rect 500138 385102 503214 385338
rect 503450 385102 503492 385338
rect 499860 385060 503492 385102
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect 78132 382618 84340 382660
rect 78132 382382 78174 382618
rect 78410 382382 84062 382618
rect 84298 382382 84340 382618
rect 78132 382340 84340 382382
rect 499308 382618 503492 382660
rect 499308 382382 499350 382618
rect 499586 382382 503214 382618
rect 503450 382382 503492 382618
rect 499308 382340 503492 382382
rect 498572 381258 499628 381300
rect 498572 381022 498614 381258
rect 498850 381022 499350 381258
rect 499586 381022 499628 381258
rect 498572 380980 499628 381022
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect 101316 378538 101820 378580
rect 101316 378302 101542 378538
rect 101778 378302 101820 378538
rect 101316 378260 101820 378302
rect 82732 377858 83972 377900
rect 82732 377622 82774 377858
rect 83010 377622 83694 377858
rect 83930 377622 83972 377858
rect 82732 377580 83972 377622
rect 84020 377178 85076 377220
rect 84020 376942 84062 377178
rect 84298 376942 85076 377178
rect 84020 376900 85076 376942
rect 83652 376498 84340 376540
rect 83652 376262 84062 376498
rect 84298 376262 84340 376498
rect 83652 376220 84340 376262
rect 83652 375860 83972 376220
rect 84756 375860 85076 376900
rect 101316 376540 101636 378260
rect 101316 376498 101820 376540
rect 101316 376262 101542 376498
rect 101778 376262 101820 376498
rect 101316 376220 101820 376262
rect 78132 375818 83972 375860
rect 78132 375582 78174 375818
rect 78410 375582 83972 375818
rect 78132 375540 83972 375582
rect 84388 375818 85076 375860
rect 84388 375582 84430 375818
rect 84666 375582 85076 375818
rect 84388 375540 85076 375582
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect 82732 367658 83972 367700
rect 82732 367422 82774 367658
rect 83010 367422 83694 367658
rect 83930 367422 83972 367658
rect 82732 367380 83972 367422
rect 498020 366978 500180 367020
rect 498020 366742 498062 366978
rect 498298 366742 499902 366978
rect 500138 366742 500180 366978
rect 498020 366700 500180 366742
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect 498388 364938 500180 364980
rect 498388 364702 498430 364938
rect 498666 364702 499902 364938
rect 500138 364702 500180 364938
rect 498388 364660 500180 364702
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect 498020 360858 501652 360900
rect 498020 360622 498062 360858
rect 498298 360622 501652 360858
rect 498020 360580 501652 360622
rect 82916 359498 83236 359540
rect 82916 359262 82958 359498
rect 83194 359262 83236 359498
rect 82916 357500 83236 359262
rect 82732 357458 83236 357500
rect 82732 357222 82774 357458
rect 83010 357222 83236 357458
rect 82732 357180 83236 357222
rect 498572 358818 498892 358860
rect 498572 358582 498614 358818
rect 498850 358582 498892 358818
rect 498572 357500 498892 358582
rect 498572 357458 500916 357500
rect 498572 357222 500638 357458
rect 500874 357222 500916 357458
rect 498572 357180 500916 357222
rect 501332 356820 501652 360580
rect 80708 356778 83236 356820
rect 80708 356542 80750 356778
rect 80986 356548 83236 356778
rect 499124 356778 501652 356820
rect 80986 356542 83788 356548
rect 80708 356506 83788 356542
rect 80708 356500 83510 356506
rect 82916 356270 83510 356500
rect 83746 356270 83788 356506
rect 499124 356542 499166 356778
rect 499402 356542 501652 356778
rect 499124 356500 501652 356542
rect 82916 356228 83788 356270
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect 80708 354058 83788 354100
rect 80708 353822 80750 354058
rect 80986 353822 83510 354058
rect 83746 353822 83788 354058
rect 80708 353780 83788 353822
rect 498940 354058 499628 354100
rect 498940 353822 498982 354058
rect 499218 353822 499628 354058
rect 498940 353780 499628 353822
rect 82732 353378 83788 353420
rect 82732 353142 82774 353378
rect 83010 353142 83510 353378
rect 83746 353142 83788 353378
rect 82732 353100 83788 353142
rect 499308 352740 499628 353780
rect 499308 352698 499812 352740
rect 499308 352462 499534 352698
rect 499770 352462 499812 352698
rect 499308 352420 499812 352462
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect 500228 350658 500548 350700
rect 500228 350422 500270 350658
rect 500506 350422 500548 350658
rect 80708 349978 83420 350020
rect 80708 349742 80750 349978
rect 80986 349742 83142 349978
rect 83378 349742 83420 349978
rect 80708 349700 83420 349742
rect 86596 349978 86916 350020
rect 86596 349742 86638 349978
rect 86874 349742 86916 349978
rect 80708 349298 84892 349340
rect 80708 349062 80750 349298
rect 80986 349062 84614 349298
rect 84850 349062 84892 349298
rect 80708 349020 84892 349062
rect 86596 349298 86916 349742
rect 86596 349062 86638 349298
rect 86874 349062 86916 349298
rect 86596 349020 86916 349062
rect 499124 349978 499812 350020
rect 499124 349742 499534 349978
rect 499770 349742 499812 349978
rect 499124 349700 499812 349742
rect 499124 349298 499444 349700
rect 499124 349062 499166 349298
rect 499402 349062 499444 349298
rect 499124 349020 499444 349062
rect 500228 349340 500548 350422
rect 500228 349298 501468 349340
rect 500228 349062 501190 349298
rect 501426 349062 501468 349298
rect 500228 349020 501468 349062
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect 80708 346578 84892 346620
rect 80708 346342 80750 346578
rect 80986 346342 84892 346578
rect 80708 346300 84892 346342
rect 84572 345940 84892 346300
rect 84388 345898 84892 345940
rect 84388 345662 84430 345898
rect 84666 345662 84892 345898
rect 84388 345620 84892 345662
rect 498572 345898 500548 345940
rect 498572 345662 498614 345898
rect 498850 345662 500270 345898
rect 500506 345662 500548 345898
rect 498572 345620 500548 345662
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect 84388 343178 84892 343220
rect 84388 342942 84430 343178
rect 84666 342942 84892 343178
rect 84388 342900 84892 342942
rect 82548 341138 83788 341180
rect 82548 340902 82590 341138
rect 82826 340902 83510 341138
rect 83746 340902 83788 341138
rect 82548 340860 83788 340902
rect 84572 339778 84892 342900
rect 499860 341818 500180 341860
rect 499860 341582 499902 341818
rect 500138 341582 500180 341818
rect 499860 340500 500180 341582
rect 499860 340458 500548 340500
rect 499860 340222 500270 340458
rect 500506 340222 500548 340458
rect 499860 340180 500548 340222
rect 84572 339542 84614 339778
rect 84850 339542 84892 339778
rect 84572 339500 84892 339542
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect 82364 332298 84156 332340
rect 82364 332062 82406 332298
rect 82642 332062 83878 332298
rect 84114 332062 84156 332298
rect 82364 332020 84156 332062
rect 83100 331618 83420 331660
rect 83100 331382 83142 331618
rect 83378 331382 83420 331618
rect 83100 330980 83420 331382
rect 78132 330938 83420 330980
rect 78132 330702 78174 330938
rect 78410 330702 83420 330938
rect 78132 330660 83420 330702
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect 80708 328898 83604 328940
rect 80708 328662 80750 328898
rect 80986 328662 83326 328898
rect 83562 328662 83604 328898
rect 80708 328620 83604 328662
rect 86596 328898 87652 328940
rect 86596 328662 86638 328898
rect 86874 328662 87652 328898
rect 86596 328620 87652 328662
rect 80708 328218 83972 328260
rect 80708 327982 80750 328218
rect 80986 327982 83694 328218
rect 83930 327982 83972 328218
rect 80708 327940 83972 327982
rect 84388 328218 86916 328260
rect 84388 327982 86638 328218
rect 86874 327982 86916 328218
rect 84388 327940 86916 327982
rect 84388 327580 84708 327940
rect 87332 327580 87652 328620
rect 84204 327538 84708 327580
rect 84204 327302 84246 327538
rect 84482 327302 84708 327538
rect 84204 327260 84708 327302
rect 86596 327538 87652 327580
rect 86596 327302 86638 327538
rect 86874 327302 87652 327538
rect 86596 327260 87652 327302
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect 87148 325498 87468 325540
rect 87148 325262 87190 325498
rect 87426 325262 87468 325498
rect 87148 324818 87468 325262
rect 87148 324582 87190 324818
rect 87426 324582 87468 324818
rect 87148 324540 87468 324582
rect 101132 324818 101820 324860
rect 101132 324582 101542 324818
rect 101778 324582 101820 324818
rect 101132 324540 101820 324582
rect 87516 324138 87836 324180
rect 87516 323902 87558 324138
rect 87794 323902 87836 324138
rect 87516 322820 87836 323902
rect 84204 322778 86548 322820
rect 84204 322542 84246 322778
rect 84482 322542 86548 322778
rect 84204 322500 86548 322542
rect 87516 322778 88204 322820
rect 87516 322542 87926 322778
rect 88162 322542 88204 322778
rect 87516 322500 88204 322542
rect 83652 322098 84708 322140
rect 83652 321862 83694 322098
rect 83930 321862 84708 322098
rect 83652 321820 84708 321862
rect 82916 321418 83972 321460
rect 82916 321182 82958 321418
rect 83194 321182 83694 321418
rect 83930 321182 83972 321418
rect 82916 321140 83972 321182
rect 84388 321418 84708 321820
rect 84388 321182 84430 321418
rect 84666 321182 84708 321418
rect 84388 321140 84708 321182
rect 86228 320278 86548 322500
rect 101132 322140 101452 324540
rect 498940 324138 499260 324180
rect 498940 323902 498982 324138
rect 499218 323902 499260 324138
rect 101684 322778 102004 322820
rect 101684 322542 101726 322778
rect 101962 322542 102004 322778
rect 101684 322140 102004 322542
rect 101132 321820 102004 322140
rect 498940 322140 499260 323902
rect 498940 322098 499628 322140
rect 498940 321862 499350 322098
rect 499586 321862 499628 322098
rect 498940 321820 499628 321862
rect 86228 320042 86270 320278
rect 86506 320042 86548 320278
rect 86228 320000 86548 320042
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 86270 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 86228 318462 86270 318676
rect 86506 318676 592360 318698
rect 86506 318462 86548 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect 86228 316700 86548 318462
rect 86228 316380 87284 316700
rect 86964 316138 87284 316380
rect 86964 315902 87006 316138
rect 87242 315902 87284 316138
rect 86964 315860 87284 315902
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect 80708 313258 83420 313300
rect 80708 313022 80750 313258
rect 80986 313022 83142 313258
rect 83378 313022 83420 313258
rect 80708 312980 83420 313022
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect 101500 305778 101820 305820
rect 101500 305542 101542 305778
rect 101778 305542 101820 305778
rect 101500 304460 101820 305542
rect 498204 305098 502020 305140
rect 498204 304862 498246 305098
rect 498482 304862 501742 305098
rect 501978 304862 502020 305098
rect 498204 304820 502020 304862
rect 101500 304140 102004 304460
rect 101684 303738 102004 304140
rect 101684 303502 101726 303738
rect 101962 303502 102004 303738
rect 101684 303460 102004 303502
rect 498756 303738 499076 303780
rect 498756 303502 498798 303738
rect 499034 303502 499076 303738
rect 78132 303058 84708 303100
rect 78132 302822 78174 303058
rect 78410 302822 84430 303058
rect 84666 302822 84708 303058
rect 78132 302780 84708 302822
rect 498756 302420 499076 303502
rect 84388 302378 86916 302420
rect 84388 302142 84430 302378
rect 84666 302142 86638 302378
rect 86874 302142 86916 302378
rect 84388 302100 86916 302142
rect 498756 302378 499444 302420
rect 498756 302142 499166 302378
rect 499402 302142 499444 302378
rect 498756 302100 499444 302142
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect 86780 300338 87100 300380
rect 86780 300102 86822 300338
rect 87058 300102 87100 300338
rect 80708 299658 83788 299700
rect 80708 299422 80750 299658
rect 80986 299422 83510 299658
rect 83746 299422 83788 299658
rect 80708 299380 83788 299422
rect 78132 298978 83788 299020
rect 78132 298742 78174 298978
rect 78410 298742 83510 298978
rect 83746 298742 83788 298978
rect 78132 298700 83788 298742
rect 86780 298340 87100 300102
rect 86780 298298 87652 298340
rect 86780 298062 87374 298298
rect 87610 298062 87652 298298
rect 86780 298020 87652 298062
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect 84388 296258 86916 296300
rect 84388 296022 84430 296258
rect 84666 296022 86638 296258
rect 86874 296022 86916 296258
rect 84388 295980 86916 296022
rect 78132 295578 83420 295620
rect 78132 295342 78174 295578
rect 78410 295342 83142 295578
rect 83378 295342 83420 295578
rect 78132 295300 83420 295342
rect 77764 294898 84156 294940
rect 77764 294662 77806 294898
rect 78042 294662 83878 294898
rect 84114 294662 84156 294898
rect 77764 294620 84156 294662
rect 498020 294898 502020 294940
rect 498020 294662 498062 294898
rect 498298 294662 501742 294898
rect 501978 294662 502020 294898
rect 498020 294620 502020 294662
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect 77764 292858 83236 292900
rect 77764 292622 77806 292858
rect 78042 292622 82958 292858
rect 83194 292622 83236 292858
rect 77764 292580 83236 292622
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect 499124 289458 500916 289500
rect 499124 289222 499166 289458
rect 499402 289222 500916 289458
rect 499124 289180 500916 289222
rect 86228 288538 87100 288580
rect 86228 288302 86270 288538
rect 86506 288302 87100 288538
rect 86228 288260 87100 288302
rect 86780 288140 87100 288260
rect 500596 288140 500916 289180
rect 86780 287820 88940 288140
rect 499676 288098 500916 288140
rect 499676 287862 499718 288098
rect 499954 287862 500916 288098
rect 499676 287820 500916 287862
rect 88620 286780 88940 287820
rect 87516 286738 88940 286780
rect 87516 286502 87558 286738
rect 87794 286502 88940 286738
rect 87516 286460 88940 286502
rect 498020 287418 498708 287460
rect 498020 287182 498430 287418
rect 498666 287182 498708 287418
rect 498020 287140 498708 287182
rect 499124 287418 499444 287460
rect 499124 287182 499166 287418
rect 499402 287182 499444 287418
rect 498020 285378 498340 287140
rect 499124 286058 499444 287182
rect 499124 285822 499166 286058
rect 499402 285822 499444 286058
rect 499124 285780 499444 285822
rect 498020 285142 498062 285378
rect 498298 285142 498340 285378
rect 498020 285100 498340 285142
rect 500044 285378 500364 285420
rect 500044 285142 500086 285378
rect 500322 285142 500364 285378
rect 500044 284060 500364 285142
rect 77396 284018 84524 284060
rect 77396 283782 77438 284018
rect 77674 283782 84246 284018
rect 84482 283782 84524 284018
rect 77396 283740 84524 283782
rect 498388 284018 499076 284060
rect 498388 283782 498430 284018
rect 498666 283782 498798 284018
rect 499034 283782 499076 284018
rect 498388 283740 499076 283782
rect 500044 284018 500916 284060
rect 500044 283782 500638 284018
rect 500874 283782 500916 284018
rect 500044 283740 500916 283782
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect 499124 281978 499444 282020
rect 499124 281742 499166 281978
rect 499402 281742 499444 281978
rect 84204 281298 84524 281340
rect 84204 281062 84246 281298
rect 84482 281062 84524 281298
rect 84204 280660 84524 281062
rect 499124 281298 499444 281742
rect 499124 281062 499166 281298
rect 499402 281062 499444 281298
rect 499124 281020 499444 281062
rect 84204 280618 84708 280660
rect 84204 280382 84430 280618
rect 84666 280382 84708 280618
rect 84204 280340 84708 280382
rect 498388 280618 500548 280660
rect 498388 280382 498430 280618
rect 498666 280382 500270 280618
rect 500506 280382 500548 280618
rect 498388 280340 500548 280382
rect 84020 279938 86548 279980
rect 84020 279702 84062 279938
rect 84298 279702 86270 279938
rect 86506 279702 86548 279938
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 84020 279676 86548 279702
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect 86228 278578 86548 278620
rect 86228 278342 86270 278578
rect 86506 278342 86548 278578
rect 86228 277940 86548 278342
rect 499124 278578 500916 278620
rect 499124 278342 499166 278578
rect 499402 278342 500638 278578
rect 500874 278342 500916 278578
rect 499124 278300 500916 278342
rect 78132 277898 83236 277940
rect 78132 277662 78174 277898
rect 78410 277662 83236 277898
rect 78132 277620 83236 277662
rect 82916 277218 83236 277620
rect 84020 277620 86548 277940
rect 84020 277498 84340 277620
rect 84020 277262 84062 277498
rect 84298 277262 84340 277498
rect 84020 277220 84340 277262
rect 82916 276982 82958 277218
rect 83194 276982 83236 277218
rect 82916 276940 83236 276982
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect 500596 275042 500916 275084
rect 500596 274806 500638 275042
rect 500874 274806 500916 275042
rect 500596 274540 500916 274806
rect 78132 274498 84892 274540
rect 78132 274262 78174 274498
rect 78410 274262 84892 274498
rect 78132 274220 84892 274262
rect 499124 274498 500916 274540
rect 499124 274262 499166 274498
rect 499402 274262 500916 274498
rect 499124 274220 500916 274262
rect 84572 273818 84892 274220
rect 84572 273582 84614 273818
rect 84850 273582 84892 273818
rect 84572 273540 84892 273582
rect 500044 273818 501284 273860
rect 500044 273582 501006 273818
rect 501242 273582 501284 273818
rect 500044 273540 501284 273582
rect 77396 273138 84156 273180
rect 77396 272902 77438 273138
rect 77674 272902 83878 273138
rect 84114 272902 84156 273138
rect 77396 272860 84156 272902
rect 500044 273138 500364 273540
rect 500044 272902 500086 273138
rect 500322 272902 500364 273138
rect 500044 272860 500364 272902
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect 78132 271098 84708 271140
rect 78132 270862 78174 271098
rect 78410 270862 84430 271098
rect 84666 270862 84708 271098
rect 78132 270820 84708 270862
rect 496732 271098 500732 271140
rect 496732 270862 500454 271098
rect 500690 270862 500732 271098
rect 496732 270820 500732 270862
rect 78132 269738 83604 269780
rect 78132 269502 78174 269738
rect 78410 269502 83326 269738
rect 83562 269502 83604 269738
rect 78132 269460 83604 269502
rect 496732 266380 497052 270820
rect 499124 270418 504780 270460
rect 499124 270182 499166 270418
rect 499402 270182 504502 270418
rect 504738 270182 504780 270418
rect 499124 270140 504780 270182
rect 497468 269738 500180 269780
rect 497468 269502 497510 269738
rect 497746 269502 499902 269738
rect 500138 269502 500180 269738
rect 497468 269460 500180 269502
rect 498020 269058 499812 269100
rect 498020 268822 499534 269058
rect 499770 268822 499812 269058
rect 498020 268780 499812 268822
rect 498020 267060 498340 268780
rect 498756 268378 499444 268420
rect 498756 268142 499166 268378
rect 499402 268142 499444 268378
rect 498756 268100 499444 268142
rect 498756 267698 499076 268100
rect 498756 267462 498798 267698
rect 499034 267462 499076 267698
rect 498756 267420 499076 267462
rect 498020 266740 498524 267060
rect 498204 266380 498524 266740
rect 77764 266338 83604 266380
rect 77764 266102 77806 266338
rect 78042 266102 83326 266338
rect 83562 266102 83604 266338
rect 77764 266060 83604 266102
rect 496732 266338 497788 266380
rect 496732 266102 497510 266338
rect 497746 266102 497788 266338
rect 496732 266060 497788 266102
rect 498204 266338 500732 266380
rect 498204 266102 500454 266338
rect 500690 266102 500732 266338
rect 498204 266060 500732 266102
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect 77764 264298 83604 264340
rect 77764 264062 77806 264298
rect 78042 264062 83326 264298
rect 83562 264062 83604 264298
rect 77764 264020 83604 264062
rect 497100 264298 498156 264340
rect 497100 264062 497878 264298
rect 498114 264062 498156 264298
rect 497100 264020 498156 264062
rect 500044 264298 500364 264340
rect 500044 264062 500086 264298
rect 500322 264062 500364 264298
rect 497100 262980 497420 264020
rect 500044 263660 500364 264062
rect 497836 263618 500364 263660
rect 497836 263382 497878 263618
rect 498114 263382 500364 263618
rect 497836 263340 500364 263382
rect 500780 264298 501100 264340
rect 500780 264062 500822 264298
rect 501058 264062 501100 264298
rect 500780 262980 501100 264062
rect 497100 262938 499628 262980
rect 497100 262702 499350 262938
rect 499586 262702 499628 262938
rect 497100 262660 499628 262702
rect 500412 262938 501100 262980
rect 500412 262702 500454 262938
rect 500690 262702 501100 262938
rect 500412 262660 501100 262702
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect 77764 260218 83236 260260
rect 77764 259982 77806 260218
rect 78042 259982 82958 260218
rect 83194 259982 83236 260218
rect 77764 259940 83236 259982
rect 497468 260218 497972 260260
rect 497468 259982 497510 260218
rect 497746 259982 497972 260218
rect 497468 259940 497972 259982
rect 497652 258900 497972 259940
rect 499308 259538 501284 259580
rect 499308 259302 499350 259538
rect 499586 259302 501006 259538
rect 501242 259302 501284 259538
rect 499308 259260 501284 259302
rect 77764 258858 84340 258900
rect 77764 258622 77806 258858
rect 78042 258622 84062 258858
rect 84298 258622 84340 258858
rect 77764 258580 84340 258622
rect 497652 258858 498340 258900
rect 497652 258622 498062 258858
rect 498298 258622 498340 258858
rect 497652 258580 498340 258622
rect 499308 258858 500364 258900
rect 499308 258622 499350 258858
rect 499586 258622 500086 258858
rect 500322 258622 500364 258858
rect 499308 258580 500364 258622
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect 499492 256138 501284 256180
rect 499492 255902 501006 256138
rect 501242 255902 501284 256138
rect 499492 255860 501284 255902
rect 499492 255730 499812 255860
rect 82916 255458 83972 255500
rect 82916 255222 82958 255458
rect 83194 255222 83694 255458
rect 83930 255222 83972 255458
rect 499492 255494 499534 255730
rect 499770 255494 499812 255730
rect 499492 255452 499812 255494
rect 82916 255180 83972 255222
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect 498020 253418 501284 253460
rect 498020 253182 498062 253418
rect 498298 253182 501284 253418
rect 498020 253140 501284 253182
rect 78132 252738 83788 252780
rect 78132 252502 78174 252738
rect 78410 252502 83510 252738
rect 83746 252502 83788 252738
rect 78132 252460 83788 252502
rect 497652 252738 498340 252780
rect 497652 252502 497694 252738
rect 497930 252502 498062 252738
rect 498298 252502 498340 252738
rect 497652 252460 498340 252502
rect 500964 252738 501284 253140
rect 500964 252502 501006 252738
rect 501242 252502 501284 252738
rect 500964 252460 501284 252502
rect 77396 247978 84156 248020
rect 77396 247742 77438 247978
rect 77674 247742 83878 247978
rect 84114 247742 84156 247978
rect 77396 247700 84156 247742
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect 498572 246210 498892 246252
rect 498572 245980 498614 246210
rect 497100 245974 498614 245980
rect 498850 245974 498892 246210
rect 497100 245660 498892 245974
rect 78132 245258 84156 245300
rect 78132 245022 78174 245258
rect 78410 245022 83878 245258
rect 84114 245022 84156 245258
rect 78132 244980 84156 245022
rect 497100 244620 497420 245660
rect 497836 245258 501284 245300
rect 497836 245022 497878 245258
rect 498114 245022 501006 245258
rect 501242 245022 501284 245258
rect 497836 244980 501284 245022
rect 497100 244578 500548 244620
rect 497100 244342 500270 244578
rect 500506 244342 500548 244578
rect 497100 244300 500548 244342
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect 77764 242538 83420 242580
rect 77764 242302 77806 242538
rect 78042 242302 83142 242538
rect 83378 242302 83420 242538
rect 77764 242260 83420 242302
rect 99844 242260 108996 242580
rect 83468 241858 87284 241900
rect 83468 241622 83510 241858
rect 83746 241622 87006 241858
rect 87242 241622 87284 241858
rect 83468 241580 87284 241622
rect 99844 241220 100164 242260
rect 78132 241178 100164 241220
rect 78132 240942 78174 241178
rect 78410 240942 100164 241178
rect 78132 240900 100164 240942
rect 108676 241220 108996 242260
rect 195892 242260 205596 242580
rect 195892 241220 196212 242260
rect 108676 240900 196212 241220
rect 205276 241220 205596 242260
rect 215212 242260 224916 242580
rect 215212 241220 215532 242260
rect 205276 240900 215532 241220
rect 224596 241220 224916 242260
rect 234532 242260 244236 242580
rect 234532 241220 234852 242260
rect 224596 240900 234852 241220
rect 243916 241220 244236 242260
rect 253852 242260 263556 242580
rect 253852 241220 254172 242260
rect 243916 240900 254172 241220
rect 263236 241220 263556 242260
rect 273172 242260 282876 242580
rect 273172 241220 273492 242260
rect 263236 240900 273492 241220
rect 282556 241220 282876 242260
rect 292492 242260 302196 242580
rect 292492 241220 292812 242260
rect 282556 240900 292812 241220
rect 301876 241220 302196 242260
rect 311812 242260 321516 242580
rect 311812 241220 312132 242260
rect 301876 240900 312132 241220
rect 321196 241220 321516 242260
rect 331132 242260 340836 242580
rect 331132 241220 331452 242260
rect 321196 240900 331452 241220
rect 340516 241220 340836 242260
rect 350452 242260 360156 242580
rect 350452 241220 350772 242260
rect 340516 240900 350772 241220
rect 359836 241220 360156 242260
rect 369772 242260 379476 242580
rect 369772 241220 370092 242260
rect 359836 240900 370092 241220
rect 379156 241220 379476 242260
rect 389092 242260 398796 242580
rect 389092 241220 389412 242260
rect 379156 240900 389412 241220
rect 398476 241220 398796 242260
rect 408412 242260 418116 242580
rect 408412 241220 408732 242260
rect 398476 240900 408732 241220
rect 417796 241220 418116 242260
rect 427732 242260 437436 242580
rect 427732 241220 428052 242260
rect 417796 240900 428052 241220
rect 437116 241220 437436 242260
rect 447052 242260 456756 242580
rect 447052 241220 447372 242260
rect 437116 240900 447372 241220
rect 456436 241220 456756 242260
rect 466372 242260 470004 242580
rect 466372 241220 466692 242260
rect 456436 240900 466692 241220
rect 469684 241220 470004 242260
rect 497652 241900 499076 242172
rect 493236 241858 501652 241900
rect 493236 241852 501374 241858
rect 493236 241580 497972 241852
rect 498756 241622 501374 241852
rect 501610 241622 501652 241858
rect 498756 241580 501652 241622
rect 493236 241220 493556 241580
rect 469684 240900 493556 241220
rect 498204 241178 499444 241220
rect 498204 240942 498246 241178
rect 498482 240942 499166 241178
rect 499402 240942 499444 241178
rect 498204 240900 499444 240942
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect 86780 239138 87836 239180
rect 86780 238902 87558 239138
rect 87794 238902 87836 239138
rect 86780 238860 87836 238902
rect 86780 238500 87100 238860
rect 77258 238458 83788 238500
rect 77258 238222 83510 238458
rect 83746 238222 83788 238458
rect 77258 238180 83788 238222
rect 84204 238180 87100 238500
rect 87516 238458 87836 238500
rect 87516 238222 87558 238458
rect 87794 238222 87836 238458
rect 77258 237140 77578 238180
rect 77948 237778 83052 237820
rect 77948 237542 77990 237778
rect 78226 237542 82774 237778
rect 83010 237542 83052 237778
rect 77948 237500 83052 237542
rect 84204 237140 84524 238180
rect 77258 237098 80476 237140
rect 77258 236862 80198 237098
rect 80434 236862 80476 237098
rect 77258 236820 80476 236862
rect 83836 237098 84524 237140
rect 83836 236862 83878 237098
rect 84114 236862 84524 237098
rect 83836 236820 84524 236862
rect 87516 237098 87836 238222
rect 498756 238458 500548 238500
rect 498756 238222 498798 238458
rect 499034 238222 500270 238458
rect 500506 238222 500548 238458
rect 498756 238180 500548 238222
rect 500964 238458 501284 238500
rect 500964 238222 501006 238458
rect 501242 238222 501284 238458
rect 87516 236862 87558 237098
rect 87794 236862 87836 237098
rect 87516 236820 87836 236862
rect 500964 237098 501284 238222
rect 500964 236862 501006 237098
rect 501242 236862 501284 237098
rect 500964 236820 501284 236862
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 82364 235874 82730 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect 82364 235638 82452 235874
rect 82688 235638 82730 235874
rect 82364 235596 82730 235638
rect 82364 235100 82684 235596
rect 82364 234780 88066 235100
rect 498756 235058 501836 235100
rect 498756 234822 498798 235058
rect 499034 234822 501836 235058
rect 498756 234780 501836 234822
rect 82548 234378 87422 234420
rect 82548 234142 82590 234378
rect 82826 234142 87144 234378
rect 87380 234142 87422 234378
rect 82548 234100 87422 234142
rect 87746 233740 88066 234780
rect 78132 233698 83236 233740
rect 78132 233462 78174 233698
rect 78410 233462 82958 233698
rect 83194 233462 83236 233698
rect 78132 233420 83236 233462
rect 83836 233420 88066 233740
rect 101500 234378 101820 234420
rect 101500 234142 101542 234378
rect 101778 234142 101820 234378
rect 83836 232380 84156 233420
rect 86228 233018 87652 233060
rect 86228 232782 86270 233018
rect 86506 232782 87374 233018
rect 87610 232782 87652 233018
rect 86228 232740 87652 232782
rect 82364 232338 84156 232380
rect 82364 232102 82406 232338
rect 82642 232102 84156 232338
rect 82364 232060 84156 232102
rect 86412 232338 87652 232380
rect 86412 232102 86454 232338
rect 86690 232102 87652 232338
rect 86412 232060 87652 232102
rect 82732 231658 86916 231700
rect 82732 231422 82774 231658
rect 83010 231422 86638 231658
rect 86874 231422 86916 231658
rect 82732 231380 86916 231422
rect 87332 231020 87652 232060
rect 88252 231658 88940 231700
rect 88252 231422 88294 231658
rect 88530 231422 88940 231658
rect 88252 231380 88940 231422
rect 77764 230978 87652 231020
rect 77764 230742 77806 230978
rect 78042 230742 87652 230978
rect 77764 230700 87652 230742
rect 82410 230298 86732 230340
rect 82410 230062 86454 230298
rect 86690 230062 86732 230298
rect 82410 230020 86732 230062
rect 82410 229618 82730 230020
rect 88620 229660 88940 231380
rect 101500 230298 101820 234142
rect 497284 234378 500732 234420
rect 497284 234142 500454 234378
rect 500690 234142 500732 234378
rect 497284 234100 500732 234142
rect 497284 232380 497604 234100
rect 498020 233018 498708 233060
rect 498020 232782 498062 233018
rect 498298 232782 498430 233018
rect 498666 232782 498708 233018
rect 498020 232740 498708 232782
rect 500044 233018 501100 233060
rect 500044 232782 500086 233018
rect 500322 232782 500822 233018
rect 501058 232782 501100 233018
rect 500044 232740 501100 232782
rect 501516 232380 501836 234780
rect 497284 232338 498156 232380
rect 497284 232102 497878 232338
rect 498114 232102 498156 232338
rect 497284 232060 498156 232102
rect 499308 232060 501836 232380
rect 499308 231700 499628 232060
rect 499308 231658 502388 231700
rect 499308 231422 502110 231658
rect 502346 231422 502388 231658
rect 499308 231380 502388 231422
rect 101500 230062 101542 230298
rect 101778 230062 101820 230298
rect 101500 230020 101820 230062
rect 82410 229382 82452 229618
rect 82688 229382 82730 229618
rect 82410 229340 82730 229382
rect 86228 229618 88940 229660
rect 86228 229382 86270 229618
rect 86506 229382 88940 229618
rect 86228 229340 88940 229382
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect 82364 228258 86548 228300
rect 82364 228022 82406 228258
rect 82642 228022 86548 228258
rect 82364 227980 86548 228022
rect 83836 227578 84340 227620
rect 83836 227342 83878 227578
rect 84114 227342 84340 227578
rect 83836 227300 84340 227342
rect 86228 227578 86548 227980
rect 86228 227342 86270 227578
rect 86506 227342 86548 227578
rect 86228 227300 86548 227342
rect 498388 227578 498708 227620
rect 498388 227342 498430 227578
rect 498666 227342 498708 227578
rect 84020 226668 84340 227300
rect 498388 226940 498708 227342
rect 498388 226898 500180 226940
rect 84020 226626 84524 226668
rect 84020 226390 84246 226626
rect 84482 226390 84524 226626
rect 498388 226662 499902 226898
rect 500138 226662 500180 226898
rect 498388 226620 500180 226662
rect 84020 226348 84524 226390
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect 82548 224178 86916 224220
rect 82548 223942 82590 224178
rect 82826 223942 86916 224178
rect 82548 223900 86916 223942
rect 86596 223498 86916 223900
rect 86596 223262 86638 223498
rect 86874 223262 86916 223498
rect 86596 223220 86916 223262
rect 499860 224178 500180 224220
rect 499860 223942 499902 224178
rect 500138 223942 500180 224178
rect 499860 223498 500180 223942
rect 499860 223262 499902 223498
rect 500138 223262 500180 223498
rect 499860 223220 500180 223262
rect 500780 223498 501100 223540
rect 500780 223262 500822 223498
rect 501058 223262 501100 223498
rect 500780 222860 501100 223262
rect 77764 222818 86180 222860
rect 77764 222582 77806 222818
rect 78042 222582 86180 222818
rect 77764 222540 86180 222582
rect 85860 222340 86180 222540
rect 86596 222818 86916 222860
rect 86596 222582 86638 222818
rect 86874 222582 86916 222818
rect 86596 222340 86916 222582
rect 498940 222818 501100 222860
rect 498940 222582 498982 222818
rect 499218 222582 501100 222818
rect 498940 222540 501100 222582
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 85860 222076 86916 222340
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect 497836 220778 499812 220820
rect 497836 220542 499534 220778
rect 499770 220542 499812 220778
rect 497836 220500 499812 220542
rect 77764 220098 84524 220140
rect 77764 219862 77806 220098
rect 78042 219862 84524 220098
rect 77764 219820 84524 219862
rect 82916 219418 83604 219460
rect 82916 219182 82958 219418
rect 83194 219182 83326 219418
rect 83562 219182 83604 219418
rect 82916 219140 83604 219182
rect 84204 219418 84524 219820
rect 84204 219182 84246 219418
rect 84482 219182 84524 219418
rect 84204 219140 84524 219182
rect 85308 219418 87652 219460
rect 85308 219182 87374 219418
rect 87610 219182 87652 219418
rect 85308 219140 87652 219182
rect 497836 219418 498156 220500
rect 499308 220098 501468 220140
rect 499308 219862 499350 220098
rect 499586 219862 501190 220098
rect 501426 219862 501468 220098
rect 499308 219820 501468 219862
rect 497836 219182 497878 219418
rect 498114 219182 498156 219418
rect 497836 219140 498156 219182
rect 499492 219418 504780 219460
rect 499492 219182 499534 219418
rect 499770 219182 504502 219418
rect 504738 219182 504780 219418
rect 499492 219140 504780 219182
rect 85308 218916 85628 219140
rect 84756 218780 85628 218916
rect 84388 218738 85628 218780
rect 84388 218502 84430 218738
rect 84666 218596 85628 218738
rect 84666 218502 85076 218596
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 84388 218476 85076 218502
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect 84020 217378 89676 217420
rect 84020 217142 84062 217378
rect 84298 217142 89676 217378
rect 84020 217100 89676 217142
rect 75924 216698 83972 216740
rect 75924 216462 75966 216698
rect 76202 216462 83694 216698
rect 83930 216462 83972 216698
rect 75924 216420 83972 216462
rect 84756 216698 88756 216740
rect 84756 216462 84798 216698
rect 85034 216462 88756 216698
rect 84756 216420 88756 216462
rect 77764 216018 84156 216060
rect 77764 215782 77806 216018
rect 78042 215782 83878 216018
rect 84114 215782 84156 216018
rect 77764 215740 84156 215782
rect 84756 216018 88020 216060
rect 84756 215782 84798 216018
rect 85034 215782 87742 216018
rect 87978 215782 88020 216018
rect 84756 215740 88020 215782
rect 88436 215380 88756 216420
rect 83468 215338 88756 215380
rect 83468 215102 83510 215338
rect 83746 215102 88756 215338
rect 83468 215060 88756 215102
rect 84388 214658 84708 214700
rect 84388 214422 84430 214658
rect 84666 214422 84708 214658
rect 84388 214020 84708 214422
rect 83284 213978 84708 214020
rect 83284 213742 83326 213978
rect 83562 213742 84708 213978
rect 83284 213700 84708 213742
rect 85124 214658 86548 214700
rect 85124 214422 86270 214658
rect 86506 214422 86548 214658
rect 85124 214380 86548 214422
rect 87516 214658 87836 214700
rect 87516 214422 87558 214658
rect 87794 214422 87836 214658
rect 85124 213340 85444 214380
rect 82732 213020 85444 213340
rect 87516 213340 87836 214422
rect 88252 214658 88940 214700
rect 88252 214422 88294 214658
rect 88530 214422 88940 214658
rect 88252 214380 88940 214422
rect 87516 213298 88204 213340
rect 87516 213062 87926 213298
rect 88162 213062 88204 213298
rect 87516 213020 88204 213062
rect 82732 212660 83052 213020
rect 88620 212660 88940 214380
rect 77764 212618 83052 212660
rect 77764 212382 77806 212618
rect 78042 212382 83052 212618
rect 77764 212340 83052 212382
rect 88206 212618 88940 212660
rect 88206 212382 88248 212618
rect 88484 212382 88940 212618
rect 88206 212340 88940 212382
rect 89356 211980 89676 217100
rect 497468 217378 497788 217420
rect 497468 217142 497510 217378
rect 497746 217142 497788 217378
rect 497468 216740 497788 217142
rect 497468 216420 499076 216740
rect 90460 215338 90964 215380
rect 90460 215102 90502 215338
rect 90738 215102 90964 215338
rect 90460 215060 90964 215102
rect 90644 213978 90964 215060
rect 90644 213742 90686 213978
rect 90922 213742 90964 213978
rect 90644 213700 90964 213742
rect 498756 212618 499076 216420
rect 499492 216698 499812 216740
rect 499492 216462 499534 216698
rect 499770 216462 499812 216698
rect 499492 214020 499812 216462
rect 500228 215338 501284 215380
rect 500228 215102 500270 215338
rect 500506 215102 501006 215338
rect 501242 215102 501284 215338
rect 500228 215060 501284 215102
rect 504460 215338 504780 215380
rect 504460 215102 504502 215338
rect 504738 215102 504780 215338
rect 504460 214700 504780 215102
rect 500228 214658 504780 214700
rect 500228 214422 500270 214658
rect 500506 214422 504780 214658
rect 500228 214380 504780 214422
rect 499492 213978 500364 214020
rect 499492 213742 500086 213978
rect 500322 213742 500364 213978
rect 499492 213700 500364 213742
rect 498756 212382 498798 212618
rect 499034 212382 499076 212618
rect 498756 212340 499076 212382
rect 84572 211938 89676 211980
rect 84572 211702 84614 211938
rect 84850 211702 89676 211938
rect 84572 211660 89676 211702
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect 84572 210578 86916 210620
rect 84572 210342 84614 210578
rect 84850 210342 86638 210578
rect 86874 210342 86916 210578
rect 84572 210300 86916 210342
rect 84756 209898 85076 209940
rect 84756 209662 84798 209898
rect 85034 209662 85076 209898
rect 84756 209260 85076 209662
rect 498756 209898 499444 209940
rect 498756 209662 498798 209898
rect 499034 209662 499166 209898
rect 499402 209662 499444 209898
rect 498756 209620 499444 209662
rect 82364 209218 85076 209260
rect 82364 208982 82406 209218
rect 82642 208982 85076 209218
rect 82364 208940 85076 208982
rect 498756 209218 499812 209260
rect 498756 208982 498798 209218
rect 499034 208982 499534 209218
rect 499770 208982 499812 209218
rect 498756 208940 499812 208982
rect 77396 208538 86180 208580
rect 77396 208302 77438 208538
rect 77674 208302 85902 208538
rect 86138 208302 86180 208538
rect 77396 208260 86180 208302
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect 82916 206498 83972 206540
rect 82916 206262 82958 206498
rect 83194 206262 83694 206498
rect 83930 206262 83972 206498
rect 82916 206220 83972 206262
rect 85860 206498 87652 206540
rect 85860 206262 85902 206498
rect 86138 206362 87652 206498
rect 86138 206262 87374 206362
rect 85860 206220 87374 206262
rect 87332 206126 87374 206220
rect 87610 206126 87652 206362
rect 87332 206084 87652 206126
rect 78132 205818 85444 205860
rect 78132 205582 78174 205818
rect 78410 205582 85166 205818
rect 85402 205582 85444 205818
rect 78132 205540 85444 205582
rect 86228 205818 86916 205860
rect 86228 205582 86270 205818
rect 86506 205582 86638 205818
rect 86874 205582 86916 205818
rect 86228 205540 86916 205582
rect 498204 205818 499812 205860
rect 498204 205582 498246 205818
rect 498482 205582 499534 205818
rect 499770 205582 499812 205818
rect 498204 205540 499812 205582
rect 84204 205138 85812 205180
rect 84204 204902 84246 205138
rect 84482 204902 85534 205138
rect 85770 204902 85812 205138
rect 84204 204860 85812 204902
rect 86780 205138 88020 205180
rect 86780 204902 86822 205138
rect 87058 204902 87742 205138
rect 87978 204902 88020 205138
rect 86780 204860 88020 204902
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect 78132 203098 102556 203140
rect 78132 202862 78174 203098
rect 78410 202862 102556 203098
rect 78132 202820 102556 202862
rect 84756 202418 85444 202460
rect 84756 202182 84798 202418
rect 85034 202182 85444 202418
rect 84756 202140 85444 202182
rect 85860 202418 87468 202460
rect 85860 202182 85902 202418
rect 86138 202182 87190 202418
rect 87426 202182 87468 202418
rect 85860 202140 87468 202182
rect 85124 201738 85444 202140
rect 102236 201780 102556 202820
rect 169580 202820 179468 203140
rect 169580 201780 169900 202820
rect 85124 201502 85166 201738
rect 85402 201502 85444 201738
rect 85124 201460 85444 201502
rect 85860 201738 88020 201780
rect 85860 201502 85902 201738
rect 86138 201502 87742 201738
rect 87978 201502 88020 201738
rect 85860 201460 88020 201502
rect 102236 201460 169900 201780
rect 179148 201780 179468 202820
rect 208220 202820 218108 203140
rect 187060 202140 189956 202460
rect 187060 201780 187380 202140
rect 179148 201460 187380 201780
rect 189636 201780 189956 202140
rect 208220 201780 208540 202820
rect 189636 201460 208540 201780
rect 217788 201780 218108 202820
rect 227540 202820 237428 203140
rect 227540 201780 227860 202820
rect 217788 201460 227860 201780
rect 237108 201780 237428 202820
rect 246860 202820 256748 203140
rect 246860 201780 247180 202820
rect 237108 201460 247180 201780
rect 256428 201780 256748 202820
rect 266180 202820 276068 203140
rect 266180 201780 266500 202820
rect 256428 201460 266500 201780
rect 275748 201780 276068 202820
rect 285500 202820 295388 203140
rect 285500 201780 285820 202820
rect 275748 201460 285820 201780
rect 295068 201780 295388 202820
rect 304820 202820 314708 203140
rect 304820 201780 305140 202820
rect 295068 201460 305140 201780
rect 314388 201780 314708 202820
rect 324140 202820 334028 203140
rect 324140 201780 324460 202820
rect 314388 201460 324460 201780
rect 333708 201780 334028 202820
rect 339412 202820 346724 203140
rect 339412 201780 339732 202820
rect 333708 201460 339732 201780
rect 346404 201780 346724 202820
rect 394980 202820 403948 203140
rect 394980 201780 395300 202820
rect 346404 201460 395300 201780
rect 403628 201780 403948 202820
rect 414300 202820 423268 203140
rect 414300 201780 414620 202820
rect 403628 201460 414620 201780
rect 422948 201780 423268 202820
rect 433620 202820 442588 203140
rect 433620 201780 433940 202820
rect 422948 201460 433940 201780
rect 442268 201780 442588 202820
rect 452940 202820 461908 203140
rect 452940 201780 453260 202820
rect 442268 201460 453260 201780
rect 461588 201780 461908 202820
rect 472260 202820 480492 203140
rect 499124 203098 501468 203140
rect 499124 202862 499166 203098
rect 499402 202862 501190 203098
rect 501426 202862 501468 203098
rect 499124 202820 501468 202862
rect 472260 201780 472580 202820
rect 461588 201460 472580 201780
rect 480172 201780 480492 202820
rect 493236 202140 498156 202460
rect 493236 201780 493556 202140
rect 480172 201460 493556 201780
rect 497836 201780 498156 202140
rect 499124 202418 501284 202460
rect 499124 202182 501006 202418
rect 501242 202182 501284 202418
rect 499124 202140 501284 202182
rect 499124 201780 499444 202140
rect 497836 201460 499444 201780
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect 101316 199698 101636 199740
rect 101316 199462 101358 199698
rect 101594 199462 101636 199698
rect 84756 199018 86180 199060
rect 84756 198782 84798 199018
rect 85034 198782 85902 199018
rect 86138 198782 86180 199018
rect 84756 198740 86180 198782
rect 82548 196978 86916 197020
rect 82548 196742 82590 196978
rect 82826 196742 86638 196978
rect 86874 196742 86916 196978
rect 82548 196700 86916 196742
rect 101316 196340 101636 199462
rect 499676 199018 500916 199060
rect 499676 198782 499718 199018
rect 499954 198782 500638 199018
rect 500874 198782 500916 199018
rect 499676 198740 500916 198782
rect 497468 197658 498708 197700
rect 497468 197422 498430 197658
rect 498666 197422 498708 197658
rect 497468 197380 498708 197422
rect 83100 196298 84892 196340
rect 83100 196062 83142 196298
rect 83378 196062 84614 196298
rect 84850 196062 84892 196298
rect 83100 196020 84892 196062
rect 87700 196298 88020 196340
rect 87700 196062 87742 196298
rect 87978 196062 88020 196298
rect 87700 195660 88020 196062
rect 101316 196298 101820 196340
rect 101316 196062 101542 196298
rect 101778 196062 101820 196298
rect 101316 196020 101820 196062
rect 77948 195618 83052 195660
rect 77948 195382 77990 195618
rect 78226 195382 82774 195618
rect 83010 195382 83052 195618
rect 77948 195340 83052 195382
rect 86228 195618 88020 195660
rect 86228 195382 86270 195618
rect 86506 195382 88020 195618
rect 86228 195340 88020 195382
rect 82732 194938 84524 194980
rect 82732 194702 82774 194938
rect 83010 194702 84246 194938
rect 84482 194702 84524 194938
rect 82732 194660 84524 194702
rect 77396 194258 83052 194300
rect 77396 194022 77438 194258
rect 77674 194022 82774 194258
rect 83010 194022 83052 194258
rect 77396 193980 83052 194022
rect 83468 194258 86916 194300
rect 83468 194022 83510 194258
rect 83746 194022 86638 194258
rect 86874 194022 86916 194258
rect 83468 193980 86916 194022
rect 497468 194258 497788 197380
rect 498388 196978 500364 197020
rect 498388 196742 500086 196978
rect 500322 196742 500364 196978
rect 498388 196700 500364 196742
rect 498388 195618 498708 196700
rect 498388 195382 498430 195618
rect 498666 195382 498708 195618
rect 498388 195340 498708 195382
rect 500044 195618 500364 195660
rect 500044 195382 500086 195618
rect 500322 195382 500364 195618
rect 500044 194980 500364 195382
rect 500044 194938 501652 194980
rect 500044 194702 501374 194938
rect 501610 194702 501652 194938
rect 500044 194660 501652 194702
rect 497468 194022 497510 194258
rect 497746 194022 497788 194258
rect 497468 193980 497788 194022
rect 500044 194258 501652 194300
rect 500044 194022 500086 194258
rect 500322 194022 501374 194258
rect 501610 194022 501652 194258
rect 500044 193980 501652 194022
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect 83836 192218 86916 192260
rect 83836 191982 83878 192218
rect 84114 191982 86638 192218
rect 86874 191982 86916 192218
rect 83836 191940 86916 191982
rect 88068 192218 89308 192260
rect 88068 191982 88110 192218
rect 88346 191982 89308 192218
rect 88068 191940 89308 191982
rect 77764 191538 83788 191580
rect 77764 191302 77806 191538
rect 78042 191302 83510 191538
rect 83746 191302 83788 191538
rect 77764 191260 83788 191302
rect 84204 191538 88572 191580
rect 84204 191302 84246 191538
rect 84482 191302 88572 191538
rect 84204 191260 88572 191302
rect 82364 190858 85076 190900
rect 82364 190622 82406 190858
rect 82642 190622 84798 190858
rect 85034 190622 85076 190858
rect 82364 190580 85076 190622
rect 88252 190858 88572 191260
rect 88252 190622 88294 190858
rect 88530 190622 88572 190858
rect 88252 190580 88572 190622
rect 88988 190220 89308 191940
rect 499860 191538 500180 191580
rect 499860 191302 499902 191538
rect 500138 191302 500180 191538
rect 499860 190900 500180 191302
rect 499308 190858 500180 190900
rect 499308 190622 499350 190858
rect 499586 190622 500180 190858
rect 499308 190580 500180 190622
rect 88068 190178 89308 190220
rect 88068 189942 88110 190178
rect 88346 189942 89308 190178
rect 88068 189900 89308 189942
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect 82548 188138 85076 188180
rect 82548 187902 82590 188138
rect 82826 187902 84798 188138
rect 85034 187902 85076 188138
rect 82548 187860 85076 187902
rect 83652 187458 88204 187500
rect 83652 187222 83694 187458
rect 83930 187222 87926 187458
rect 88162 187222 88204 187458
rect 83652 187180 88204 187222
rect 83836 186778 84892 186820
rect 83836 186542 83878 186778
rect 84114 186542 84614 186778
rect 84850 186542 84892 186778
rect 83836 186500 84892 186542
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect 77396 184738 85444 184780
rect 77396 184502 77438 184738
rect 77674 184502 85444 184738
rect 77396 184460 85444 184502
rect 77764 184058 82132 184100
rect 77764 183822 77806 184058
rect 78042 183822 82132 184058
rect 77764 183780 82132 183822
rect 81812 183420 82132 183780
rect 85124 183420 85444 184460
rect 81812 183378 83604 183420
rect 81812 183142 83326 183378
rect 83562 183142 83604 183378
rect 81812 183100 83604 183142
rect 84388 183378 85444 183420
rect 84388 183142 84430 183378
rect 84666 183142 85444 183378
rect 84388 183100 85444 183142
rect 498204 183378 499996 183420
rect 498204 183142 498246 183378
rect 498482 183142 499718 183378
rect 499954 183142 499996 183378
rect 498204 183100 499996 183142
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect 82548 181338 86916 181380
rect 82548 181102 86638 181338
rect 86874 181102 86916 181338
rect 82548 181060 86916 181102
rect 90276 181338 90780 181380
rect 90276 181102 90502 181338
rect 90738 181102 90780 181338
rect 90276 181060 90780 181102
rect 82548 179298 82868 181060
rect 86596 180658 87284 180700
rect 86596 180422 86638 180658
rect 86874 180422 87006 180658
rect 87242 180422 87284 180658
rect 86596 180380 87284 180422
rect 82548 179062 82590 179298
rect 82826 179062 82868 179298
rect 82548 179020 82868 179062
rect 83284 179978 83604 180020
rect 83284 179742 83326 179978
rect 83562 179742 83604 179978
rect 83284 178618 83604 179742
rect 84020 179978 87468 180020
rect 84020 179742 84062 179978
rect 84298 179742 87468 179978
rect 84020 179700 87468 179742
rect 83284 178382 83326 178618
rect 83562 178382 83604 178618
rect 83284 178340 83604 178382
rect 84204 179298 84524 179340
rect 84204 179062 84246 179298
rect 84482 179062 84524 179298
rect 77764 177258 83788 177300
rect 77764 177022 77806 177258
rect 78042 177022 83510 177258
rect 83746 177022 83788 177258
rect 77764 176980 83788 177022
rect 84204 176620 84524 179062
rect 78132 176578 84524 176620
rect 78132 176342 78174 176578
rect 78410 176342 84524 176578
rect 78132 176300 84524 176342
rect 87148 176578 87468 179700
rect 90276 178660 90596 181060
rect 101500 179978 102004 180020
rect 101500 179742 101726 179978
rect 101962 179742 102004 179978
rect 101500 179700 102004 179742
rect 497652 179978 499076 180020
rect 497652 179742 498798 179978
rect 499034 179742 499076 179978
rect 497652 179700 499076 179742
rect 101500 179340 101820 179700
rect 101132 179020 101820 179340
rect 90276 178618 90964 178660
rect 90276 178382 90686 178618
rect 90922 178382 90964 178618
rect 90276 178340 90964 178382
rect 101132 177980 101452 179020
rect 101132 177938 101820 177980
rect 101132 177702 101542 177938
rect 101778 177702 101820 177938
rect 101132 177660 101820 177702
rect 87884 177258 88940 177300
rect 87884 177022 87926 177258
rect 88162 177022 88940 177258
rect 87884 176980 88940 177022
rect 87148 176342 87190 176578
rect 87426 176342 87468 176578
rect 87148 176300 87468 176342
rect 88620 175940 88940 176980
rect 497652 176620 497972 179700
rect 498572 178618 499260 178660
rect 498572 178382 498982 178618
rect 499218 178382 499260 178618
rect 498572 178340 499260 178382
rect 500412 178618 500732 178660
rect 500412 178382 500454 178618
rect 500690 178382 500732 178618
rect 498572 177980 498892 178340
rect 498572 177938 499996 177980
rect 498572 177702 499718 177938
rect 499954 177702 499996 177938
rect 498572 177660 499996 177702
rect 500412 177300 500732 178382
rect 500228 177258 500732 177300
rect 500228 177022 500270 177258
rect 500506 177022 500732 177258
rect 500228 176980 500732 177022
rect 497652 176300 499260 176620
rect 87148 175898 88940 175940
rect 87148 175662 87190 175898
rect 87426 175662 88940 175898
rect 87148 175620 88940 175662
rect 498940 175898 499260 176300
rect 498940 175662 498982 175898
rect 499218 175662 499260 175898
rect 498940 175620 499260 175662
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect 87194 174538 87514 174580
rect 87194 174302 87236 174538
rect 87472 174302 87514 174538
rect 87194 173900 87514 174302
rect 87194 173580 88020 173900
rect 85676 173178 87284 173220
rect 85676 172942 87006 173178
rect 87242 172942 87284 173178
rect 85676 172900 87284 172942
rect 85676 172540 85996 172900
rect 87700 172540 88020 173580
rect 88942 173858 89262 173900
rect 88942 173622 88984 173858
rect 89220 173622 89262 173858
rect 88942 172540 89262 173622
rect 498572 173858 500548 173900
rect 498572 173622 498614 173858
rect 498850 173622 500270 173858
rect 500506 173622 500548 173858
rect 498572 173580 500548 173622
rect 83284 172498 85996 172540
rect 83284 172262 83326 172498
rect 83562 172262 85996 172498
rect 83284 172220 85996 172262
rect 87194 172498 88020 172540
rect 87194 172262 87236 172498
rect 87472 172262 88020 172498
rect 87194 172220 88020 172262
rect 88620 172498 89262 172540
rect 88620 172262 88662 172498
rect 88898 172262 89262 172498
rect 88620 172220 89262 172262
rect 498204 172498 499628 172540
rect 498204 172262 498246 172498
rect 498482 172262 499350 172498
rect 499586 172262 499628 172498
rect 498204 172220 499628 172262
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect 499308 170594 499628 170636
rect 83836 170458 86916 170500
rect 83836 170222 83878 170458
rect 84114 170222 86916 170458
rect 83836 170180 86916 170222
rect 88252 170458 89676 170500
rect 88252 170222 88294 170458
rect 88530 170222 89676 170458
rect 88252 170180 89676 170222
rect 90460 170458 90964 170500
rect 90460 170222 90502 170458
rect 90738 170222 90964 170458
rect 90460 170180 90964 170222
rect 499308 170358 499350 170594
rect 499586 170500 499628 170594
rect 499586 170358 500916 170500
rect 499308 170180 500916 170358
rect 84020 169778 84340 169820
rect 84020 169542 84062 169778
rect 84298 169542 84340 169778
rect 84020 169140 84340 169542
rect 78132 169098 84340 169140
rect 78132 168862 78174 169098
rect 78410 168862 84340 169098
rect 78132 168820 84340 168862
rect 86596 169098 86916 170180
rect 86596 168862 86638 169098
rect 86874 168862 86916 169098
rect 86596 168820 86916 168862
rect 87516 169778 88940 169820
rect 87516 169542 88662 169778
rect 88898 169542 88940 169778
rect 87516 169500 88940 169542
rect 87516 168460 87836 169500
rect 89356 169140 89676 170180
rect 90644 169778 90964 170180
rect 90644 169542 90686 169778
rect 90922 169542 90964 169778
rect 90644 169500 90964 169542
rect 500596 169778 500916 170180
rect 500596 169542 500638 169778
rect 500874 169542 500916 169778
rect 500596 169500 500916 169542
rect 88574 169098 89676 169140
rect 88574 168862 88616 169098
rect 88852 168862 89676 169098
rect 88574 168820 89676 168862
rect 498204 169098 499444 169140
rect 498204 168862 498246 169098
rect 498482 168862 499166 169098
rect 499402 168862 499444 169098
rect 498204 168820 499444 168862
rect 87378 168418 87836 168460
rect 87378 168182 87420 168418
rect 87656 168182 87836 168418
rect 87378 168140 87836 168182
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect 78132 167058 84524 167100
rect 78132 166822 78174 167058
rect 78410 166822 84246 167058
rect 84482 166822 84524 167058
rect 78132 166780 84524 166822
rect 498020 167058 500916 167100
rect 498020 166822 498062 167058
rect 498298 166822 500638 167058
rect 500874 166822 500916 167058
rect 498020 166780 500916 166822
rect 86964 166378 87698 166420
rect 86964 166142 87420 166378
rect 87656 166142 87698 166378
rect 86964 166100 87698 166142
rect 88436 166378 88756 166420
rect 88436 166142 88478 166378
rect 88714 166142 88756 166378
rect 78132 165698 84156 165740
rect 78132 165462 78174 165698
rect 78410 165462 83878 165698
rect 84114 165462 84156 165698
rect 78132 165420 84156 165462
rect 86964 165060 87284 166100
rect 88436 165698 88756 166142
rect 88436 165462 88478 165698
rect 88714 165462 88756 165698
rect 88436 165420 88756 165462
rect 499676 165698 500916 165740
rect 499676 165462 499718 165698
rect 499954 165462 500638 165698
rect 500874 165462 500916 165698
rect 499676 165420 500916 165462
rect 86964 165018 87422 165060
rect 86964 164782 87144 165018
rect 87380 164782 87422 165018
rect 86964 164740 87422 164782
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect 86228 163658 86548 163700
rect 86228 163422 86270 163658
rect 86506 163422 86548 163658
rect 77764 162978 83972 163020
rect 77764 162742 77806 162978
rect 78042 162742 83694 162978
rect 83930 162742 83972 162978
rect 77764 162700 83972 162742
rect 86228 161660 86548 163422
rect 87516 163658 87836 163700
rect 87516 163422 87558 163658
rect 87794 163422 87836 163658
rect 87516 162340 87836 163422
rect 88574 163658 88894 163700
rect 88574 163422 88616 163658
rect 88852 163422 88894 163658
rect 87516 162020 88204 162340
rect 88574 162298 88894 163422
rect 499308 162978 499996 163020
rect 499308 162742 499350 162978
rect 499586 162742 499996 162978
rect 499308 162700 499996 162742
rect 88574 162062 88616 162298
rect 88852 162062 88894 162298
rect 88574 162020 88894 162062
rect 86228 161618 87468 161660
rect 86228 161382 87190 161618
rect 87426 161382 87468 161618
rect 86228 161340 87468 161382
rect 87884 160980 88204 162020
rect 84204 160938 84708 160980
rect 84204 160702 84246 160938
rect 84482 160702 84708 160938
rect 84204 160660 84708 160702
rect 78132 158898 83972 158940
rect 78132 158662 78174 158898
rect 78410 158662 83694 158898
rect 83930 158662 83972 158898
rect 78132 158620 83972 158662
rect 84388 158260 84708 160660
rect 87332 160660 88204 160980
rect 499676 160938 499996 162700
rect 499676 160702 499718 160938
rect 499954 160702 499996 160938
rect 499676 160660 499996 160702
rect 87332 160258 87652 160660
rect 87332 160022 87374 160258
rect 87610 160022 87652 160258
rect 87332 159980 87652 160022
rect 83836 158218 84708 158260
rect 83836 157982 83878 158218
rect 84114 157982 84708 158218
rect 83836 157940 84708 157982
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect 498388 156178 499996 156220
rect 498388 155942 499718 156178
rect 499954 155942 499996 156178
rect 498388 155900 499996 155942
rect 498388 155540 498708 155900
rect 77764 155498 83972 155540
rect 77764 155262 77806 155498
rect 78042 155262 83694 155498
rect 83930 155262 83972 155498
rect 77764 155220 83972 155262
rect 498388 155498 499996 155540
rect 498388 155262 499718 155498
rect 499954 155262 499996 155498
rect 498388 155220 499996 155262
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect 78132 152098 83788 152140
rect 78132 151862 78174 152098
rect 78410 151862 83510 152098
rect 83746 151862 83788 152098
rect 78132 151820 83788 151862
rect 77764 150738 83788 150780
rect 77764 150502 77806 150738
rect 78042 150502 83510 150738
rect 83746 150502 83788 150738
rect 77764 150460 83788 150502
rect 499308 150738 500548 150780
rect 499308 150502 499350 150738
rect 499586 150502 500270 150738
rect 500506 150502 500548 150738
rect 499308 150460 500548 150502
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect 499124 148970 499444 149012
rect 497652 148698 498340 148740
rect 497652 148462 498062 148698
rect 498298 148462 498340 148698
rect 497652 148420 498340 148462
rect 499124 148734 499166 148970
rect 499402 148740 499444 148970
rect 499402 148734 500548 148740
rect 499124 148698 500548 148734
rect 499124 148462 500270 148698
rect 500506 148462 500548 148698
rect 499124 148420 500548 148462
rect 497652 147380 497972 148420
rect 498388 148018 499628 148060
rect 498388 147782 498430 148018
rect 498666 147782 499350 148018
rect 499586 147782 499628 148018
rect 498388 147740 499628 147782
rect 497652 147338 498524 147380
rect 497652 147102 498246 147338
rect 498482 147102 498524 147338
rect 497652 147060 498524 147102
rect 499860 147338 501284 147380
rect 499860 147102 499902 147338
rect 500138 147102 501006 147338
rect 501242 147102 501284 147338
rect 499860 147060 501284 147102
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect 498204 145298 499490 145340
rect 498204 145062 498246 145298
rect 498482 145062 499212 145298
rect 499448 145062 499490 145298
rect 498204 145020 499490 145062
rect 499860 145298 500916 145340
rect 499860 145062 499902 145298
rect 500138 145062 500638 145298
rect 500874 145062 500916 145298
rect 499860 145020 500916 145062
rect 84020 144618 84892 144660
rect 84020 144382 84062 144618
rect 84298 144382 84892 144618
rect 84020 144340 84892 144382
rect 498572 144618 500180 144660
rect 498572 144382 498614 144618
rect 498850 144382 499902 144618
rect 500138 144382 500180 144618
rect 498572 144340 500180 144382
rect 78132 141898 83972 141940
rect 78132 141662 78174 141898
rect 78410 141662 83694 141898
rect 83930 141662 83972 141898
rect 78132 141620 83972 141662
rect 83468 141218 84156 141260
rect 83468 140982 83878 141218
rect 84114 140982 84156 141218
rect 83468 140940 84156 140982
rect 83468 140538 83788 140940
rect 84572 140580 84892 144340
rect 86964 143938 87284 143980
rect 86964 143702 87006 143938
rect 87242 143702 87284 143938
rect 86964 142578 87284 143702
rect 86964 142342 87006 142578
rect 87242 142342 87284 142578
rect 86964 142300 87284 142342
rect 83468 140302 83510 140538
rect 83746 140302 83788 140538
rect 83468 140260 83788 140302
rect 84204 140538 84892 140580
rect 84204 140302 84246 140538
rect 84482 140302 84892 140538
rect 84204 140260 84892 140302
rect 498940 140538 499628 140580
rect 498940 140302 498982 140538
rect 499218 140302 499350 140538
rect 499586 140302 499628 140538
rect 498940 140260 499628 140302
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect 86596 137818 86916 137860
rect 86596 137582 86638 137818
rect 86874 137582 86916 137818
rect 86596 137180 86916 137582
rect 86596 137138 87284 137180
rect 86596 136902 87006 137138
rect 87242 136902 87284 137138
rect 86596 136860 87284 136902
rect 499860 137138 501468 137180
rect 499860 136902 499902 137138
rect 500138 136902 501190 137138
rect 501426 136902 501468 137138
rect 499860 136860 501468 136902
rect 499170 136458 501100 136500
rect 499170 136222 499212 136458
rect 499448 136222 500822 136458
rect 501058 136222 501100 136458
rect 499170 136180 501100 136222
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect 497652 134418 499490 134460
rect 497652 134182 499212 134418
rect 499448 134182 499490 134418
rect 497652 134140 499490 134182
rect 497652 133100 497972 134140
rect 498388 133738 499490 133780
rect 498388 133502 498430 133738
rect 498666 133502 499212 133738
rect 499448 133502 499490 133738
rect 498388 133460 499490 133502
rect 84204 133058 86916 133100
rect 84204 132822 84246 133058
rect 84482 132822 86638 133058
rect 86874 132822 86916 133058
rect 84204 132780 86916 132822
rect 497652 133058 498340 133100
rect 497652 132822 498062 133058
rect 498298 132822 498340 133058
rect 497652 132780 498340 132822
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect 77396 131018 84156 131060
rect 77396 130782 77438 131018
rect 77674 130782 83878 131018
rect 84114 130782 84156 131018
rect 77396 130740 84156 130782
rect 498388 131018 499490 131060
rect 498388 130782 498430 131018
rect 498666 130782 499212 131018
rect 499448 130782 499490 131018
rect 498388 130740 499490 130782
rect 499860 131018 500364 131060
rect 499860 130782 499902 131018
rect 500138 130782 500364 131018
rect 499860 130740 500364 130782
rect 77396 130338 83788 130380
rect 77396 130102 77438 130338
rect 77674 130102 83510 130338
rect 83746 130102 83788 130338
rect 77396 130060 83788 130102
rect 500044 129700 500364 130740
rect 78132 129658 84340 129700
rect 78132 129422 78174 129658
rect 78410 129422 84062 129658
rect 84298 129422 84340 129658
rect 78132 129380 84340 129422
rect 499308 129658 500364 129700
rect 499308 129422 499350 129658
rect 499586 129422 500364 129658
rect 499308 129380 500364 129422
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect 201412 125980 203388 126300
rect 201412 124940 201732 125980
rect 203068 124940 203388 125980
rect 108308 124620 109364 124940
rect 108308 122900 108628 124620
rect 99108 122858 108628 122900
rect 99108 122622 99150 122858
rect 99386 122622 108628 122858
rect 99108 122580 108628 122622
rect 109044 122900 109364 124620
rect 185956 124620 201732 124940
rect 202700 124620 203388 124940
rect 224596 124620 229148 124940
rect 185956 123580 186276 124620
rect 202700 124260 203020 124620
rect 202700 123940 210012 124260
rect 176020 123538 186276 123580
rect 176020 123302 176062 123538
rect 176298 123302 186276 123538
rect 176020 123260 186276 123302
rect 209692 123538 210012 123940
rect 224596 123580 224916 124620
rect 209692 123302 209734 123538
rect 209970 123302 210012 123538
rect 209692 123260 210012 123302
rect 219076 123538 224916 123580
rect 219076 123302 219118 123538
rect 219354 123302 224916 123538
rect 219076 123260 224916 123302
rect 228828 123580 229148 124620
rect 371796 124620 381684 124940
rect 371796 124260 372116 124620
rect 235084 123940 240372 124260
rect 228828 123538 234300 123580
rect 228828 123302 234022 123538
rect 234258 123302 234300 123538
rect 228828 123260 234300 123302
rect 235084 123538 235404 123940
rect 235084 123302 235126 123538
rect 235362 123302 235404 123538
rect 235084 123260 235404 123302
rect 240052 123538 240372 123940
rect 240052 123302 240094 123538
rect 240330 123302 240372 123538
rect 240052 123260 240372 123302
rect 252932 123940 258220 124260
rect 252932 123538 253252 123940
rect 252932 123302 252974 123538
rect 253210 123302 253252 123538
rect 252932 123260 253252 123302
rect 257900 123538 258220 123940
rect 272988 123940 289132 124260
rect 272988 123716 273308 123940
rect 272436 123580 273308 123716
rect 257900 123302 257942 123538
rect 258178 123302 258220 123538
rect 257900 123260 258220 123302
rect 259924 123538 273308 123580
rect 259924 123302 259966 123538
rect 260202 123396 273308 123538
rect 288812 123580 289132 123940
rect 302060 123940 315996 124260
rect 302060 123580 302380 123940
rect 260202 123302 272756 123396
rect 259924 123260 272756 123302
rect 288812 123260 302380 123580
rect 315676 123580 315996 123940
rect 321564 123940 331452 124260
rect 321564 123580 321884 123940
rect 315676 123260 321884 123580
rect 331132 123580 331452 123940
rect 344932 123940 350772 124260
rect 344932 123580 345252 123940
rect 331132 123260 345252 123580
rect 350452 123580 350772 123940
rect 360020 123940 372116 124260
rect 381364 124260 381684 124620
rect 381364 123940 394196 124260
rect 360020 123580 360340 123940
rect 350452 123260 360340 123580
rect 393876 123580 394196 123940
rect 398660 123940 408732 124260
rect 398660 123580 398980 123940
rect 393876 123260 398980 123580
rect 408412 122900 408732 123940
rect 427732 123940 437620 124260
rect 427732 123580 428052 123940
rect 420004 123538 428052 123580
rect 420004 123302 420046 123538
rect 420282 123302 428052 123538
rect 420004 123260 428052 123302
rect 437300 123580 437620 123940
rect 447052 123940 466508 124260
rect 447052 123580 447372 123940
rect 437300 123260 447372 123580
rect 466188 123538 466508 123940
rect 466188 123302 466230 123538
rect 466466 123302 466508 123538
rect 466188 123260 466508 123302
rect 473916 123538 483252 123580
rect 473916 123302 473958 123538
rect 474194 123302 483252 123538
rect 473916 123260 483252 123302
rect 482932 123036 483252 123260
rect 485140 123538 496684 123580
rect 485140 123302 496406 123538
rect 496642 123302 496684 123538
rect 485140 123260 496684 123302
rect 497100 123538 498340 123580
rect 497100 123302 497142 123538
rect 497378 123302 498340 123538
rect 497100 123260 498340 123302
rect 482932 122900 483436 123036
rect 485140 122900 485460 123260
rect 498020 122900 498340 123260
rect 109044 122858 258772 122900
rect 109044 122622 258494 122858
rect 258730 122622 258772 122858
rect 109044 122580 258772 122622
rect 259188 122858 342492 122900
rect 259188 122622 259230 122858
rect 259466 122622 342214 122858
rect 342450 122622 342492 122858
rect 259188 122580 342492 122622
rect 350452 122580 360340 122900
rect 379156 122858 379844 122900
rect 379156 122622 379198 122858
rect 379434 122622 379844 122858
rect 379156 122580 379844 122622
rect 408412 122858 417748 122900
rect 408412 122622 417470 122858
rect 417706 122622 417748 122858
rect 408412 122580 417748 122622
rect 434356 122858 434860 122900
rect 434356 122622 434398 122858
rect 434634 122622 434860 122858
rect 434356 122580 434860 122622
rect 350452 122220 350772 122580
rect 148052 122178 157204 122220
rect 148052 121942 148094 122178
rect 148330 121948 157204 122178
rect 157620 122084 166588 122220
rect 167372 122084 176524 122220
rect 176940 122084 185908 122220
rect 186692 122084 195844 122220
rect 196260 122084 205228 122220
rect 206012 122178 215348 122220
rect 206012 122084 215070 122178
rect 157620 121948 215070 122084
rect 148330 121942 215070 121948
rect 215306 121942 215348 122178
rect 148052 121900 215348 121942
rect 215396 122178 224548 122220
rect 215396 121942 215438 122178
rect 215674 122084 224548 122178
rect 229196 122178 243684 122220
rect 229196 122084 243406 122178
rect 215674 121942 243406 122084
rect 243642 121942 243684 122178
rect 215396 121900 243684 121942
rect 259188 122178 273124 122220
rect 259188 121942 259230 122178
rect 259466 121948 273124 122178
rect 273540 122178 281404 122220
rect 273540 121948 281126 122178
rect 259466 121942 281126 121948
rect 281362 121942 281404 122178
rect 259188 121900 281404 121942
rect 293044 122178 301644 122220
rect 293044 121942 293086 122178
rect 293322 121942 301366 122178
rect 301602 121942 301644 122178
rect 293044 121900 301644 121942
rect 322484 122178 331268 122220
rect 322484 121942 322526 122178
rect 322762 121942 330990 122178
rect 331226 121942 331268 122178
rect 322484 121900 331268 121942
rect 344748 122178 350772 122220
rect 344748 121942 344790 122178
rect 345026 121942 350772 122178
rect 344748 121900 350772 121942
rect 360020 122220 360340 122580
rect 379524 122220 379844 122580
rect 360020 122178 370092 122220
rect 360020 121942 369814 122178
rect 370050 121942 370092 122178
rect 360020 121900 370092 121942
rect 379524 122178 398428 122220
rect 379524 121942 398150 122178
rect 398386 121942 398428 122178
rect 379524 121900 398428 121942
rect 399028 122178 425292 122220
rect 399028 121942 399070 122178
rect 399306 121942 425014 122178
rect 425250 121942 425292 122178
rect 399028 121900 425292 121942
rect 434540 122178 434860 122580
rect 434540 121942 434582 122178
rect 434818 121942 434860 122178
rect 434540 121900 434860 121942
rect 444108 122858 444428 122900
rect 444108 122622 444150 122858
rect 444386 122622 444428 122858
rect 444108 122220 444428 122622
rect 447052 122580 456940 122900
rect 447052 122220 447372 122580
rect 444108 121900 447372 122220
rect 456620 122220 456940 122580
rect 466372 122580 476260 122900
rect 482932 122716 485460 122900
rect 483116 122580 485460 122716
rect 495812 122858 498340 122900
rect 495812 122622 495854 122858
rect 496090 122622 498340 122858
rect 495812 122580 498340 122622
rect 501516 122858 510300 122900
rect 501516 122622 510022 122858
rect 510258 122622 510300 122858
rect 501516 122580 510300 122622
rect 466372 122220 466692 122580
rect 456620 121900 466692 122220
rect 475940 122220 476260 122580
rect 501516 122220 501836 122580
rect 475940 121900 501836 122220
rect 156884 121628 157940 121900
rect 166268 121764 167692 121900
rect 176204 121764 177260 121900
rect 185588 121764 187012 121900
rect 195524 121764 196580 121900
rect 204908 121764 206332 121900
rect 224228 121764 229516 121900
rect 272804 121628 273860 121900
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect 163876 120138 174684 120180
rect 163876 119902 163918 120138
rect 164154 119902 174406 120138
rect 174642 119902 174684 120138
rect 163876 119860 174684 119902
rect 190372 120138 193452 120180
rect 190372 119902 193174 120138
rect 193410 119902 193452 120138
rect 190372 119860 193452 119902
rect 229012 120138 251412 120180
rect 229012 119902 251134 120138
rect 251370 119902 251412 120138
rect 229012 119860 251412 119902
rect 282740 119860 297596 120180
rect 183196 118778 186460 118820
rect 183196 118542 183238 118778
rect 183474 118542 186182 118778
rect 186418 118542 186460 118778
rect 183196 118500 186460 118542
rect 190372 118778 190692 119860
rect 229012 119500 229332 119860
rect 282740 119500 283060 119860
rect 196444 119458 229332 119500
rect 196444 119222 196486 119458
rect 196722 119222 229332 119458
rect 196444 119180 229332 119222
rect 273540 119458 283060 119500
rect 273540 119222 273582 119458
rect 273818 119222 283060 119458
rect 273540 119180 283060 119222
rect 297276 119500 297596 119860
rect 302244 119860 316180 120180
rect 326716 120138 331452 120180
rect 326716 119902 326758 120138
rect 326994 119902 331174 120138
rect 331410 119902 331452 120138
rect 326716 119860 331452 119902
rect 344932 119860 355556 120180
rect 302244 119500 302564 119860
rect 297276 119180 302564 119500
rect 190372 118542 190414 118778
rect 190650 118542 190692 118778
rect 190372 118500 190692 118542
rect 265444 118778 269996 118820
rect 265444 118542 265486 118778
rect 265722 118542 269718 118778
rect 269954 118542 269996 118778
rect 265444 118500 269996 118542
rect 315860 118778 316180 119860
rect 344932 119500 345252 119860
rect 340516 119458 345252 119500
rect 340516 119222 340558 119458
rect 340794 119222 345252 119458
rect 340516 119180 345252 119222
rect 355236 119500 355556 119860
rect 360020 120138 376900 120180
rect 360020 119902 376622 120138
rect 376858 119902 376900 120138
rect 360020 119860 376900 119902
rect 434172 120138 446820 120180
rect 434172 119902 446542 120138
rect 446778 119902 446820 120138
rect 434172 119860 446820 119902
rect 466372 119860 476260 120180
rect 360020 119500 360340 119860
rect 355236 119180 360340 119500
rect 394428 119458 395088 119500
rect 394428 119222 394654 119458
rect 394890 119222 395088 119458
rect 394428 119180 395088 119222
rect 399396 119458 408732 119500
rect 399396 119222 399438 119458
rect 399674 119222 408454 119458
rect 408690 119222 408732 119458
rect 399396 119180 408732 119222
rect 422764 119458 425476 119500
rect 422764 119222 422806 119458
rect 423042 119222 425476 119458
rect 422764 119180 425476 119222
rect 434172 119458 434492 119860
rect 466372 119500 466692 119860
rect 434172 119222 434214 119458
rect 434450 119222 434492 119458
rect 434172 119180 434492 119222
rect 453492 119458 454180 119500
rect 453492 119222 453534 119458
rect 453770 119222 453902 119458
rect 454138 119222 454180 119458
rect 453492 119180 454180 119222
rect 457172 119458 466692 119500
rect 457172 119222 457214 119458
rect 457450 119222 466692 119458
rect 457172 119180 466692 119222
rect 475940 119500 476260 119860
rect 475940 119458 507172 119500
rect 475940 119222 506894 119458
rect 507130 119222 507172 119458
rect 475940 119180 507172 119222
rect 315860 118542 315902 118778
rect 316138 118542 316180 118778
rect 315860 118500 316180 118542
rect 394428 118778 394748 119180
rect 425156 118820 425476 119180
rect 394428 118542 394470 118778
rect 394706 118542 394748 118778
rect 394428 118500 394748 118542
rect 424972 118778 425476 118820
rect 424972 118542 425014 118778
rect 425250 118542 425476 118778
rect 424972 118500 425476 118542
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect 87930 106538 88572 106580
rect 87930 106302 88294 106538
rect 88530 106302 88572 106538
rect 87930 106260 88572 106302
rect 87930 105900 88250 106260
rect 87930 105858 88572 105900
rect 87930 105622 88294 105858
rect 88530 105622 88572 105858
rect 87930 105580 88572 105622
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect 89356 4260 106236 4580
rect 89356 3900 89676 4260
rect 77028 3858 89676 3900
rect 77028 3622 77070 3858
rect 77306 3622 89676 3858
rect 77028 3580 89676 3622
rect 105916 3220 106236 4260
rect 114012 4260 128500 4580
rect 114012 3220 114332 4260
rect 128180 3900 128500 4260
rect 147316 4538 164564 4580
rect 147316 4302 164286 4538
rect 164522 4302 164564 4538
rect 147316 4260 164564 4302
rect 181908 4538 216452 4580
rect 181908 4302 181950 4538
rect 182186 4302 216452 4538
rect 181908 4260 216452 4302
rect 147316 3900 147636 4260
rect 216132 3900 216452 4260
rect 128180 3580 147636 3900
rect 169028 3858 172660 3900
rect 169028 3622 169070 3858
rect 169306 3622 172382 3858
rect 172618 3622 172660 3858
rect 169028 3580 172660 3622
rect 215028 3220 215532 3900
rect 216132 3858 243868 3900
rect 216132 3622 243590 3858
rect 243826 3622 243868 3858
rect 216132 3580 243868 3622
rect 253668 3220 254172 4580
rect 273172 4538 292812 4580
rect 273172 4302 273214 4538
rect 273450 4302 292812 4538
rect 273172 4260 292812 4302
rect 292492 3900 292812 4260
rect 306292 4260 316180 4580
rect 306292 3900 306612 4260
rect 268756 3858 272940 3900
rect 268756 3622 268798 3858
rect 269034 3622 272662 3858
rect 272898 3622 272940 3858
rect 268756 3580 272940 3622
rect 282188 3444 283244 3764
rect 292492 3580 306612 3900
rect 315860 3900 316180 4260
rect 325612 4538 329428 4580
rect 325612 4302 329150 4538
rect 329386 4302 329428 4538
rect 325612 4260 329428 4302
rect 337756 4538 367332 4580
rect 337756 4302 337798 4538
rect 338034 4302 367054 4538
rect 367290 4302 367332 4538
rect 337756 4260 367332 4302
rect 385964 4538 396220 4580
rect 385964 4302 395942 4538
rect 396178 4302 396220 4538
rect 385964 4260 396220 4302
rect 405468 4538 415908 4580
rect 405468 4302 405510 4538
rect 405746 4302 415630 4538
rect 415866 4302 415908 4538
rect 405468 4260 415908 4302
rect 424788 4538 434860 4580
rect 424788 4302 424830 4538
rect 425066 4302 434582 4538
rect 434818 4302 434860 4538
rect 424788 4260 434860 4302
rect 443188 4538 443508 4580
rect 443188 4302 443230 4538
rect 443466 4444 443508 4538
rect 444108 4538 444612 4580
rect 444108 4444 444334 4538
rect 443466 4302 444334 4444
rect 444570 4302 444612 4538
rect 443188 4260 444612 4302
rect 462324 4538 495396 4580
rect 462324 4302 462366 4538
rect 462602 4302 495118 4538
rect 495354 4302 495396 4538
rect 462324 4260 495396 4302
rect 325612 3900 325932 4260
rect 385964 3900 386284 4260
rect 443188 4124 444428 4260
rect 315860 3580 325932 3900
rect 367564 3858 386284 3900
rect 367564 3622 367606 3858
rect 367842 3622 386284 3858
rect 367564 3580 386284 3622
rect 457356 3858 461172 3900
rect 457356 3622 457398 3858
rect 457634 3622 460894 3858
rect 461130 3622 461172 3858
rect 457356 3580 461172 3622
rect 519916 3858 521892 3900
rect 519916 3622 519958 3858
rect 520194 3622 521614 3858
rect 521850 3622 521892 3858
rect 519916 3580 521892 3622
rect 547884 3858 558140 3900
rect 547884 3622 557862 3858
rect 558098 3622 558140 3858
rect 547884 3580 558140 3622
rect 282188 3220 282508 3444
rect 105916 2900 114332 3220
rect 114748 3178 127948 3220
rect 114748 2942 114790 3178
rect 115026 2942 127670 3178
rect 127906 2942 127948 3178
rect 114748 2900 127948 2942
rect 128364 3178 147268 3220
rect 128364 2942 128406 3178
rect 128642 2942 146990 3178
rect 147226 2942 147268 3178
rect 128364 2900 147268 2942
rect 147684 3178 205228 3220
rect 147684 2942 147726 3178
rect 147962 2942 204950 3178
rect 205186 2942 205228 3178
rect 147684 2900 205228 2942
rect 205644 3178 243684 3220
rect 205644 2942 205686 3178
rect 205922 2942 243406 3178
rect 243642 2942 243684 3178
rect 205644 2900 243684 2942
rect 244100 3178 264660 3220
rect 244100 2942 244142 3178
rect 244378 2942 264382 3178
rect 264618 2942 264660 3178
rect 244100 2900 264660 2942
rect 267468 3178 282508 3220
rect 267468 2942 267510 3178
rect 267746 2942 282508 3178
rect 267468 2900 282508 2942
rect 282924 3220 283244 3444
rect 547884 3220 548204 3580
rect 282924 3178 302196 3220
rect 282924 2942 301918 3178
rect 302154 2942 302196 3178
rect 282924 2900 302196 2942
rect 306108 3178 316180 3220
rect 306108 2942 306150 3178
rect 306386 2942 315902 3178
rect 316138 2942 316180 3178
rect 306108 2900 316180 2942
rect 325428 3178 335500 3220
rect 325428 2942 325470 3178
rect 325706 2942 335222 3178
rect 335458 2942 335500 3178
rect 325428 2900 335500 2942
rect 340700 3178 378740 3220
rect 340700 2942 340742 3178
rect 340978 2942 378462 3178
rect 378698 2942 378740 3178
rect 340700 2900 378740 2942
rect 379524 3178 398428 3220
rect 379524 2942 379566 3178
rect 379802 2942 398150 3178
rect 398386 2942 398428 3178
rect 379524 2900 398428 2942
rect 398844 3178 417748 3220
rect 398844 2942 398886 3178
rect 399122 2942 417470 3178
rect 417706 2942 417748 3178
rect 398844 2900 417748 2942
rect 419084 3178 436332 3220
rect 419084 2942 419126 3178
rect 419362 2942 436054 3178
rect 436290 2942 436332 3178
rect 419084 2900 436332 2942
rect 437300 3178 451788 3220
rect 437300 2942 437342 3178
rect 437578 2942 451510 3178
rect 451746 2942 451788 3178
rect 437300 2900 451788 2942
rect 461220 3178 470740 3220
rect 461220 2942 461262 3178
rect 461498 2942 470462 3178
rect 470698 2942 470740 3178
rect 461220 2900 470740 2942
rect 485508 3178 498892 3220
rect 485508 2942 485550 3178
rect 485786 2942 498614 3178
rect 498850 2942 498892 3178
rect 485508 2900 498892 2942
rect 507588 3178 514164 3220
rect 507588 2942 507630 3178
rect 507866 2942 513886 3178
rect 514122 2942 514164 3178
rect 507588 2900 514164 2942
rect 530956 3178 548204 3220
rect 530956 2942 530998 3178
rect 531234 2942 548204 3178
rect 530956 2900 548204 2942
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use Ibtida_top_dffram_cv  mprj
timestamp 1607298761
transform 1 0 82000 0 1 122000
box 0 0 420000 460000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 4 analog_io[0]
port 1 nsew
rlabel metal3 s 583520 474996 584960 475236 4 analog_io[10]
port 2 nsew
rlabel metal3 s 583520 521916 584960 522156 4 analog_io[11]
port 3 nsew
rlabel metal3 s 583520 568836 584960 569076 4 analog_io[12]
port 4 nsew
rlabel metal3 s 583520 615756 584960 615996 4 analog_io[13]
port 5 nsew
rlabel metal3 s 583520 662676 584960 662916 4 analog_io[14]
port 6 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[16]
port 8 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[17]
port 9 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[18]
port 10 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 52716 584960 52956 4 analog_io[1]
port 12 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[20]
port 13 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[21]
port 14 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[22]
port 15 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 21 nsew
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 22 nsew
rlabel metal3 s 583520 99636 584960 99876 4 analog_io[2]
port 23 nsew
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 24 nsew
rlabel metal3 s 583520 146556 584960 146796 4 analog_io[3]
port 25 nsew
rlabel metal3 s 583520 193476 584960 193716 4 analog_io[4]
port 26 nsew
rlabel metal3 s 583520 240396 584960 240636 4 analog_io[5]
port 27 nsew
rlabel metal3 s 583520 287316 584960 287556 4 analog_io[6]
port 28 nsew
rlabel metal3 s 583520 334236 584960 334476 4 analog_io[7]
port 29 nsew
rlabel metal3 s 583520 381156 584960 381396 4 analog_io[8]
port 30 nsew
rlabel metal3 s 583520 428076 584960 428316 4 analog_io[9]
port 31 nsew
rlabel metal3 s 583520 17492 584960 17732 4 io_in[0]
port 32 nsew
rlabel metal3 s 583520 486692 584960 486932 4 io_in[10]
port 33 nsew
rlabel metal3 s 583520 533748 584960 533988 4 io_in[11]
port 34 nsew
rlabel metal3 s 583520 580668 584960 580908 4 io_in[12]
port 35 nsew
rlabel metal3 s 583520 627588 584960 627828 4 io_in[13]
port 36 nsew
rlabel metal3 s 583520 674508 584960 674748 4 io_in[14]
port 37 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 38 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 39 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 40 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 41 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 42 nsew
rlabel metal3 s 583520 64412 584960 64652 4 io_in[1]
port 43 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 44 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 45 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 46 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 47 nsew
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 48 nsew
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 49 nsew
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 50 nsew
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 51 nsew
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 52 nsew
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 53 nsew
rlabel metal3 s 583520 111332 584960 111572 4 io_in[2]
port 54 nsew
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 55 nsew
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 56 nsew
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 57 nsew
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 58 nsew
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 59 nsew
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 60 nsew
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 61 nsew
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 62 nsew
rlabel metal3 s 583520 158252 584960 158492 4 io_in[3]
port 63 nsew
rlabel metal3 s 583520 205172 584960 205412 4 io_in[4]
port 64 nsew
rlabel metal3 s 583520 252092 584960 252332 4 io_in[5]
port 65 nsew
rlabel metal3 s 583520 299012 584960 299252 4 io_in[6]
port 66 nsew
rlabel metal3 s 583520 345932 584960 346172 4 io_in[7]
port 67 nsew
rlabel metal3 s 583520 392852 584960 393092 4 io_in[8]
port 68 nsew
rlabel metal3 s 583520 439772 584960 440012 4 io_in[9]
port 69 nsew
rlabel metal3 s 583520 40884 584960 41124 4 io_oeb[0]
port 70 nsew
rlabel metal3 s 583520 510220 584960 510460 4 io_oeb[10]
port 71 nsew
rlabel metal3 s 583520 557140 584960 557380 4 io_oeb[11]
port 72 nsew
rlabel metal3 s 583520 604060 584960 604300 4 io_oeb[12]
port 73 nsew
rlabel metal3 s 583520 650980 584960 651220 4 io_oeb[13]
port 74 nsew
rlabel metal3 s 583520 697900 584960 698140 4 io_oeb[14]
port 75 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 76 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 77 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 78 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 79 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 80 nsew
rlabel metal3 s 583520 87804 584960 88044 4 io_oeb[1]
port 81 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 82 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 83 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 84 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 85 nsew
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 86 nsew
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 87 nsew
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 88 nsew
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 89 nsew
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 90 nsew
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 91 nsew
rlabel metal3 s 583520 134724 584960 134964 4 io_oeb[2]
port 92 nsew
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 93 nsew
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 94 nsew
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 95 nsew
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 96 nsew
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 97 nsew
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 98 nsew
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 99 nsew
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 100 nsew
rlabel metal3 s 583520 181780 584960 182020 4 io_oeb[3]
port 101 nsew
rlabel metal3 s 583520 228700 584960 228940 4 io_oeb[4]
port 102 nsew
rlabel metal3 s 583520 275620 584960 275860 4 io_oeb[5]
port 103 nsew
rlabel metal3 s 583520 322540 584960 322780 4 io_oeb[6]
port 104 nsew
rlabel metal3 s 583520 369460 584960 369700 4 io_oeb[7]
port 105 nsew
rlabel metal3 s 583520 416380 584960 416620 4 io_oeb[8]
port 106 nsew
rlabel metal3 s 583520 463300 584960 463540 4 io_oeb[9]
port 107 nsew
rlabel metal3 s 583520 29188 584960 29428 4 io_out[0]
port 108 nsew
rlabel metal3 s 583520 498524 584960 498764 4 io_out[10]
port 109 nsew
rlabel metal3 s 583520 545444 584960 545684 4 io_out[11]
port 110 nsew
rlabel metal3 s 583520 592364 584960 592604 4 io_out[12]
port 111 nsew
rlabel metal3 s 583520 639284 584960 639524 4 io_out[13]
port 112 nsew
rlabel metal3 s 583520 686204 584960 686444 4 io_out[14]
port 113 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 114 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 115 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 116 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 117 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 118 nsew
rlabel metal3 s 583520 76108 584960 76348 4 io_out[1]
port 119 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 120 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 121 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 122 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 123 nsew
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 124 nsew
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 125 nsew
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 126 nsew
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 127 nsew
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 128 nsew
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 129 nsew
rlabel metal3 s 583520 123028 584960 123268 4 io_out[2]
port 130 nsew
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 131 nsew
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 132 nsew
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 133 nsew
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 134 nsew
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 135 nsew
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 136 nsew
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 137 nsew
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 138 nsew
rlabel metal3 s 583520 169948 584960 170188 4 io_out[3]
port 139 nsew
rlabel metal3 s 583520 216868 584960 217108 4 io_out[4]
port 140 nsew
rlabel metal3 s 583520 263788 584960 264028 4 io_out[5]
port 141 nsew
rlabel metal3 s 583520 310708 584960 310948 4 io_out[6]
port 142 nsew
rlabel metal3 s 583520 357764 584960 358004 4 io_out[7]
port 143 nsew
rlabel metal3 s 583520 404684 584960 404924 4 io_out[8]
port 144 nsew
rlabel metal3 s 583520 451604 584960 451844 4 io_out[9]
port 145 nsew
rlabel metal2 s 126582 -960 126694 480 4 la_data_in[0]
port 146 nsew
rlabel metal2 s 483450 -960 483562 480 4 la_data_in[100]
port 147 nsew
rlabel metal2 s 486946 -960 487058 480 4 la_data_in[101]
port 148 nsew
rlabel metal2 s 490534 -960 490646 480 4 la_data_in[102]
port 149 nsew
rlabel metal2 s 494122 -960 494234 480 4 la_data_in[103]
port 150 nsew
rlabel metal2 s 497710 -960 497822 480 4 la_data_in[104]
port 151 nsew
rlabel metal2 s 501206 -960 501318 480 4 la_data_in[105]
port 152 nsew
rlabel metal2 s 504794 -960 504906 480 4 la_data_in[106]
port 153 nsew
rlabel metal2 s 508382 -960 508494 480 4 la_data_in[107]
port 154 nsew
rlabel metal2 s 511970 -960 512082 480 4 la_data_in[108]
port 155 nsew
rlabel metal2 s 515558 -960 515670 480 4 la_data_in[109]
port 156 nsew
rlabel metal2 s 162278 -960 162390 480 4 la_data_in[10]
port 157 nsew
rlabel metal2 s 519054 -960 519166 480 4 la_data_in[110]
port 158 nsew
rlabel metal2 s 522642 -960 522754 480 4 la_data_in[111]
port 159 nsew
rlabel metal2 s 526230 -960 526342 480 4 la_data_in[112]
port 160 nsew
rlabel metal2 s 529818 -960 529930 480 4 la_data_in[113]
port 161 nsew
rlabel metal2 s 533406 -960 533518 480 4 la_data_in[114]
port 162 nsew
rlabel metal2 s 536902 -960 537014 480 4 la_data_in[115]
port 163 nsew
rlabel metal2 s 540490 -960 540602 480 4 la_data_in[116]
port 164 nsew
rlabel metal2 s 544078 -960 544190 480 4 la_data_in[117]
port 165 nsew
rlabel metal2 s 547666 -960 547778 480 4 la_data_in[118]
port 166 nsew
rlabel metal2 s 551162 -960 551274 480 4 la_data_in[119]
port 167 nsew
rlabel metal2 s 165866 -960 165978 480 4 la_data_in[11]
port 168 nsew
rlabel metal2 s 554750 -960 554862 480 4 la_data_in[120]
port 169 nsew
rlabel metal2 s 558338 -960 558450 480 4 la_data_in[121]
port 170 nsew
rlabel metal2 s 561926 -960 562038 480 4 la_data_in[122]
port 171 nsew
rlabel metal2 s 565514 -960 565626 480 4 la_data_in[123]
port 172 nsew
rlabel metal2 s 569010 -960 569122 480 4 la_data_in[124]
port 173 nsew
rlabel metal2 s 572598 -960 572710 480 4 la_data_in[125]
port 174 nsew
rlabel metal2 s 576186 -960 576298 480 4 la_data_in[126]
port 175 nsew
rlabel metal2 s 579774 -960 579886 480 4 la_data_in[127]
port 176 nsew
rlabel metal2 s 169362 -960 169474 480 4 la_data_in[12]
port 177 nsew
rlabel metal2 s 172950 -960 173062 480 4 la_data_in[13]
port 178 nsew
rlabel metal2 s 176538 -960 176650 480 4 la_data_in[14]
port 179 nsew
rlabel metal2 s 180126 -960 180238 480 4 la_data_in[15]
port 180 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_in[16]
port 181 nsew
rlabel metal2 s 187210 -960 187322 480 4 la_data_in[17]
port 182 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_in[18]
port 183 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_in[19]
port 184 nsew
rlabel metal2 s 130170 -960 130282 480 4 la_data_in[1]
port 185 nsew
rlabel metal2 s 197974 -960 198086 480 4 la_data_in[20]
port 186 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_in[21]
port 187 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_in[22]
port 188 nsew
rlabel metal2 s 208646 -960 208758 480 4 la_data_in[23]
port 189 nsew
rlabel metal2 s 212234 -960 212346 480 4 la_data_in[24]
port 190 nsew
rlabel metal2 s 215822 -960 215934 480 4 la_data_in[25]
port 191 nsew
rlabel metal2 s 219318 -960 219430 480 4 la_data_in[26]
port 192 nsew
rlabel metal2 s 222906 -960 223018 480 4 la_data_in[27]
port 193 nsew
rlabel metal2 s 226494 -960 226606 480 4 la_data_in[28]
port 194 nsew
rlabel metal2 s 230082 -960 230194 480 4 la_data_in[29]
port 195 nsew
rlabel metal2 s 133758 -960 133870 480 4 la_data_in[2]
port 196 nsew
rlabel metal2 s 233670 -960 233782 480 4 la_data_in[30]
port 197 nsew
rlabel metal2 s 237166 -960 237278 480 4 la_data_in[31]
port 198 nsew
rlabel metal2 s 240754 -960 240866 480 4 la_data_in[32]
port 199 nsew
rlabel metal2 s 244342 -960 244454 480 4 la_data_in[33]
port 200 nsew
rlabel metal2 s 247930 -960 248042 480 4 la_data_in[34]
port 201 nsew
rlabel metal2 s 251426 -960 251538 480 4 la_data_in[35]
port 202 nsew
rlabel metal2 s 255014 -960 255126 480 4 la_data_in[36]
port 203 nsew
rlabel metal2 s 258602 -960 258714 480 4 la_data_in[37]
port 204 nsew
rlabel metal2 s 262190 -960 262302 480 4 la_data_in[38]
port 205 nsew
rlabel metal2 s 265778 -960 265890 480 4 la_data_in[39]
port 206 nsew
rlabel metal2 s 137254 -960 137366 480 4 la_data_in[3]
port 207 nsew
rlabel metal2 s 269274 -960 269386 480 4 la_data_in[40]
port 208 nsew
rlabel metal2 s 272862 -960 272974 480 4 la_data_in[41]
port 209 nsew
rlabel metal2 s 276450 -960 276562 480 4 la_data_in[42]
port 210 nsew
rlabel metal2 s 280038 -960 280150 480 4 la_data_in[43]
port 211 nsew
rlabel metal2 s 283626 -960 283738 480 4 la_data_in[44]
port 212 nsew
rlabel metal2 s 287122 -960 287234 480 4 la_data_in[45]
port 213 nsew
rlabel metal2 s 290710 -960 290822 480 4 la_data_in[46]
port 214 nsew
rlabel metal2 s 294298 -960 294410 480 4 la_data_in[47]
port 215 nsew
rlabel metal2 s 297886 -960 297998 480 4 la_data_in[48]
port 216 nsew
rlabel metal2 s 301382 -960 301494 480 4 la_data_in[49]
port 217 nsew
rlabel metal2 s 140842 -960 140954 480 4 la_data_in[4]
port 218 nsew
rlabel metal2 s 304970 -960 305082 480 4 la_data_in[50]
port 219 nsew
rlabel metal2 s 308558 -960 308670 480 4 la_data_in[51]
port 220 nsew
rlabel metal2 s 312146 -960 312258 480 4 la_data_in[52]
port 221 nsew
rlabel metal2 s 315734 -960 315846 480 4 la_data_in[53]
port 222 nsew
rlabel metal2 s 319230 -960 319342 480 4 la_data_in[54]
port 223 nsew
rlabel metal2 s 322818 -960 322930 480 4 la_data_in[55]
port 224 nsew
rlabel metal2 s 326406 -960 326518 480 4 la_data_in[56]
port 225 nsew
rlabel metal2 s 329994 -960 330106 480 4 la_data_in[57]
port 226 nsew
rlabel metal2 s 333582 -960 333694 480 4 la_data_in[58]
port 227 nsew
rlabel metal2 s 337078 -960 337190 480 4 la_data_in[59]
port 228 nsew
rlabel metal2 s 144430 -960 144542 480 4 la_data_in[5]
port 229 nsew
rlabel metal2 s 340666 -960 340778 480 4 la_data_in[60]
port 230 nsew
rlabel metal2 s 344254 -960 344366 480 4 la_data_in[61]
port 231 nsew
rlabel metal2 s 347842 -960 347954 480 4 la_data_in[62]
port 232 nsew
rlabel metal2 s 351338 -960 351450 480 4 la_data_in[63]
port 233 nsew
rlabel metal2 s 354926 -960 355038 480 4 la_data_in[64]
port 234 nsew
rlabel metal2 s 358514 -960 358626 480 4 la_data_in[65]
port 235 nsew
rlabel metal2 s 362102 -960 362214 480 4 la_data_in[66]
port 236 nsew
rlabel metal2 s 365690 -960 365802 480 4 la_data_in[67]
port 237 nsew
rlabel metal2 s 369186 -960 369298 480 4 la_data_in[68]
port 238 nsew
rlabel metal2 s 372774 -960 372886 480 4 la_data_in[69]
port 239 nsew
rlabel metal2 s 148018 -960 148130 480 4 la_data_in[6]
port 240 nsew
rlabel metal2 s 376362 -960 376474 480 4 la_data_in[70]
port 241 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_data_in[71]
port 242 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_data_in[72]
port 243 nsew
rlabel metal2 s 387034 -960 387146 480 4 la_data_in[73]
port 244 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_data_in[74]
port 245 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_data_in[75]
port 246 nsew
rlabel metal2 s 397798 -960 397910 480 4 la_data_in[76]
port 247 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_data_in[77]
port 248 nsew
rlabel metal2 s 404882 -960 404994 480 4 la_data_in[78]
port 249 nsew
rlabel metal2 s 408470 -960 408582 480 4 la_data_in[79]
port 250 nsew
rlabel metal2 s 151514 -960 151626 480 4 la_data_in[7]
port 251 nsew
rlabel metal2 s 412058 -960 412170 480 4 la_data_in[80]
port 252 nsew
rlabel metal2 s 415646 -960 415758 480 4 la_data_in[81]
port 253 nsew
rlabel metal2 s 419142 -960 419254 480 4 la_data_in[82]
port 254 nsew
rlabel metal2 s 422730 -960 422842 480 4 la_data_in[83]
port 255 nsew
rlabel metal2 s 426318 -960 426430 480 4 la_data_in[84]
port 256 nsew
rlabel metal2 s 429906 -960 430018 480 4 la_data_in[85]
port 257 nsew
rlabel metal2 s 433494 -960 433606 480 4 la_data_in[86]
port 258 nsew
rlabel metal2 s 436990 -960 437102 480 4 la_data_in[87]
port 259 nsew
rlabel metal2 s 440578 -960 440690 480 4 la_data_in[88]
port 260 nsew
rlabel metal2 s 444166 -960 444278 480 4 la_data_in[89]
port 261 nsew
rlabel metal2 s 155102 -960 155214 480 4 la_data_in[8]
port 262 nsew
rlabel metal2 s 447754 -960 447866 480 4 la_data_in[90]
port 263 nsew
rlabel metal2 s 451250 -960 451362 480 4 la_data_in[91]
port 264 nsew
rlabel metal2 s 454838 -960 454950 480 4 la_data_in[92]
port 265 nsew
rlabel metal2 s 458426 -960 458538 480 4 la_data_in[93]
port 266 nsew
rlabel metal2 s 462014 -960 462126 480 4 la_data_in[94]
port 267 nsew
rlabel metal2 s 465602 -960 465714 480 4 la_data_in[95]
port 268 nsew
rlabel metal2 s 469098 -960 469210 480 4 la_data_in[96]
port 269 nsew
rlabel metal2 s 472686 -960 472798 480 4 la_data_in[97]
port 270 nsew
rlabel metal2 s 476274 -960 476386 480 4 la_data_in[98]
port 271 nsew
rlabel metal2 s 479862 -960 479974 480 4 la_data_in[99]
port 272 nsew
rlabel metal2 s 158690 -960 158802 480 4 la_data_in[9]
port 273 nsew
rlabel metal2 s 127778 -960 127890 480 4 la_data_out[0]
port 274 nsew
rlabel metal2 s 484554 -960 484666 480 4 la_data_out[100]
port 275 nsew
rlabel metal2 s 488142 -960 488254 480 4 la_data_out[101]
port 276 nsew
rlabel metal2 s 491730 -960 491842 480 4 la_data_out[102]
port 277 nsew
rlabel metal2 s 495318 -960 495430 480 4 la_data_out[103]
port 278 nsew
rlabel metal2 s 498906 -960 499018 480 4 la_data_out[104]
port 279 nsew
rlabel metal2 s 502402 -960 502514 480 4 la_data_out[105]
port 280 nsew
rlabel metal2 s 505990 -960 506102 480 4 la_data_out[106]
port 281 nsew
rlabel metal2 s 509578 -960 509690 480 4 la_data_out[107]
port 282 nsew
rlabel metal2 s 513166 -960 513278 480 4 la_data_out[108]
port 283 nsew
rlabel metal2 s 516754 -960 516866 480 4 la_data_out[109]
port 284 nsew
rlabel metal2 s 163474 -960 163586 480 4 la_data_out[10]
port 285 nsew
rlabel metal2 s 520250 -960 520362 480 4 la_data_out[110]
port 286 nsew
rlabel metal2 s 523838 -960 523950 480 4 la_data_out[111]
port 287 nsew
rlabel metal2 s 527426 -960 527538 480 4 la_data_out[112]
port 288 nsew
rlabel metal2 s 531014 -960 531126 480 4 la_data_out[113]
port 289 nsew
rlabel metal2 s 534510 -960 534622 480 4 la_data_out[114]
port 290 nsew
rlabel metal2 s 538098 -960 538210 480 4 la_data_out[115]
port 291 nsew
rlabel metal2 s 541686 -960 541798 480 4 la_data_out[116]
port 292 nsew
rlabel metal2 s 545274 -960 545386 480 4 la_data_out[117]
port 293 nsew
rlabel metal2 s 548862 -960 548974 480 4 la_data_out[118]
port 294 nsew
rlabel metal2 s 552358 -960 552470 480 4 la_data_out[119]
port 295 nsew
rlabel metal2 s 167062 -960 167174 480 4 la_data_out[11]
port 296 nsew
rlabel metal2 s 555946 -960 556058 480 4 la_data_out[120]
port 297 nsew
rlabel metal2 s 559534 -960 559646 480 4 la_data_out[121]
port 298 nsew
rlabel metal2 s 563122 -960 563234 480 4 la_data_out[122]
port 299 nsew
rlabel metal2 s 566710 -960 566822 480 4 la_data_out[123]
port 300 nsew
rlabel metal2 s 570206 -960 570318 480 4 la_data_out[124]
port 301 nsew
rlabel metal2 s 573794 -960 573906 480 4 la_data_out[125]
port 302 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[126]
port 303 nsew
rlabel metal2 s 580970 -960 581082 480 4 la_data_out[127]
port 304 nsew
rlabel metal2 s 170558 -960 170670 480 4 la_data_out[12]
port 305 nsew
rlabel metal2 s 174146 -960 174258 480 4 la_data_out[13]
port 306 nsew
rlabel metal2 s 177734 -960 177846 480 4 la_data_out[14]
port 307 nsew
rlabel metal2 s 181322 -960 181434 480 4 la_data_out[15]
port 308 nsew
rlabel metal2 s 184818 -960 184930 480 4 la_data_out[16]
port 309 nsew
rlabel metal2 s 188406 -960 188518 480 4 la_data_out[17]
port 310 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_data_out[18]
port 311 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_data_out[19]
port 312 nsew
rlabel metal2 s 131366 -960 131478 480 4 la_data_out[1]
port 313 nsew
rlabel metal2 s 199170 -960 199282 480 4 la_data_out[20]
port 314 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_data_out[21]
port 315 nsew
rlabel metal2 s 206254 -960 206366 480 4 la_data_out[22]
port 316 nsew
rlabel metal2 s 209842 -960 209954 480 4 la_data_out[23]
port 317 nsew
rlabel metal2 s 213430 -960 213542 480 4 la_data_out[24]
port 318 nsew
rlabel metal2 s 217018 -960 217130 480 4 la_data_out[25]
port 319 nsew
rlabel metal2 s 220514 -960 220626 480 4 la_data_out[26]
port 320 nsew
rlabel metal2 s 224102 -960 224214 480 4 la_data_out[27]
port 321 nsew
rlabel metal2 s 227690 -960 227802 480 4 la_data_out[28]
port 322 nsew
rlabel metal2 s 231278 -960 231390 480 4 la_data_out[29]
port 323 nsew
rlabel metal2 s 134862 -960 134974 480 4 la_data_out[2]
port 324 nsew
rlabel metal2 s 234774 -960 234886 480 4 la_data_out[30]
port 325 nsew
rlabel metal2 s 238362 -960 238474 480 4 la_data_out[31]
port 326 nsew
rlabel metal2 s 241950 -960 242062 480 4 la_data_out[32]
port 327 nsew
rlabel metal2 s 245538 -960 245650 480 4 la_data_out[33]
port 328 nsew
rlabel metal2 s 249126 -960 249238 480 4 la_data_out[34]
port 329 nsew
rlabel metal2 s 252622 -960 252734 480 4 la_data_out[35]
port 330 nsew
rlabel metal2 s 256210 -960 256322 480 4 la_data_out[36]
port 331 nsew
rlabel metal2 s 259798 -960 259910 480 4 la_data_out[37]
port 332 nsew
rlabel metal2 s 263386 -960 263498 480 4 la_data_out[38]
port 333 nsew
rlabel metal2 s 266974 -960 267086 480 4 la_data_out[39]
port 334 nsew
rlabel metal2 s 138450 -960 138562 480 4 la_data_out[3]
port 335 nsew
rlabel metal2 s 270470 -960 270582 480 4 la_data_out[40]
port 336 nsew
rlabel metal2 s 274058 -960 274170 480 4 la_data_out[41]
port 337 nsew
rlabel metal2 s 277646 -960 277758 480 4 la_data_out[42]
port 338 nsew
rlabel metal2 s 281234 -960 281346 480 4 la_data_out[43]
port 339 nsew
rlabel metal2 s 284730 -960 284842 480 4 la_data_out[44]
port 340 nsew
rlabel metal2 s 288318 -960 288430 480 4 la_data_out[45]
port 341 nsew
rlabel metal2 s 291906 -960 292018 480 4 la_data_out[46]
port 342 nsew
rlabel metal2 s 295494 -960 295606 480 4 la_data_out[47]
port 343 nsew
rlabel metal2 s 299082 -960 299194 480 4 la_data_out[48]
port 344 nsew
rlabel metal2 s 302578 -960 302690 480 4 la_data_out[49]
port 345 nsew
rlabel metal2 s 142038 -960 142150 480 4 la_data_out[4]
port 346 nsew
rlabel metal2 s 306166 -960 306278 480 4 la_data_out[50]
port 347 nsew
rlabel metal2 s 309754 -960 309866 480 4 la_data_out[51]
port 348 nsew
rlabel metal2 s 313342 -960 313454 480 4 la_data_out[52]
port 349 nsew
rlabel metal2 s 316930 -960 317042 480 4 la_data_out[53]
port 350 nsew
rlabel metal2 s 320426 -960 320538 480 4 la_data_out[54]
port 351 nsew
rlabel metal2 s 324014 -960 324126 480 4 la_data_out[55]
port 352 nsew
rlabel metal2 s 327602 -960 327714 480 4 la_data_out[56]
port 353 nsew
rlabel metal2 s 331190 -960 331302 480 4 la_data_out[57]
port 354 nsew
rlabel metal2 s 334686 -960 334798 480 4 la_data_out[58]
port 355 nsew
rlabel metal2 s 338274 -960 338386 480 4 la_data_out[59]
port 356 nsew
rlabel metal2 s 145626 -960 145738 480 4 la_data_out[5]
port 357 nsew
rlabel metal2 s 341862 -960 341974 480 4 la_data_out[60]
port 358 nsew
rlabel metal2 s 345450 -960 345562 480 4 la_data_out[61]
port 359 nsew
rlabel metal2 s 349038 -960 349150 480 4 la_data_out[62]
port 360 nsew
rlabel metal2 s 352534 -960 352646 480 4 la_data_out[63]
port 361 nsew
rlabel metal2 s 356122 -960 356234 480 4 la_data_out[64]
port 362 nsew
rlabel metal2 s 359710 -960 359822 480 4 la_data_out[65]
port 363 nsew
rlabel metal2 s 363298 -960 363410 480 4 la_data_out[66]
port 364 nsew
rlabel metal2 s 366886 -960 366998 480 4 la_data_out[67]
port 365 nsew
rlabel metal2 s 370382 -960 370494 480 4 la_data_out[68]
port 366 nsew
rlabel metal2 s 373970 -960 374082 480 4 la_data_out[69]
port 367 nsew
rlabel metal2 s 149214 -960 149326 480 4 la_data_out[6]
port 368 nsew
rlabel metal2 s 377558 -960 377670 480 4 la_data_out[70]
port 369 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_out[71]
port 370 nsew
rlabel metal2 s 384642 -960 384754 480 4 la_data_out[72]
port 371 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_out[73]
port 372 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_out[74]
port 373 nsew
rlabel metal2 s 395406 -960 395518 480 4 la_data_out[75]
port 374 nsew
rlabel metal2 s 398994 -960 399106 480 4 la_data_out[76]
port 375 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_out[77]
port 376 nsew
rlabel metal2 s 406078 -960 406190 480 4 la_data_out[78]
port 377 nsew
rlabel metal2 s 409666 -960 409778 480 4 la_data_out[79]
port 378 nsew
rlabel metal2 s 152710 -960 152822 480 4 la_data_out[7]
port 379 nsew
rlabel metal2 s 413254 -960 413366 480 4 la_data_out[80]
port 380 nsew
rlabel metal2 s 416842 -960 416954 480 4 la_data_out[81]
port 381 nsew
rlabel metal2 s 420338 -960 420450 480 4 la_data_out[82]
port 382 nsew
rlabel metal2 s 423926 -960 424038 480 4 la_data_out[83]
port 383 nsew
rlabel metal2 s 427514 -960 427626 480 4 la_data_out[84]
port 384 nsew
rlabel metal2 s 431102 -960 431214 480 4 la_data_out[85]
port 385 nsew
rlabel metal2 s 434598 -960 434710 480 4 la_data_out[86]
port 386 nsew
rlabel metal2 s 438186 -960 438298 480 4 la_data_out[87]
port 387 nsew
rlabel metal2 s 441774 -960 441886 480 4 la_data_out[88]
port 388 nsew
rlabel metal2 s 445362 -960 445474 480 4 la_data_out[89]
port 389 nsew
rlabel metal2 s 156298 -960 156410 480 4 la_data_out[8]
port 390 nsew
rlabel metal2 s 448950 -960 449062 480 4 la_data_out[90]
port 391 nsew
rlabel metal2 s 452446 -960 452558 480 4 la_data_out[91]
port 392 nsew
rlabel metal2 s 456034 -960 456146 480 4 la_data_out[92]
port 393 nsew
rlabel metal2 s 459622 -960 459734 480 4 la_data_out[93]
port 394 nsew
rlabel metal2 s 463210 -960 463322 480 4 la_data_out[94]
port 395 nsew
rlabel metal2 s 466798 -960 466910 480 4 la_data_out[95]
port 396 nsew
rlabel metal2 s 470294 -960 470406 480 4 la_data_out[96]
port 397 nsew
rlabel metal2 s 473882 -960 473994 480 4 la_data_out[97]
port 398 nsew
rlabel metal2 s 477470 -960 477582 480 4 la_data_out[98]
port 399 nsew
rlabel metal2 s 481058 -960 481170 480 4 la_data_out[99]
port 400 nsew
rlabel metal2 s 159886 -960 159998 480 4 la_data_out[9]
port 401 nsew
rlabel metal2 s 128974 -960 129086 480 4 la_oen[0]
port 402 nsew
rlabel metal2 s 485750 -960 485862 480 4 la_oen[100]
port 403 nsew
rlabel metal2 s 489338 -960 489450 480 4 la_oen[101]
port 404 nsew
rlabel metal2 s 492926 -960 493038 480 4 la_oen[102]
port 405 nsew
rlabel metal2 s 496514 -960 496626 480 4 la_oen[103]
port 406 nsew
rlabel metal2 s 500102 -960 500214 480 4 la_oen[104]
port 407 nsew
rlabel metal2 s 503598 -960 503710 480 4 la_oen[105]
port 408 nsew
rlabel metal2 s 507186 -960 507298 480 4 la_oen[106]
port 409 nsew
rlabel metal2 s 510774 -960 510886 480 4 la_oen[107]
port 410 nsew
rlabel metal2 s 514362 -960 514474 480 4 la_oen[108]
port 411 nsew
rlabel metal2 s 517858 -960 517970 480 4 la_oen[109]
port 412 nsew
rlabel metal2 s 164670 -960 164782 480 4 la_oen[10]
port 413 nsew
rlabel metal2 s 521446 -960 521558 480 4 la_oen[110]
port 414 nsew
rlabel metal2 s 525034 -960 525146 480 4 la_oen[111]
port 415 nsew
rlabel metal2 s 528622 -960 528734 480 4 la_oen[112]
port 416 nsew
rlabel metal2 s 532210 -960 532322 480 4 la_oen[113]
port 417 nsew
rlabel metal2 s 535706 -960 535818 480 4 la_oen[114]
port 418 nsew
rlabel metal2 s 539294 -960 539406 480 4 la_oen[115]
port 419 nsew
rlabel metal2 s 542882 -960 542994 480 4 la_oen[116]
port 420 nsew
rlabel metal2 s 546470 -960 546582 480 4 la_oen[117]
port 421 nsew
rlabel metal2 s 550058 -960 550170 480 4 la_oen[118]
port 422 nsew
rlabel metal2 s 553554 -960 553666 480 4 la_oen[119]
port 423 nsew
rlabel metal2 s 168166 -960 168278 480 4 la_oen[11]
port 424 nsew
rlabel metal2 s 557142 -960 557254 480 4 la_oen[120]
port 425 nsew
rlabel metal2 s 560730 -960 560842 480 4 la_oen[121]
port 426 nsew
rlabel metal2 s 564318 -960 564430 480 4 la_oen[122]
port 427 nsew
rlabel metal2 s 567814 -960 567926 480 4 la_oen[123]
port 428 nsew
rlabel metal2 s 571402 -960 571514 480 4 la_oen[124]
port 429 nsew
rlabel metal2 s 574990 -960 575102 480 4 la_oen[125]
port 430 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oen[126]
port 431 nsew
rlabel metal2 s 582166 -960 582278 480 4 la_oen[127]
port 432 nsew
rlabel metal2 s 171754 -960 171866 480 4 la_oen[12]
port 433 nsew
rlabel metal2 s 175342 -960 175454 480 4 la_oen[13]
port 434 nsew
rlabel metal2 s 178930 -960 179042 480 4 la_oen[14]
port 435 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_oen[15]
port 436 nsew
rlabel metal2 s 186014 -960 186126 480 4 la_oen[16]
port 437 nsew
rlabel metal2 s 189602 -960 189714 480 4 la_oen[17]
port 438 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_oen[18]
port 439 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_oen[19]
port 440 nsew
rlabel metal2 s 132562 -960 132674 480 4 la_oen[1]
port 441 nsew
rlabel metal2 s 200366 -960 200478 480 4 la_oen[20]
port 442 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_oen[21]
port 443 nsew
rlabel metal2 s 207450 -960 207562 480 4 la_oen[22]
port 444 nsew
rlabel metal2 s 211038 -960 211150 480 4 la_oen[23]
port 445 nsew
rlabel metal2 s 214626 -960 214738 480 4 la_oen[24]
port 446 nsew
rlabel metal2 s 218122 -960 218234 480 4 la_oen[25]
port 447 nsew
rlabel metal2 s 221710 -960 221822 480 4 la_oen[26]
port 448 nsew
rlabel metal2 s 225298 -960 225410 480 4 la_oen[27]
port 449 nsew
rlabel metal2 s 228886 -960 228998 480 4 la_oen[28]
port 450 nsew
rlabel metal2 s 232474 -960 232586 480 4 la_oen[29]
port 451 nsew
rlabel metal2 s 136058 -960 136170 480 4 la_oen[2]
port 452 nsew
rlabel metal2 s 235970 -960 236082 480 4 la_oen[30]
port 453 nsew
rlabel metal2 s 239558 -960 239670 480 4 la_oen[31]
port 454 nsew
rlabel metal2 s 243146 -960 243258 480 4 la_oen[32]
port 455 nsew
rlabel metal2 s 246734 -960 246846 480 4 la_oen[33]
port 456 nsew
rlabel metal2 s 250322 -960 250434 480 4 la_oen[34]
port 457 nsew
rlabel metal2 s 253818 -960 253930 480 4 la_oen[35]
port 458 nsew
rlabel metal2 s 257406 -960 257518 480 4 la_oen[36]
port 459 nsew
rlabel metal2 s 260994 -960 261106 480 4 la_oen[37]
port 460 nsew
rlabel metal2 s 264582 -960 264694 480 4 la_oen[38]
port 461 nsew
rlabel metal2 s 268078 -960 268190 480 4 la_oen[39]
port 462 nsew
rlabel metal2 s 139646 -960 139758 480 4 la_oen[3]
port 463 nsew
rlabel metal2 s 271666 -960 271778 480 4 la_oen[40]
port 464 nsew
rlabel metal2 s 275254 -960 275366 480 4 la_oen[41]
port 465 nsew
rlabel metal2 s 278842 -960 278954 480 4 la_oen[42]
port 466 nsew
rlabel metal2 s 282430 -960 282542 480 4 la_oen[43]
port 467 nsew
rlabel metal2 s 285926 -960 286038 480 4 la_oen[44]
port 468 nsew
rlabel metal2 s 289514 -960 289626 480 4 la_oen[45]
port 469 nsew
rlabel metal2 s 293102 -960 293214 480 4 la_oen[46]
port 470 nsew
rlabel metal2 s 296690 -960 296802 480 4 la_oen[47]
port 471 nsew
rlabel metal2 s 300278 -960 300390 480 4 la_oen[48]
port 472 nsew
rlabel metal2 s 303774 -960 303886 480 4 la_oen[49]
port 473 nsew
rlabel metal2 s 143234 -960 143346 480 4 la_oen[4]
port 474 nsew
rlabel metal2 s 307362 -960 307474 480 4 la_oen[50]
port 475 nsew
rlabel metal2 s 310950 -960 311062 480 4 la_oen[51]
port 476 nsew
rlabel metal2 s 314538 -960 314650 480 4 la_oen[52]
port 477 nsew
rlabel metal2 s 318034 -960 318146 480 4 la_oen[53]
port 478 nsew
rlabel metal2 s 321622 -960 321734 480 4 la_oen[54]
port 479 nsew
rlabel metal2 s 325210 -960 325322 480 4 la_oen[55]
port 480 nsew
rlabel metal2 s 328798 -960 328910 480 4 la_oen[56]
port 481 nsew
rlabel metal2 s 332386 -960 332498 480 4 la_oen[57]
port 482 nsew
rlabel metal2 s 335882 -960 335994 480 4 la_oen[58]
port 483 nsew
rlabel metal2 s 339470 -960 339582 480 4 la_oen[59]
port 484 nsew
rlabel metal2 s 146822 -960 146934 480 4 la_oen[5]
port 485 nsew
rlabel metal2 s 343058 -960 343170 480 4 la_oen[60]
port 486 nsew
rlabel metal2 s 346646 -960 346758 480 4 la_oen[61]
port 487 nsew
rlabel metal2 s 350234 -960 350346 480 4 la_oen[62]
port 488 nsew
rlabel metal2 s 353730 -960 353842 480 4 la_oen[63]
port 489 nsew
rlabel metal2 s 357318 -960 357430 480 4 la_oen[64]
port 490 nsew
rlabel metal2 s 360906 -960 361018 480 4 la_oen[65]
port 491 nsew
rlabel metal2 s 364494 -960 364606 480 4 la_oen[66]
port 492 nsew
rlabel metal2 s 367990 -960 368102 480 4 la_oen[67]
port 493 nsew
rlabel metal2 s 371578 -960 371690 480 4 la_oen[68]
port 494 nsew
rlabel metal2 s 375166 -960 375278 480 4 la_oen[69]
port 495 nsew
rlabel metal2 s 150410 -960 150522 480 4 la_oen[6]
port 496 nsew
rlabel metal2 s 378754 -960 378866 480 4 la_oen[70]
port 497 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_oen[71]
port 498 nsew
rlabel metal2 s 385838 -960 385950 480 4 la_oen[72]
port 499 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_oen[73]
port 500 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_oen[74]
port 501 nsew
rlabel metal2 s 396602 -960 396714 480 4 la_oen[75]
port 502 nsew
rlabel metal2 s 400190 -960 400302 480 4 la_oen[76]
port 503 nsew
rlabel metal2 s 403686 -960 403798 480 4 la_oen[77]
port 504 nsew
rlabel metal2 s 407274 -960 407386 480 4 la_oen[78]
port 505 nsew
rlabel metal2 s 410862 -960 410974 480 4 la_oen[79]
port 506 nsew
rlabel metal2 s 153906 -960 154018 480 4 la_oen[7]
port 507 nsew
rlabel metal2 s 414450 -960 414562 480 4 la_oen[80]
port 508 nsew
rlabel metal2 s 417946 -960 418058 480 4 la_oen[81]
port 509 nsew
rlabel metal2 s 421534 -960 421646 480 4 la_oen[82]
port 510 nsew
rlabel metal2 s 425122 -960 425234 480 4 la_oen[83]
port 511 nsew
rlabel metal2 s 428710 -960 428822 480 4 la_oen[84]
port 512 nsew
rlabel metal2 s 432298 -960 432410 480 4 la_oen[85]
port 513 nsew
rlabel metal2 s 435794 -960 435906 480 4 la_oen[86]
port 514 nsew
rlabel metal2 s 439382 -960 439494 480 4 la_oen[87]
port 515 nsew
rlabel metal2 s 442970 -960 443082 480 4 la_oen[88]
port 516 nsew
rlabel metal2 s 446558 -960 446670 480 4 la_oen[89]
port 517 nsew
rlabel metal2 s 157494 -960 157606 480 4 la_oen[8]
port 518 nsew
rlabel metal2 s 450146 -960 450258 480 4 la_oen[90]
port 519 nsew
rlabel metal2 s 453642 -960 453754 480 4 la_oen[91]
port 520 nsew
rlabel metal2 s 457230 -960 457342 480 4 la_oen[92]
port 521 nsew
rlabel metal2 s 460818 -960 460930 480 4 la_oen[93]
port 522 nsew
rlabel metal2 s 464406 -960 464518 480 4 la_oen[94]
port 523 nsew
rlabel metal2 s 467902 -960 468014 480 4 la_oen[95]
port 524 nsew
rlabel metal2 s 471490 -960 471602 480 4 la_oen[96]
port 525 nsew
rlabel metal2 s 475078 -960 475190 480 4 la_oen[97]
port 526 nsew
rlabel metal2 s 478666 -960 478778 480 4 la_oen[98]
port 527 nsew
rlabel metal2 s 482254 -960 482366 480 4 la_oen[99]
port 528 nsew
rlabel metal2 s 161082 -960 161194 480 4 la_oen[9]
port 529 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_clock2
port 530 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 531 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 532 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 533 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 534 nsew
rlabel metal2 s 48106 -960 48218 480 4 wbs_adr_i[10]
port 535 nsew
rlabel metal2 s 51602 -960 51714 480 4 wbs_adr_i[11]
port 536 nsew
rlabel metal2 s 55190 -960 55302 480 4 wbs_adr_i[12]
port 537 nsew
rlabel metal2 s 58778 -960 58890 480 4 wbs_adr_i[13]
port 538 nsew
rlabel metal2 s 62366 -960 62478 480 4 wbs_adr_i[14]
port 539 nsew
rlabel metal2 s 65954 -960 66066 480 4 wbs_adr_i[15]
port 540 nsew
rlabel metal2 s 69450 -960 69562 480 4 wbs_adr_i[16]
port 541 nsew
rlabel metal2 s 73038 -960 73150 480 4 wbs_adr_i[17]
port 542 nsew
rlabel metal2 s 76626 -960 76738 480 4 wbs_adr_i[18]
port 543 nsew
rlabel metal2 s 80214 -960 80326 480 4 wbs_adr_i[19]
port 544 nsew
rlabel metal2 s 12410 -960 12522 480 4 wbs_adr_i[1]
port 545 nsew
rlabel metal2 s 83802 -960 83914 480 4 wbs_adr_i[20]
port 546 nsew
rlabel metal2 s 87298 -960 87410 480 4 wbs_adr_i[21]
port 547 nsew
rlabel metal2 s 90886 -960 90998 480 4 wbs_adr_i[22]
port 548 nsew
rlabel metal2 s 94474 -960 94586 480 4 wbs_adr_i[23]
port 549 nsew
rlabel metal2 s 98062 -960 98174 480 4 wbs_adr_i[24]
port 550 nsew
rlabel metal2 s 101558 -960 101670 480 4 wbs_adr_i[25]
port 551 nsew
rlabel metal2 s 105146 -960 105258 480 4 wbs_adr_i[26]
port 552 nsew
rlabel metal2 s 108734 -960 108846 480 4 wbs_adr_i[27]
port 553 nsew
rlabel metal2 s 112322 -960 112434 480 4 wbs_adr_i[28]
port 554 nsew
rlabel metal2 s 115910 -960 116022 480 4 wbs_adr_i[29]
port 555 nsew
rlabel metal2 s 17194 -960 17306 480 4 wbs_adr_i[2]
port 556 nsew
rlabel metal2 s 119406 -960 119518 480 4 wbs_adr_i[30]
port 557 nsew
rlabel metal2 s 122994 -960 123106 480 4 wbs_adr_i[31]
port 558 nsew
rlabel metal2 s 21886 -960 21998 480 4 wbs_adr_i[3]
port 559 nsew
rlabel metal2 s 26670 -960 26782 480 4 wbs_adr_i[4]
port 560 nsew
rlabel metal2 s 30258 -960 30370 480 4 wbs_adr_i[5]
port 561 nsew
rlabel metal2 s 33846 -960 33958 480 4 wbs_adr_i[6]
port 562 nsew
rlabel metal2 s 37342 -960 37454 480 4 wbs_adr_i[7]
port 563 nsew
rlabel metal2 s 40930 -960 41042 480 4 wbs_adr_i[8]
port 564 nsew
rlabel metal2 s 44518 -960 44630 480 4 wbs_adr_i[9]
port 565 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 566 nsew
rlabel metal2 s 8822 -960 8934 480 4 wbs_dat_i[0]
port 567 nsew
rlabel metal2 s 49302 -960 49414 480 4 wbs_dat_i[10]
port 568 nsew
rlabel metal2 s 52798 -960 52910 480 4 wbs_dat_i[11]
port 569 nsew
rlabel metal2 s 56386 -960 56498 480 4 wbs_dat_i[12]
port 570 nsew
rlabel metal2 s 59974 -960 60086 480 4 wbs_dat_i[13]
port 571 nsew
rlabel metal2 s 63562 -960 63674 480 4 wbs_dat_i[14]
port 572 nsew
rlabel metal2 s 67150 -960 67262 480 4 wbs_dat_i[15]
port 573 nsew
rlabel metal2 s 70646 -960 70758 480 4 wbs_dat_i[16]
port 574 nsew
rlabel metal2 s 74234 -960 74346 480 4 wbs_dat_i[17]
port 575 nsew
rlabel metal2 s 77822 -960 77934 480 4 wbs_dat_i[18]
port 576 nsew
rlabel metal2 s 81410 -960 81522 480 4 wbs_dat_i[19]
port 577 nsew
rlabel metal2 s 13606 -960 13718 480 4 wbs_dat_i[1]
port 578 nsew
rlabel metal2 s 84906 -960 85018 480 4 wbs_dat_i[20]
port 579 nsew
rlabel metal2 s 88494 -960 88606 480 4 wbs_dat_i[21]
port 580 nsew
rlabel metal2 s 92082 -960 92194 480 4 wbs_dat_i[22]
port 581 nsew
rlabel metal2 s 95670 -960 95782 480 4 wbs_dat_i[23]
port 582 nsew
rlabel metal2 s 99258 -960 99370 480 4 wbs_dat_i[24]
port 583 nsew
rlabel metal2 s 102754 -960 102866 480 4 wbs_dat_i[25]
port 584 nsew
rlabel metal2 s 106342 -960 106454 480 4 wbs_dat_i[26]
port 585 nsew
rlabel metal2 s 109930 -960 110042 480 4 wbs_dat_i[27]
port 586 nsew
rlabel metal2 s 113518 -960 113630 480 4 wbs_dat_i[28]
port 587 nsew
rlabel metal2 s 117106 -960 117218 480 4 wbs_dat_i[29]
port 588 nsew
rlabel metal2 s 18298 -960 18410 480 4 wbs_dat_i[2]
port 589 nsew
rlabel metal2 s 120602 -960 120714 480 4 wbs_dat_i[30]
port 590 nsew
rlabel metal2 s 124190 -960 124302 480 4 wbs_dat_i[31]
port 591 nsew
rlabel metal2 s 23082 -960 23194 480 4 wbs_dat_i[3]
port 592 nsew
rlabel metal2 s 27866 -960 27978 480 4 wbs_dat_i[4]
port 593 nsew
rlabel metal2 s 31454 -960 31566 480 4 wbs_dat_i[5]
port 594 nsew
rlabel metal2 s 34950 -960 35062 480 4 wbs_dat_i[6]
port 595 nsew
rlabel metal2 s 38538 -960 38650 480 4 wbs_dat_i[7]
port 596 nsew
rlabel metal2 s 42126 -960 42238 480 4 wbs_dat_i[8]
port 597 nsew
rlabel metal2 s 45714 -960 45826 480 4 wbs_dat_i[9]
port 598 nsew
rlabel metal2 s 10018 -960 10130 480 4 wbs_dat_o[0]
port 599 nsew
rlabel metal2 s 50498 -960 50610 480 4 wbs_dat_o[10]
port 600 nsew
rlabel metal2 s 53994 -960 54106 480 4 wbs_dat_o[11]
port 601 nsew
rlabel metal2 s 57582 -960 57694 480 4 wbs_dat_o[12]
port 602 nsew
rlabel metal2 s 61170 -960 61282 480 4 wbs_dat_o[13]
port 603 nsew
rlabel metal2 s 64758 -960 64870 480 4 wbs_dat_o[14]
port 604 nsew
rlabel metal2 s 68254 -960 68366 480 4 wbs_dat_o[15]
port 605 nsew
rlabel metal2 s 71842 -960 71954 480 4 wbs_dat_o[16]
port 606 nsew
rlabel metal2 s 75430 -960 75542 480 4 wbs_dat_o[17]
port 607 nsew
rlabel metal2 s 79018 -960 79130 480 4 wbs_dat_o[18]
port 608 nsew
rlabel metal2 s 82606 -960 82718 480 4 wbs_dat_o[19]
port 609 nsew
rlabel metal2 s 14802 -960 14914 480 4 wbs_dat_o[1]
port 610 nsew
rlabel metal2 s 86102 -960 86214 480 4 wbs_dat_o[20]
port 611 nsew
rlabel metal2 s 89690 -960 89802 480 4 wbs_dat_o[21]
port 612 nsew
rlabel metal2 s 93278 -960 93390 480 4 wbs_dat_o[22]
port 613 nsew
rlabel metal2 s 96866 -960 96978 480 4 wbs_dat_o[23]
port 614 nsew
rlabel metal2 s 100454 -960 100566 480 4 wbs_dat_o[24]
port 615 nsew
rlabel metal2 s 103950 -960 104062 480 4 wbs_dat_o[25]
port 616 nsew
rlabel metal2 s 107538 -960 107650 480 4 wbs_dat_o[26]
port 617 nsew
rlabel metal2 s 111126 -960 111238 480 4 wbs_dat_o[27]
port 618 nsew
rlabel metal2 s 114714 -960 114826 480 4 wbs_dat_o[28]
port 619 nsew
rlabel metal2 s 118210 -960 118322 480 4 wbs_dat_o[29]
port 620 nsew
rlabel metal2 s 19494 -960 19606 480 4 wbs_dat_o[2]
port 621 nsew
rlabel metal2 s 121798 -960 121910 480 4 wbs_dat_o[30]
port 622 nsew
rlabel metal2 s 125386 -960 125498 480 4 wbs_dat_o[31]
port 623 nsew
rlabel metal2 s 24278 -960 24390 480 4 wbs_dat_o[3]
port 624 nsew
rlabel metal2 s 29062 -960 29174 480 4 wbs_dat_o[4]
port 625 nsew
rlabel metal2 s 32650 -960 32762 480 4 wbs_dat_o[5]
port 626 nsew
rlabel metal2 s 36146 -960 36258 480 4 wbs_dat_o[6]
port 627 nsew
rlabel metal2 s 39734 -960 39846 480 4 wbs_dat_o[7]
port 628 nsew
rlabel metal2 s 43322 -960 43434 480 4 wbs_dat_o[8]
port 629 nsew
rlabel metal2 s 46910 -960 47022 480 4 wbs_dat_o[9]
port 630 nsew
rlabel metal2 s 11214 -960 11326 480 4 wbs_sel_i[0]
port 631 nsew
rlabel metal2 s 15998 -960 16110 480 4 wbs_sel_i[1]
port 632 nsew
rlabel metal2 s 20690 -960 20802 480 4 wbs_sel_i[2]
port 633 nsew
rlabel metal2 s 25474 -960 25586 480 4 wbs_sel_i[3]
port 634 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 635 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 636 nsew
rlabel metal5 s -1996 -924 585920 -324 4 vccd1
port 637 nsew
rlabel metal5 s -2916 -1844 586840 -1244 4 vssd1
port 638 nsew
rlabel metal5 s -3836 -2764 587760 -2164 4 vccd2
port 639 nsew
rlabel metal5 s -4756 -3684 588680 -3084 4 vssd2
port 640 nsew
rlabel metal5 s -5676 -4604 589600 -4004 4 vdda1
port 641 nsew
rlabel metal5 s -6596 -5524 590520 -4924 4 vssa1
port 642 nsew
rlabel metal5 s -7516 -6444 591440 -5844 4 vdda2
port 643 nsew
rlabel metal5 s -8436 -7364 592360 -6764 4 vssa2
port 644 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 221762806
string GDS_START 218527394
<< end >>
