magic
tech sky130A
magscale 1 2
timestamp 1607587669
<< obsli1 >>
rect 1104 2159 418876 497777
<< obsm1 >>
rect 474 892 418876 497808
<< metal2 >>
rect 7746 499200 7802 500000
rect 23294 499200 23350 500000
rect 38842 499200 38898 500000
rect 54390 499200 54446 500000
rect 69938 499200 69994 500000
rect 85486 499200 85542 500000
rect 101034 499200 101090 500000
rect 116582 499200 116638 500000
rect 132130 499200 132186 500000
rect 147678 499200 147734 500000
rect 163226 499200 163282 500000
rect 178774 499200 178830 500000
rect 194322 499200 194378 500000
rect 209870 499200 209926 500000
rect 225510 499200 225566 500000
rect 241058 499200 241114 500000
rect 256606 499200 256662 500000
rect 272154 499200 272210 500000
rect 287702 499200 287758 500000
rect 303250 499200 303306 500000
rect 318798 499200 318854 500000
rect 334346 499200 334402 500000
rect 349894 499200 349950 500000
rect 365442 499200 365498 500000
rect 380990 499200 381046 500000
rect 396538 499200 396594 500000
rect 412086 499200 412142 500000
rect 478 0 534 800
rect 1490 0 1546 800
rect 2594 0 2650 800
rect 3698 0 3754 800
rect 4802 0 4858 800
rect 5906 0 5962 800
rect 6918 0 6974 800
rect 8022 0 8078 800
rect 9126 0 9182 800
rect 10230 0 10286 800
rect 11334 0 11390 800
rect 12438 0 12494 800
rect 13450 0 13506 800
rect 14554 0 14610 800
rect 15658 0 15714 800
rect 16762 0 16818 800
rect 17866 0 17922 800
rect 18970 0 19026 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26514 0 26570 800
rect 27618 0 27674 800
rect 28722 0 28778 800
rect 29826 0 29882 800
rect 30930 0 30986 800
rect 31942 0 31998 800
rect 33046 0 33102 800
rect 34150 0 34206 800
rect 35254 0 35310 800
rect 36358 0 36414 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39578 0 39634 800
rect 40682 0 40738 800
rect 41786 0 41842 800
rect 42890 0 42946 800
rect 43994 0 44050 800
rect 45006 0 45062 800
rect 46110 0 46166 800
rect 47214 0 47270 800
rect 48318 0 48374 800
rect 49422 0 49478 800
rect 50526 0 50582 800
rect 51538 0 51594 800
rect 52642 0 52698 800
rect 53746 0 53802 800
rect 54850 0 54906 800
rect 55954 0 56010 800
rect 56966 0 57022 800
rect 58070 0 58126 800
rect 59174 0 59230 800
rect 60278 0 60334 800
rect 61382 0 61438 800
rect 62486 0 62542 800
rect 63498 0 63554 800
rect 64602 0 64658 800
rect 65706 0 65762 800
rect 66810 0 66866 800
rect 67914 0 67970 800
rect 69018 0 69074 800
rect 70030 0 70086 800
rect 71134 0 71190 800
rect 72238 0 72294 800
rect 73342 0 73398 800
rect 74446 0 74502 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77666 0 77722 800
rect 78770 0 78826 800
rect 79874 0 79930 800
rect 80978 0 81034 800
rect 81990 0 82046 800
rect 83094 0 83150 800
rect 84198 0 84254 800
rect 85302 0 85358 800
rect 86406 0 86462 800
rect 87510 0 87566 800
rect 88522 0 88578 800
rect 89626 0 89682 800
rect 90730 0 90786 800
rect 91834 0 91890 800
rect 92938 0 92994 800
rect 94042 0 94098 800
rect 95054 0 95110 800
rect 96158 0 96214 800
rect 97262 0 97318 800
rect 98366 0 98422 800
rect 99470 0 99526 800
rect 100574 0 100630 800
rect 101586 0 101642 800
rect 102690 0 102746 800
rect 103794 0 103850 800
rect 104898 0 104954 800
rect 106002 0 106058 800
rect 107014 0 107070 800
rect 108118 0 108174 800
rect 109222 0 109278 800
rect 110326 0 110382 800
rect 111430 0 111486 800
rect 112534 0 112590 800
rect 113546 0 113602 800
rect 114650 0 114706 800
rect 115754 0 115810 800
rect 116858 0 116914 800
rect 117962 0 118018 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121182 0 121238 800
rect 122286 0 122342 800
rect 123390 0 123446 800
rect 124494 0 124550 800
rect 125598 0 125654 800
rect 126610 0 126666 800
rect 127714 0 127770 800
rect 128818 0 128874 800
rect 129922 0 129978 800
rect 131026 0 131082 800
rect 132038 0 132094 800
rect 133142 0 133198 800
rect 134246 0 134302 800
rect 135350 0 135406 800
rect 136454 0 136510 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139674 0 139730 800
rect 140778 0 140834 800
rect 141882 0 141938 800
rect 142986 0 143042 800
rect 144090 0 144146 800
rect 145102 0 145158 800
rect 146206 0 146262 800
rect 147310 0 147366 800
rect 148414 0 148470 800
rect 149518 0 149574 800
rect 150622 0 150678 800
rect 151634 0 151690 800
rect 152738 0 152794 800
rect 153842 0 153898 800
rect 154946 0 155002 800
rect 156050 0 156106 800
rect 157154 0 157210 800
rect 158166 0 158222 800
rect 159270 0 159326 800
rect 160374 0 160430 800
rect 161478 0 161534 800
rect 162582 0 162638 800
rect 163594 0 163650 800
rect 164698 0 164754 800
rect 165802 0 165858 800
rect 166906 0 166962 800
rect 168010 0 168066 800
rect 169114 0 169170 800
rect 170126 0 170182 800
rect 171230 0 171286 800
rect 172334 0 172390 800
rect 173438 0 173494 800
rect 174542 0 174598 800
rect 175646 0 175702 800
rect 176658 0 176714 800
rect 177762 0 177818 800
rect 178866 0 178922 800
rect 179970 0 180026 800
rect 181074 0 181130 800
rect 182178 0 182234 800
rect 183190 0 183246 800
rect 184294 0 184350 800
rect 185398 0 185454 800
rect 186502 0 186558 800
rect 187606 0 187662 800
rect 188618 0 188674 800
rect 189722 0 189778 800
rect 190826 0 190882 800
rect 191930 0 191986 800
rect 193034 0 193090 800
rect 194138 0 194194 800
rect 195150 0 195206 800
rect 196254 0 196310 800
rect 197358 0 197414 800
rect 198462 0 198518 800
rect 199566 0 199622 800
rect 200670 0 200726 800
rect 201682 0 201738 800
rect 202786 0 202842 800
rect 203890 0 203946 800
rect 204994 0 205050 800
rect 206098 0 206154 800
rect 207202 0 207258 800
rect 208214 0 208270 800
rect 209318 0 209374 800
rect 210422 0 210478 800
rect 211526 0 211582 800
rect 212630 0 212686 800
rect 213642 0 213698 800
rect 214746 0 214802 800
rect 215850 0 215906 800
rect 216954 0 217010 800
rect 218058 0 218114 800
rect 219162 0 219218 800
rect 220174 0 220230 800
rect 221278 0 221334 800
rect 222382 0 222438 800
rect 223486 0 223542 800
rect 224590 0 224646 800
rect 225694 0 225750 800
rect 226706 0 226762 800
rect 227810 0 227866 800
rect 228914 0 228970 800
rect 230018 0 230074 800
rect 231122 0 231178 800
rect 232226 0 232282 800
rect 233238 0 233294 800
rect 234342 0 234398 800
rect 235446 0 235502 800
rect 236550 0 236606 800
rect 237654 0 237710 800
rect 238666 0 238722 800
rect 239770 0 239826 800
rect 240874 0 240930 800
rect 241978 0 242034 800
rect 243082 0 243138 800
rect 244186 0 244242 800
rect 245198 0 245254 800
rect 246302 0 246358 800
rect 247406 0 247462 800
rect 248510 0 248566 800
rect 249614 0 249670 800
rect 250718 0 250774 800
rect 251730 0 251786 800
rect 252834 0 252890 800
rect 253938 0 253994 800
rect 255042 0 255098 800
rect 256146 0 256202 800
rect 257250 0 257306 800
rect 258262 0 258318 800
rect 259366 0 259422 800
rect 260470 0 260526 800
rect 261574 0 261630 800
rect 262678 0 262734 800
rect 263690 0 263746 800
rect 264794 0 264850 800
rect 265898 0 265954 800
rect 267002 0 267058 800
rect 268106 0 268162 800
rect 269210 0 269266 800
rect 270222 0 270278 800
rect 271326 0 271382 800
rect 272430 0 272486 800
rect 273534 0 273590 800
rect 274638 0 274694 800
rect 275742 0 275798 800
rect 276754 0 276810 800
rect 277858 0 277914 800
rect 278962 0 279018 800
rect 280066 0 280122 800
rect 281170 0 281226 800
rect 282274 0 282330 800
rect 283286 0 283342 800
rect 284390 0 284446 800
rect 285494 0 285550 800
rect 286598 0 286654 800
rect 287702 0 287758 800
rect 288806 0 288862 800
rect 289818 0 289874 800
rect 290922 0 290978 800
rect 292026 0 292082 800
rect 293130 0 293186 800
rect 294234 0 294290 800
rect 295246 0 295302 800
rect 296350 0 296406 800
rect 297454 0 297510 800
rect 298558 0 298614 800
rect 299662 0 299718 800
rect 300766 0 300822 800
rect 301778 0 301834 800
rect 302882 0 302938 800
rect 303986 0 304042 800
rect 305090 0 305146 800
rect 306194 0 306250 800
rect 307298 0 307354 800
rect 308310 0 308366 800
rect 309414 0 309470 800
rect 310518 0 310574 800
rect 311622 0 311678 800
rect 312726 0 312782 800
rect 313830 0 313886 800
rect 314842 0 314898 800
rect 315946 0 316002 800
rect 317050 0 317106 800
rect 318154 0 318210 800
rect 319258 0 319314 800
rect 320270 0 320326 800
rect 321374 0 321430 800
rect 322478 0 322534 800
rect 323582 0 323638 800
rect 324686 0 324742 800
rect 325790 0 325846 800
rect 326802 0 326858 800
rect 327906 0 327962 800
rect 329010 0 329066 800
rect 330114 0 330170 800
rect 331218 0 331274 800
rect 332322 0 332378 800
rect 333334 0 333390 800
rect 334438 0 334494 800
rect 335542 0 335598 800
rect 336646 0 336702 800
rect 337750 0 337806 800
rect 338854 0 338910 800
rect 339866 0 339922 800
rect 340970 0 341026 800
rect 342074 0 342130 800
rect 343178 0 343234 800
rect 344282 0 344338 800
rect 345294 0 345350 800
rect 346398 0 346454 800
rect 347502 0 347558 800
rect 348606 0 348662 800
rect 349710 0 349766 800
rect 350814 0 350870 800
rect 351826 0 351882 800
rect 352930 0 352986 800
rect 354034 0 354090 800
rect 355138 0 355194 800
rect 356242 0 356298 800
rect 357346 0 357402 800
rect 358358 0 358414 800
rect 359462 0 359518 800
rect 360566 0 360622 800
rect 361670 0 361726 800
rect 362774 0 362830 800
rect 363878 0 363934 800
rect 364890 0 364946 800
rect 365994 0 366050 800
rect 367098 0 367154 800
rect 368202 0 368258 800
rect 369306 0 369362 800
rect 370318 0 370374 800
rect 371422 0 371478 800
rect 372526 0 372582 800
rect 373630 0 373686 800
rect 374734 0 374790 800
rect 375838 0 375894 800
rect 376850 0 376906 800
rect 377954 0 378010 800
rect 379058 0 379114 800
rect 380162 0 380218 800
rect 381266 0 381322 800
rect 382370 0 382426 800
rect 383382 0 383438 800
rect 384486 0 384542 800
rect 385590 0 385646 800
rect 386694 0 386750 800
rect 387798 0 387854 800
rect 388902 0 388958 800
rect 389914 0 389970 800
rect 391018 0 391074 800
rect 392122 0 392178 800
rect 393226 0 393282 800
rect 394330 0 394386 800
rect 395342 0 395398 800
rect 396446 0 396502 800
rect 397550 0 397606 800
rect 398654 0 398710 800
rect 399758 0 399814 800
rect 400862 0 400918 800
rect 401874 0 401930 800
rect 402978 0 403034 800
rect 404082 0 404138 800
rect 405186 0 405242 800
rect 406290 0 406346 800
rect 407394 0 407450 800
rect 408406 0 408462 800
rect 409510 0 409566 800
rect 410614 0 410670 800
rect 411718 0 411774 800
rect 412822 0 412878 800
rect 413926 0 413982 800
rect 414938 0 414994 800
rect 416042 0 416098 800
rect 417146 0 417202 800
rect 418250 0 418306 800
rect 419354 0 419410 800
<< obsm2 >>
rect 480 499144 7690 499202
rect 7858 499144 23238 499202
rect 23406 499144 38786 499202
rect 38954 499144 54334 499202
rect 54502 499144 69882 499202
rect 70050 499144 85430 499202
rect 85598 499144 100978 499202
rect 101146 499144 116526 499202
rect 116694 499144 132074 499202
rect 132242 499144 147622 499202
rect 147790 499144 163170 499202
rect 163338 499144 178718 499202
rect 178886 499144 194266 499202
rect 194434 499144 209814 499202
rect 209982 499144 225454 499202
rect 225622 499144 241002 499202
rect 241170 499144 256550 499202
rect 256718 499144 272098 499202
rect 272266 499144 287646 499202
rect 287814 499144 303194 499202
rect 303362 499144 318742 499202
rect 318910 499144 334290 499202
rect 334458 499144 349838 499202
rect 350006 499144 365386 499202
rect 365554 499144 380934 499202
rect 381102 499144 396482 499202
rect 396650 499144 412030 499202
rect 412198 499144 418304 499202
rect 480 856 418304 499144
rect 590 800 1434 856
rect 1602 800 2538 856
rect 2706 800 3642 856
rect 3810 800 4746 856
rect 4914 800 5850 856
rect 6018 800 6862 856
rect 7030 800 7966 856
rect 8134 800 9070 856
rect 9238 800 10174 856
rect 10342 800 11278 856
rect 11446 800 12382 856
rect 12550 800 13394 856
rect 13562 800 14498 856
rect 14666 800 15602 856
rect 15770 800 16706 856
rect 16874 800 17810 856
rect 17978 800 18914 856
rect 19082 800 19926 856
rect 20094 800 21030 856
rect 21198 800 22134 856
rect 22302 800 23238 856
rect 23406 800 24342 856
rect 24510 800 25446 856
rect 25614 800 26458 856
rect 26626 800 27562 856
rect 27730 800 28666 856
rect 28834 800 29770 856
rect 29938 800 30874 856
rect 31042 800 31886 856
rect 32054 800 32990 856
rect 33158 800 34094 856
rect 34262 800 35198 856
rect 35366 800 36302 856
rect 36470 800 37406 856
rect 37574 800 38418 856
rect 38586 800 39522 856
rect 39690 800 40626 856
rect 40794 800 41730 856
rect 41898 800 42834 856
rect 43002 800 43938 856
rect 44106 800 44950 856
rect 45118 800 46054 856
rect 46222 800 47158 856
rect 47326 800 48262 856
rect 48430 800 49366 856
rect 49534 800 50470 856
rect 50638 800 51482 856
rect 51650 800 52586 856
rect 52754 800 53690 856
rect 53858 800 54794 856
rect 54962 800 55898 856
rect 56066 800 56910 856
rect 57078 800 58014 856
rect 58182 800 59118 856
rect 59286 800 60222 856
rect 60390 800 61326 856
rect 61494 800 62430 856
rect 62598 800 63442 856
rect 63610 800 64546 856
rect 64714 800 65650 856
rect 65818 800 66754 856
rect 66922 800 67858 856
rect 68026 800 68962 856
rect 69130 800 69974 856
rect 70142 800 71078 856
rect 71246 800 72182 856
rect 72350 800 73286 856
rect 73454 800 74390 856
rect 74558 800 75494 856
rect 75662 800 76506 856
rect 76674 800 77610 856
rect 77778 800 78714 856
rect 78882 800 79818 856
rect 79986 800 80922 856
rect 81090 800 81934 856
rect 82102 800 83038 856
rect 83206 800 84142 856
rect 84310 800 85246 856
rect 85414 800 86350 856
rect 86518 800 87454 856
rect 87622 800 88466 856
rect 88634 800 89570 856
rect 89738 800 90674 856
rect 90842 800 91778 856
rect 91946 800 92882 856
rect 93050 800 93986 856
rect 94154 800 94998 856
rect 95166 800 96102 856
rect 96270 800 97206 856
rect 97374 800 98310 856
rect 98478 800 99414 856
rect 99582 800 100518 856
rect 100686 800 101530 856
rect 101698 800 102634 856
rect 102802 800 103738 856
rect 103906 800 104842 856
rect 105010 800 105946 856
rect 106114 800 106958 856
rect 107126 800 108062 856
rect 108230 800 109166 856
rect 109334 800 110270 856
rect 110438 800 111374 856
rect 111542 800 112478 856
rect 112646 800 113490 856
rect 113658 800 114594 856
rect 114762 800 115698 856
rect 115866 800 116802 856
rect 116970 800 117906 856
rect 118074 800 119010 856
rect 119178 800 120022 856
rect 120190 800 121126 856
rect 121294 800 122230 856
rect 122398 800 123334 856
rect 123502 800 124438 856
rect 124606 800 125542 856
rect 125710 800 126554 856
rect 126722 800 127658 856
rect 127826 800 128762 856
rect 128930 800 129866 856
rect 130034 800 130970 856
rect 131138 800 131982 856
rect 132150 800 133086 856
rect 133254 800 134190 856
rect 134358 800 135294 856
rect 135462 800 136398 856
rect 136566 800 137502 856
rect 137670 800 138514 856
rect 138682 800 139618 856
rect 139786 800 140722 856
rect 140890 800 141826 856
rect 141994 800 142930 856
rect 143098 800 144034 856
rect 144202 800 145046 856
rect 145214 800 146150 856
rect 146318 800 147254 856
rect 147422 800 148358 856
rect 148526 800 149462 856
rect 149630 800 150566 856
rect 150734 800 151578 856
rect 151746 800 152682 856
rect 152850 800 153786 856
rect 153954 800 154890 856
rect 155058 800 155994 856
rect 156162 800 157098 856
rect 157266 800 158110 856
rect 158278 800 159214 856
rect 159382 800 160318 856
rect 160486 800 161422 856
rect 161590 800 162526 856
rect 162694 800 163538 856
rect 163706 800 164642 856
rect 164810 800 165746 856
rect 165914 800 166850 856
rect 167018 800 167954 856
rect 168122 800 169058 856
rect 169226 800 170070 856
rect 170238 800 171174 856
rect 171342 800 172278 856
rect 172446 800 173382 856
rect 173550 800 174486 856
rect 174654 800 175590 856
rect 175758 800 176602 856
rect 176770 800 177706 856
rect 177874 800 178810 856
rect 178978 800 179914 856
rect 180082 800 181018 856
rect 181186 800 182122 856
rect 182290 800 183134 856
rect 183302 800 184238 856
rect 184406 800 185342 856
rect 185510 800 186446 856
rect 186614 800 187550 856
rect 187718 800 188562 856
rect 188730 800 189666 856
rect 189834 800 190770 856
rect 190938 800 191874 856
rect 192042 800 192978 856
rect 193146 800 194082 856
rect 194250 800 195094 856
rect 195262 800 196198 856
rect 196366 800 197302 856
rect 197470 800 198406 856
rect 198574 800 199510 856
rect 199678 800 200614 856
rect 200782 800 201626 856
rect 201794 800 202730 856
rect 202898 800 203834 856
rect 204002 800 204938 856
rect 205106 800 206042 856
rect 206210 800 207146 856
rect 207314 800 208158 856
rect 208326 800 209262 856
rect 209430 800 210366 856
rect 210534 800 211470 856
rect 211638 800 212574 856
rect 212742 800 213586 856
rect 213754 800 214690 856
rect 214858 800 215794 856
rect 215962 800 216898 856
rect 217066 800 218002 856
rect 218170 800 219106 856
rect 219274 800 220118 856
rect 220286 800 221222 856
rect 221390 800 222326 856
rect 222494 800 223430 856
rect 223598 800 224534 856
rect 224702 800 225638 856
rect 225806 800 226650 856
rect 226818 800 227754 856
rect 227922 800 228858 856
rect 229026 800 229962 856
rect 230130 800 231066 856
rect 231234 800 232170 856
rect 232338 800 233182 856
rect 233350 800 234286 856
rect 234454 800 235390 856
rect 235558 800 236494 856
rect 236662 800 237598 856
rect 237766 800 238610 856
rect 238778 800 239714 856
rect 239882 800 240818 856
rect 240986 800 241922 856
rect 242090 800 243026 856
rect 243194 800 244130 856
rect 244298 800 245142 856
rect 245310 800 246246 856
rect 246414 800 247350 856
rect 247518 800 248454 856
rect 248622 800 249558 856
rect 249726 800 250662 856
rect 250830 800 251674 856
rect 251842 800 252778 856
rect 252946 800 253882 856
rect 254050 800 254986 856
rect 255154 800 256090 856
rect 256258 800 257194 856
rect 257362 800 258206 856
rect 258374 800 259310 856
rect 259478 800 260414 856
rect 260582 800 261518 856
rect 261686 800 262622 856
rect 262790 800 263634 856
rect 263802 800 264738 856
rect 264906 800 265842 856
rect 266010 800 266946 856
rect 267114 800 268050 856
rect 268218 800 269154 856
rect 269322 800 270166 856
rect 270334 800 271270 856
rect 271438 800 272374 856
rect 272542 800 273478 856
rect 273646 800 274582 856
rect 274750 800 275686 856
rect 275854 800 276698 856
rect 276866 800 277802 856
rect 277970 800 278906 856
rect 279074 800 280010 856
rect 280178 800 281114 856
rect 281282 800 282218 856
rect 282386 800 283230 856
rect 283398 800 284334 856
rect 284502 800 285438 856
rect 285606 800 286542 856
rect 286710 800 287646 856
rect 287814 800 288750 856
rect 288918 800 289762 856
rect 289930 800 290866 856
rect 291034 800 291970 856
rect 292138 800 293074 856
rect 293242 800 294178 856
rect 294346 800 295190 856
rect 295358 800 296294 856
rect 296462 800 297398 856
rect 297566 800 298502 856
rect 298670 800 299606 856
rect 299774 800 300710 856
rect 300878 800 301722 856
rect 301890 800 302826 856
rect 302994 800 303930 856
rect 304098 800 305034 856
rect 305202 800 306138 856
rect 306306 800 307242 856
rect 307410 800 308254 856
rect 308422 800 309358 856
rect 309526 800 310462 856
rect 310630 800 311566 856
rect 311734 800 312670 856
rect 312838 800 313774 856
rect 313942 800 314786 856
rect 314954 800 315890 856
rect 316058 800 316994 856
rect 317162 800 318098 856
rect 318266 800 319202 856
rect 319370 800 320214 856
rect 320382 800 321318 856
rect 321486 800 322422 856
rect 322590 800 323526 856
rect 323694 800 324630 856
rect 324798 800 325734 856
rect 325902 800 326746 856
rect 326914 800 327850 856
rect 328018 800 328954 856
rect 329122 800 330058 856
rect 330226 800 331162 856
rect 331330 800 332266 856
rect 332434 800 333278 856
rect 333446 800 334382 856
rect 334550 800 335486 856
rect 335654 800 336590 856
rect 336758 800 337694 856
rect 337862 800 338798 856
rect 338966 800 339810 856
rect 339978 800 340914 856
rect 341082 800 342018 856
rect 342186 800 343122 856
rect 343290 800 344226 856
rect 344394 800 345238 856
rect 345406 800 346342 856
rect 346510 800 347446 856
rect 347614 800 348550 856
rect 348718 800 349654 856
rect 349822 800 350758 856
rect 350926 800 351770 856
rect 351938 800 352874 856
rect 353042 800 353978 856
rect 354146 800 355082 856
rect 355250 800 356186 856
rect 356354 800 357290 856
rect 357458 800 358302 856
rect 358470 800 359406 856
rect 359574 800 360510 856
rect 360678 800 361614 856
rect 361782 800 362718 856
rect 362886 800 363822 856
rect 363990 800 364834 856
rect 365002 800 365938 856
rect 366106 800 367042 856
rect 367210 800 368146 856
rect 368314 800 369250 856
rect 369418 800 370262 856
rect 370430 800 371366 856
rect 371534 800 372470 856
rect 372638 800 373574 856
rect 373742 800 374678 856
rect 374846 800 375782 856
rect 375950 800 376794 856
rect 376962 800 377898 856
rect 378066 800 379002 856
rect 379170 800 380106 856
rect 380274 800 381210 856
rect 381378 800 382314 856
rect 382482 800 383326 856
rect 383494 800 384430 856
rect 384598 800 385534 856
rect 385702 800 386638 856
rect 386806 800 387742 856
rect 387910 800 388846 856
rect 389014 800 389858 856
rect 390026 800 390962 856
rect 391130 800 392066 856
rect 392234 800 393170 856
rect 393338 800 394274 856
rect 394442 800 395286 856
rect 395454 800 396390 856
rect 396558 800 397494 856
rect 397662 800 398598 856
rect 398766 800 399702 856
rect 399870 800 400806 856
rect 400974 800 401818 856
rect 401986 800 402922 856
rect 403090 800 404026 856
rect 404194 800 405130 856
rect 405298 800 406234 856
rect 406402 800 407338 856
rect 407506 800 408350 856
rect 408518 800 409454 856
rect 409622 800 410558 856
rect 410726 800 411662 856
rect 411830 800 412766 856
rect 412934 800 413870 856
rect 414038 800 414882 856
rect 415050 800 415986 856
rect 416154 800 417090 856
rect 417258 800 418194 856
<< metal3 >>
rect 419200 494232 420000 494352
rect 0 493824 800 493944
rect 419200 483080 420000 483200
rect 0 481856 800 481976
rect 419200 471928 420000 472048
rect 0 470024 800 470144
rect 419200 460912 420000 461032
rect 0 458056 800 458176
rect 419200 449760 420000 449880
rect 0 446224 800 446344
rect 419200 438608 420000 438728
rect 0 434256 800 434376
rect 419200 427592 420000 427712
rect 0 422424 800 422544
rect 419200 416440 420000 416560
rect 0 410456 800 410576
rect 419200 405288 420000 405408
rect 0 398624 800 398744
rect 419200 394272 420000 394392
rect 0 386656 800 386776
rect 419200 383120 420000 383240
rect 0 374824 800 374944
rect 419200 371968 420000 372088
rect 0 362856 800 362976
rect 419200 360952 420000 361072
rect 0 351024 800 351144
rect 419200 349800 420000 349920
rect 0 339056 800 339176
rect 419200 338648 420000 338768
rect 419200 327496 420000 327616
rect 0 327224 800 327344
rect 419200 316480 420000 316600
rect 0 315256 800 315376
rect 419200 305328 420000 305448
rect 0 303424 800 303544
rect 419200 294176 420000 294296
rect 0 291456 800 291576
rect 419200 283160 420000 283280
rect 0 279624 800 279744
rect 419200 272008 420000 272128
rect 0 267656 800 267776
rect 419200 260856 420000 260976
rect 0 255824 800 255944
rect 419200 249840 420000 249960
rect 0 243856 800 243976
rect 419200 238688 420000 238808
rect 0 231888 800 232008
rect 419200 227536 420000 227656
rect 0 220056 800 220176
rect 419200 216520 420000 216640
rect 0 208088 800 208208
rect 419200 205368 420000 205488
rect 0 196256 800 196376
rect 419200 194216 420000 194336
rect 0 184288 800 184408
rect 419200 183200 420000 183320
rect 0 172456 800 172576
rect 419200 172048 420000 172168
rect 419200 160896 420000 161016
rect 0 160488 800 160608
rect 419200 149744 420000 149864
rect 0 148656 800 148776
rect 419200 138728 420000 138848
rect 0 136688 800 136808
rect 419200 127576 420000 127696
rect 0 124856 800 124976
rect 419200 116424 420000 116544
rect 0 112888 800 113008
rect 419200 105408 420000 105528
rect 0 101056 800 101176
rect 419200 94256 420000 94376
rect 0 89088 800 89208
rect 419200 83104 420000 83224
rect 0 77256 800 77376
rect 419200 72088 420000 72208
rect 0 65288 800 65408
rect 419200 60936 420000 61056
rect 0 53456 800 53576
rect 419200 49784 420000 49904
rect 0 41488 800 41608
rect 419200 38768 420000 38888
rect 0 29656 800 29776
rect 419200 27616 420000 27736
rect 0 17688 800 17808
rect 419200 16464 420000 16584
rect 0 5856 800 5976
rect 419200 5448 420000 5568
<< obsm3 >>
rect 800 494432 419200 497793
rect 800 494152 419120 494432
rect 800 494024 419200 494152
rect 880 493744 419200 494024
rect 800 483280 419200 493744
rect 800 483000 419120 483280
rect 800 482056 419200 483000
rect 880 481776 419200 482056
rect 800 472128 419200 481776
rect 800 471848 419120 472128
rect 800 470224 419200 471848
rect 880 469944 419200 470224
rect 800 461112 419200 469944
rect 800 460832 419120 461112
rect 800 458256 419200 460832
rect 880 457976 419200 458256
rect 800 449960 419200 457976
rect 800 449680 419120 449960
rect 800 446424 419200 449680
rect 880 446144 419200 446424
rect 800 438808 419200 446144
rect 800 438528 419120 438808
rect 800 434456 419200 438528
rect 880 434176 419200 434456
rect 800 427792 419200 434176
rect 800 427512 419120 427792
rect 800 422624 419200 427512
rect 880 422344 419200 422624
rect 800 416640 419200 422344
rect 800 416360 419120 416640
rect 800 410656 419200 416360
rect 880 410376 419200 410656
rect 800 405488 419200 410376
rect 800 405208 419120 405488
rect 800 398824 419200 405208
rect 880 398544 419200 398824
rect 800 394472 419200 398544
rect 800 394192 419120 394472
rect 800 386856 419200 394192
rect 880 386576 419200 386856
rect 800 383320 419200 386576
rect 800 383040 419120 383320
rect 800 375024 419200 383040
rect 880 374744 419200 375024
rect 800 372168 419200 374744
rect 800 371888 419120 372168
rect 800 363056 419200 371888
rect 880 362776 419200 363056
rect 800 361152 419200 362776
rect 800 360872 419120 361152
rect 800 351224 419200 360872
rect 880 350944 419200 351224
rect 800 350000 419200 350944
rect 800 349720 419120 350000
rect 800 339256 419200 349720
rect 880 338976 419200 339256
rect 800 338848 419200 338976
rect 800 338568 419120 338848
rect 800 327696 419200 338568
rect 800 327424 419120 327696
rect 880 327416 419120 327424
rect 880 327144 419200 327416
rect 800 316680 419200 327144
rect 800 316400 419120 316680
rect 800 315456 419200 316400
rect 880 315176 419200 315456
rect 800 305528 419200 315176
rect 800 305248 419120 305528
rect 800 303624 419200 305248
rect 880 303344 419200 303624
rect 800 294376 419200 303344
rect 800 294096 419120 294376
rect 800 291656 419200 294096
rect 880 291376 419200 291656
rect 800 283360 419200 291376
rect 800 283080 419120 283360
rect 800 279824 419200 283080
rect 880 279544 419200 279824
rect 800 272208 419200 279544
rect 800 271928 419120 272208
rect 800 267856 419200 271928
rect 880 267576 419200 267856
rect 800 261056 419200 267576
rect 800 260776 419120 261056
rect 800 256024 419200 260776
rect 880 255744 419200 256024
rect 800 250040 419200 255744
rect 800 249760 419120 250040
rect 800 244056 419200 249760
rect 880 243776 419200 244056
rect 800 238888 419200 243776
rect 800 238608 419120 238888
rect 800 232088 419200 238608
rect 880 231808 419200 232088
rect 800 227736 419200 231808
rect 800 227456 419120 227736
rect 800 220256 419200 227456
rect 880 219976 419200 220256
rect 800 216720 419200 219976
rect 800 216440 419120 216720
rect 800 208288 419200 216440
rect 880 208008 419200 208288
rect 800 205568 419200 208008
rect 800 205288 419120 205568
rect 800 196456 419200 205288
rect 880 196176 419200 196456
rect 800 194416 419200 196176
rect 800 194136 419120 194416
rect 800 184488 419200 194136
rect 880 184208 419200 184488
rect 800 183400 419200 184208
rect 800 183120 419120 183400
rect 800 172656 419200 183120
rect 880 172376 419200 172656
rect 800 172248 419200 172376
rect 800 171968 419120 172248
rect 800 161096 419200 171968
rect 800 160816 419120 161096
rect 800 160688 419200 160816
rect 880 160408 419200 160688
rect 800 149944 419200 160408
rect 800 149664 419120 149944
rect 800 148856 419200 149664
rect 880 148576 419200 148856
rect 800 138928 419200 148576
rect 800 138648 419120 138928
rect 800 136888 419200 138648
rect 880 136608 419200 136888
rect 800 127776 419200 136608
rect 800 127496 419120 127776
rect 800 125056 419200 127496
rect 880 124776 419200 125056
rect 800 116624 419200 124776
rect 800 116344 419120 116624
rect 800 113088 419200 116344
rect 880 112808 419200 113088
rect 800 105608 419200 112808
rect 800 105328 419120 105608
rect 800 101256 419200 105328
rect 880 100976 419200 101256
rect 800 94456 419200 100976
rect 800 94176 419120 94456
rect 800 89288 419200 94176
rect 880 89008 419200 89288
rect 800 83304 419200 89008
rect 800 83024 419120 83304
rect 800 77456 419200 83024
rect 880 77176 419200 77456
rect 800 72288 419200 77176
rect 800 72008 419120 72288
rect 800 65488 419200 72008
rect 880 65208 419200 65488
rect 800 61136 419200 65208
rect 800 60856 419120 61136
rect 800 53656 419200 60856
rect 880 53376 419200 53656
rect 800 49984 419200 53376
rect 800 49704 419120 49984
rect 800 41688 419200 49704
rect 880 41408 419200 41688
rect 800 38968 419200 41408
rect 800 38688 419120 38968
rect 800 29856 419200 38688
rect 880 29576 419200 29856
rect 800 27816 419200 29576
rect 800 27536 419120 27816
rect 800 17888 419200 27536
rect 880 17608 419200 17888
rect 800 16664 419200 17608
rect 800 16384 419120 16664
rect 800 6056 419200 16384
rect 880 5776 419200 6056
rect 800 5648 419200 5776
rect 800 5368 419120 5648
rect 800 851 419200 5368
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
<< obsm4 >>
rect 13307 2128 19488 497808
rect 19968 2128 415413 497808
<< labels >>
rlabel metal3 s 419200 5448 420000 5568 6 io_in[0]
port 1 nsew default input
rlabel metal3 s 419200 338648 420000 338768 6 io_in[10]
port 2 nsew default input
rlabel metal3 s 419200 371968 420000 372088 6 io_in[11]
port 3 nsew default input
rlabel metal3 s 419200 405288 420000 405408 6 io_in[12]
port 4 nsew default input
rlabel metal3 s 419200 438608 420000 438728 6 io_in[13]
port 5 nsew default input
rlabel metal3 s 419200 471928 420000 472048 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 412086 499200 412142 500000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 365442 499200 365498 500000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 318798 499200 318854 500000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 272154 499200 272210 500000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 225510 499200 225566 500000 6 io_in[19]
port 11 nsew default input
rlabel metal3 s 419200 38768 420000 38888 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 178774 499200 178830 500000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 132130 499200 132186 500000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 85486 499200 85542 500000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 38842 499200 38898 500000 6 io_in[23]
port 16 nsew default input
rlabel metal3 s 0 493824 800 493944 6 io_in[24]
port 17 nsew default input
rlabel metal3 s 0 458056 800 458176 6 io_in[25]
port 18 nsew default input
rlabel metal3 s 0 422424 800 422544 6 io_in[26]
port 19 nsew default input
rlabel metal3 s 0 386656 800 386776 6 io_in[27]
port 20 nsew default input
rlabel metal3 s 0 351024 800 351144 6 io_in[28]
port 21 nsew default input
rlabel metal3 s 0 315256 800 315376 6 io_in[29]
port 22 nsew default input
rlabel metal3 s 419200 72088 420000 72208 6 io_in[2]
port 23 nsew default input
rlabel metal3 s 0 279624 800 279744 6 io_in[30]
port 24 nsew default input
rlabel metal3 s 0 243856 800 243976 6 io_in[31]
port 25 nsew default input
rlabel metal3 s 0 208088 800 208208 6 io_in[32]
port 26 nsew default input
rlabel metal3 s 0 172456 800 172576 6 io_in[33]
port 27 nsew default input
rlabel metal3 s 0 136688 800 136808 6 io_in[34]
port 28 nsew default input
rlabel metal3 s 0 101056 800 101176 6 io_in[35]
port 29 nsew default input
rlabel metal3 s 0 65288 800 65408 6 io_in[36]
port 30 nsew default input
rlabel metal3 s 0 29656 800 29776 6 io_in[37]
port 31 nsew default input
rlabel metal3 s 419200 105408 420000 105528 6 io_in[3]
port 32 nsew default input
rlabel metal3 s 419200 138728 420000 138848 6 io_in[4]
port 33 nsew default input
rlabel metal3 s 419200 172048 420000 172168 6 io_in[5]
port 34 nsew default input
rlabel metal3 s 419200 205368 420000 205488 6 io_in[6]
port 35 nsew default input
rlabel metal3 s 419200 238688 420000 238808 6 io_in[7]
port 36 nsew default input
rlabel metal3 s 419200 272008 420000 272128 6 io_in[8]
port 37 nsew default input
rlabel metal3 s 419200 305328 420000 305448 6 io_in[9]
port 38 nsew default input
rlabel metal3 s 419200 27616 420000 27736 6 io_oeb[0]
port 39 nsew default output
rlabel metal3 s 419200 360952 420000 361072 6 io_oeb[10]
port 40 nsew default output
rlabel metal3 s 419200 394272 420000 394392 6 io_oeb[11]
port 41 nsew default output
rlabel metal3 s 419200 427592 420000 427712 6 io_oeb[12]
port 42 nsew default output
rlabel metal3 s 419200 460912 420000 461032 6 io_oeb[13]
port 43 nsew default output
rlabel metal3 s 419200 494232 420000 494352 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 380990 499200 381046 500000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 334346 499200 334402 500000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 287702 499200 287758 500000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 241058 499200 241114 500000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 194322 499200 194378 500000 6 io_oeb[19]
port 49 nsew default output
rlabel metal3 s 419200 60936 420000 61056 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 147678 499200 147734 500000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 101034 499200 101090 500000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 54390 499200 54446 500000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 7746 499200 7802 500000 6 io_oeb[23]
port 54 nsew default output
rlabel metal3 s 0 470024 800 470144 6 io_oeb[24]
port 55 nsew default output
rlabel metal3 s 0 434256 800 434376 6 io_oeb[25]
port 56 nsew default output
rlabel metal3 s 0 398624 800 398744 6 io_oeb[26]
port 57 nsew default output
rlabel metal3 s 0 362856 800 362976 6 io_oeb[27]
port 58 nsew default output
rlabel metal3 s 0 327224 800 327344 6 io_oeb[28]
port 59 nsew default output
rlabel metal3 s 0 291456 800 291576 6 io_oeb[29]
port 60 nsew default output
rlabel metal3 s 419200 94256 420000 94376 6 io_oeb[2]
port 61 nsew default output
rlabel metal3 s 0 255824 800 255944 6 io_oeb[30]
port 62 nsew default output
rlabel metal3 s 0 220056 800 220176 6 io_oeb[31]
port 63 nsew default output
rlabel metal3 s 0 184288 800 184408 6 io_oeb[32]
port 64 nsew default output
rlabel metal3 s 0 148656 800 148776 6 io_oeb[33]
port 65 nsew default output
rlabel metal3 s 0 112888 800 113008 6 io_oeb[34]
port 66 nsew default output
rlabel metal3 s 0 77256 800 77376 6 io_oeb[35]
port 67 nsew default output
rlabel metal3 s 0 41488 800 41608 6 io_oeb[36]
port 68 nsew default output
rlabel metal3 s 0 5856 800 5976 6 io_oeb[37]
port 69 nsew default output
rlabel metal3 s 419200 127576 420000 127696 6 io_oeb[3]
port 70 nsew default output
rlabel metal3 s 419200 160896 420000 161016 6 io_oeb[4]
port 71 nsew default output
rlabel metal3 s 419200 194216 420000 194336 6 io_oeb[5]
port 72 nsew default output
rlabel metal3 s 419200 227536 420000 227656 6 io_oeb[6]
port 73 nsew default output
rlabel metal3 s 419200 260856 420000 260976 6 io_oeb[7]
port 74 nsew default output
rlabel metal3 s 419200 294176 420000 294296 6 io_oeb[8]
port 75 nsew default output
rlabel metal3 s 419200 327496 420000 327616 6 io_oeb[9]
port 76 nsew default output
rlabel metal3 s 419200 16464 420000 16584 6 io_out[0]
port 77 nsew default output
rlabel metal3 s 419200 349800 420000 349920 6 io_out[10]
port 78 nsew default output
rlabel metal3 s 419200 383120 420000 383240 6 io_out[11]
port 79 nsew default output
rlabel metal3 s 419200 416440 420000 416560 6 io_out[12]
port 80 nsew default output
rlabel metal3 s 419200 449760 420000 449880 6 io_out[13]
port 81 nsew default output
rlabel metal3 s 419200 483080 420000 483200 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 396538 499200 396594 500000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 349894 499200 349950 500000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 303250 499200 303306 500000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 256606 499200 256662 500000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 209870 499200 209926 500000 6 io_out[19]
port 87 nsew default output
rlabel metal3 s 419200 49784 420000 49904 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 163226 499200 163282 500000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 116582 499200 116638 500000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 69938 499200 69994 500000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 23294 499200 23350 500000 6 io_out[23]
port 92 nsew default output
rlabel metal3 s 0 481856 800 481976 6 io_out[24]
port 93 nsew default output
rlabel metal3 s 0 446224 800 446344 6 io_out[25]
port 94 nsew default output
rlabel metal3 s 0 410456 800 410576 6 io_out[26]
port 95 nsew default output
rlabel metal3 s 0 374824 800 374944 6 io_out[27]
port 96 nsew default output
rlabel metal3 s 0 339056 800 339176 6 io_out[28]
port 97 nsew default output
rlabel metal3 s 0 303424 800 303544 6 io_out[29]
port 98 nsew default output
rlabel metal3 s 419200 83104 420000 83224 6 io_out[2]
port 99 nsew default output
rlabel metal3 s 0 267656 800 267776 6 io_out[30]
port 100 nsew default output
rlabel metal3 s 0 231888 800 232008 6 io_out[31]
port 101 nsew default output
rlabel metal3 s 0 196256 800 196376 6 io_out[32]
port 102 nsew default output
rlabel metal3 s 0 160488 800 160608 6 io_out[33]
port 103 nsew default output
rlabel metal3 s 0 124856 800 124976 6 io_out[34]
port 104 nsew default output
rlabel metal3 s 0 89088 800 89208 6 io_out[35]
port 105 nsew default output
rlabel metal3 s 0 53456 800 53576 6 io_out[36]
port 106 nsew default output
rlabel metal3 s 0 17688 800 17808 6 io_out[37]
port 107 nsew default output
rlabel metal3 s 419200 116424 420000 116544 6 io_out[3]
port 108 nsew default output
rlabel metal3 s 419200 149744 420000 149864 6 io_out[4]
port 109 nsew default output
rlabel metal3 s 419200 183200 420000 183320 6 io_out[5]
port 110 nsew default output
rlabel metal3 s 419200 216520 420000 216640 6 io_out[6]
port 111 nsew default output
rlabel metal3 s 419200 249840 420000 249960 6 io_out[7]
port 112 nsew default output
rlabel metal3 s 419200 283160 420000 283280 6 io_out[8]
port 113 nsew default output
rlabel metal3 s 419200 316480 420000 316600 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 2594 0 2650 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 329010 0 329066 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 332322 0 332378 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 335542 0 335598 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 338854 0 338910 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 342074 0 342130 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 345294 0 345350 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 348606 0 348662 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 351826 0 351882 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 355138 0 355194 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 358358 0 358414 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 361670 0 361726 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 364890 0 364946 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 368202 0 368258 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 371422 0 371478 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 374734 0 374790 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 377954 0 378010 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 381266 0 381322 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 384486 0 384542 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 387798 0 387854 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 391018 0 391074 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 394330 0 394386 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 397550 0 397606 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 400862 0 400918 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 404082 0 404138 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 407394 0 407450 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 410614 0 410670 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 413926 0 413982 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 417146 0 417202 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 5906 0 5962 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 9126 0 9182 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 12438 0 12494 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 15658 0 15714 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 172334 0 172390 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 182178 0 182234 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 195150 0 195206 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 18970 0 19026 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 198462 0 198518 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 201682 0 201738 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 204994 0 205050 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 214746 0 214802 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 218058 0 218114 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 221278 0 221334 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 224590 0 224646 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 227810 0 227866 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 237654 0 237710 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 240874 0 240930 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 244186 0 244242 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 247406 0 247462 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 250718 0 250774 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 260470 0 260526 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 25502 0 25558 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 263690 0 263746 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 267002 0 267058 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 270222 0 270278 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 273534 0 273590 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 280066 0 280122 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 283286 0 283342 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 286598 0 286654 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 289818 0 289874 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 293130 0 293186 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 28722 0 28778 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 296350 0 296406 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 299662 0 299718 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 302882 0 302938 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 309414 0 309470 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 312726 0 312782 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 315946 0 316002 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 319258 0 319314 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 322478 0 322534 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 325790 0 325846 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 3698 0 3754 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 330114 0 330170 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 336646 0 336702 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 339866 0 339922 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 343178 0 343234 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 346398 0 346454 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 349710 0 349766 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 352930 0 352986 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 356242 0 356298 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 359462 0 359518 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 362774 0 362830 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 365994 0 366050 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 369306 0 369362 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 372526 0 372582 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 375838 0 375894 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 379058 0 379114 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 382370 0 382426 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 385590 0 385646 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 388902 0 388958 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 392122 0 392178 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 395342 0 395398 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 398654 0 398710 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 401874 0 401930 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 405186 0 405242 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 408406 0 408462 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 411718 0 411774 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 414938 0 414994 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 418250 0 418306 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 6918 0 6974 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 10230 0 10286 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 13450 0 13506 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 157154 0 157210 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 16762 0 16818 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 176658 0 176714 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 189722 0 189778 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 193034 0 193090 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 19982 0 20038 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 199566 0 199622 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 202786 0 202842 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 206098 0 206154 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 215850 0 215906 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 222382 0 222438 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 225694 0 225750 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 23294 0 23350 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 235446 0 235502 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 238666 0 238722 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 241978 0 242034 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 245198 0 245254 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 248510 0 248566 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 255042 0 255098 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 258262 0 258318 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 261574 0 261630 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 264794 0 264850 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 268106 0 268162 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 274638 0 274694 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 281170 0 281226 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 284390 0 284446 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 287702 0 287758 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 290922 0 290978 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 294234 0 294290 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 297454 0 297510 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 300766 0 300822 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 303986 0 304042 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 307298 0 307354 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 310518 0 310574 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 313830 0 313886 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 317050 0 317106 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 320270 0 320326 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 323582 0 323638 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 326802 0 326858 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 4802 0 4858 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 331218 0 331274 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 334438 0 334494 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 337750 0 337806 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 340970 0 341026 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 344282 0 344338 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 347502 0 347558 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 350814 0 350870 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 354034 0 354090 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 357346 0 357402 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 360566 0 360622 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 37462 0 37518 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 363878 0 363934 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 367098 0 367154 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 370318 0 370374 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 373630 0 373686 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 376850 0 376906 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 380162 0 380218 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 383382 0 383438 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 386694 0 386750 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 389914 0 389970 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 393226 0 393282 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 40682 0 40738 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 396446 0 396502 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 399758 0 399814 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 402978 0 403034 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 406290 0 406346 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 409510 0 409566 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 412822 0 412878 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 416042 0 416098 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 419354 0 419410 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 43994 0 44050 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 47214 0 47270 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 50526 0 50582 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 53746 0 53802 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 56966 0 57022 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 60278 0 60334 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 63498 0 63554 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 66810 0 66866 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 8022 0 8078 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 70030 0 70086 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 73342 0 73398 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 76562 0 76618 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 79874 0 79930 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 83094 0 83150 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 86406 0 86462 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 89626 0 89682 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 92938 0 92994 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 96158 0 96214 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 99470 0 99526 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 11334 0 11390 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 102690 0 102746 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 106002 0 106058 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 109222 0 109278 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 112534 0 112590 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 115754 0 115810 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 119066 0 119122 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 122286 0 122342 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 125598 0 125654 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 128818 0 128874 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 132038 0 132094 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 14554 0 14610 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 135350 0 135406 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 138570 0 138626 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 141882 0 141938 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 145102 0 145158 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 148414 0 148470 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 151634 0 151690 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 154946 0 155002 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 158166 0 158222 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 161478 0 161534 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 164698 0 164754 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 17866 0 17922 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 168010 0 168066 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 171230 0 171286 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 174542 0 174598 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 177762 0 177818 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 181074 0 181130 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 184294 0 184350 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 187606 0 187662 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 190826 0 190882 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 194138 0 194194 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 197358 0 197414 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 21086 0 21142 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 200670 0 200726 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 203890 0 203946 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 207202 0 207258 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 210422 0 210478 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 213642 0 213698 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 216954 0 217010 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 220174 0 220230 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 223486 0 223542 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 226706 0 226762 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 230018 0 230074 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 24398 0 24454 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 233238 0 233294 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 236550 0 236606 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 239770 0 239826 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 243082 0 243138 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 246302 0 246358 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 249614 0 249670 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 252834 0 252890 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 256146 0 256202 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 259366 0 259422 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 262678 0 262734 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 27618 0 27674 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 265898 0 265954 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 269210 0 269266 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 272430 0 272486 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 275742 0 275798 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 278962 0 279018 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 282274 0 282330 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 285494 0 285550 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 288806 0 288862 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 292026 0 292082 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 295246 0 295302 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 30930 0 30986 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 298558 0 298614 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 301778 0 301834 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 305090 0 305146 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 308310 0 308366 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 311622 0 311678 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 314842 0 314898 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 318154 0 318210 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 321374 0 321430 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 324686 0 324742 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 327906 0 327962 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 34150 0 34206 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 500 nsew default input
rlabel metal4 s 4208 2128 4528 497808 6 VPWR
port 501 nsew power input
rlabel metal4 s 19568 2128 19888 497808 6 VGND
port 502 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 420000 500000
string LEFview TRUE
<< end >>
