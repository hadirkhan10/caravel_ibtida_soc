VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Ibtida_top_dffram_cv
  CLASS BLOCK ;
  FOREIGN Ibtida_top_dffram_cv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2100.000 BY 2300.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 2296.000 179.770 2300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 869.080 2100.000 869.680 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1644.130 2296.000 1644.410 2300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1587.090 0.000 1587.370 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.170 2296.000 298.450 2300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1263.250 2296.000 1263.530 2300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1896.210 0.000 1896.490 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.210 2296.000 930.490 2300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 516.840 2100.000 517.440 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1609.170 2296.000 1609.450 2300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2062.730 0.000 2063.010 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 4.000 778.560 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1059.480 4.000 1060.080 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1766.680 2100.000 1767.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2275.320 4.000 2275.920 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1860.330 0.000 1860.610 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.250 2296.000 918.530 2300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.010 2296.000 1013.290 2300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.410 2296.000 870.690 2300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1819.720 2100.000 1820.320 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2037.890 2296.000 2038.170 2300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1274.360 2100.000 1274.960 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2225.000 2100.000 2225.600 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1227.370 2296.000 1227.650 2300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.250 2296.000 251.530 2300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 512.530 2296.000 512.810 2300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1256.680 2100.000 1257.280 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2012.840 2100.000 2013.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1009.160 2100.000 1009.760 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 536.450 2296.000 536.730 2300.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 217.640 2100.000 218.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 973.800 2100.000 974.400 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.170 2296.000 620.450 2300.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1977.480 2100.000 1978.080 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1525.450 2296.000 1525.730 2300.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1598.130 0.000 1598.410 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2260.360 2100.000 2260.960 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1906.330 2296.000 1906.610 2300.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1920.130 0.000 1920.410 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.450 2296.000 1180.730 2300.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.290 2296.000 239.570 2300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 2296.000 60.170 2300.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.610 2296.000 143.890 2300.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1343.720 2100.000 1344.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2002.010 2296.000 2002.290 2300.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 691.930 2296.000 692.210 2300.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2096.770 2296.000 2097.050 2300.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1014.850 0.000 1015.130 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1715.890 2296.000 1716.170 2300.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 572.330 2296.000 572.610 2300.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 477.570 2296.000 477.850 2300.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1479.450 0.000 1479.730 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1203.640 2100.000 1204.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2065.880 2100.000 2066.480 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.160 4.000 2063.760 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.090 2296.000 1311.370 2300.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1193.330 0.000 1193.610 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1729.690 0.000 1729.970 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1396.760 2100.000 1397.360 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1781.640 4.000 1782.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 584.290 2296.000 584.570 2300.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.920 4.000 1201.520 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2154.280 2100.000 2154.880 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 2296.000 989.370 2300.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 393.080 2100.000 393.680 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1358.930 2296.000 1359.210 2300.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.290 2296.000 906.570 2300.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 417.770 2296.000 418.050 2300.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 499.160 2100.000 499.760 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1429.400 4.000 1430.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2118.920 2100.000 2119.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1394.810 2296.000 1395.090 2300.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 780.680 2100.000 781.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1763.730 2296.000 1764.010 2300.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1181.370 0.000 1181.650 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 310.130 2296.000 310.410 2300.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 340.040 2100.000 340.640 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 5.480 2100.000 6.080 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 703.890 2296.000 704.170 2300.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1870.450 2296.000 1870.730 2300.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.770 2296.000 1430.050 2300.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1657.930 0.000 1658.210 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 639.240 2100.000 639.840 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1990.050 2296.000 1990.330 2300.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1728.600 4.000 1729.200 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1765.570 0.000 1765.850 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1884.250 0.000 1884.530 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.810 2296.000 728.090 2300.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1585.250 2296.000 1585.530 2300.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 2296.000 72.130 2300.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1940.760 4.000 1941.360 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1852.360 4.000 1852.960 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 922.120 2100.000 922.720 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2039.730 0.000 2040.010 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1749.000 2100.000 1749.600 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 2296.000 131.930 2300.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2278.040 2100.000 2278.640 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.450 2296.000 858.730 2300.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.410 2296.000 548.690 2300.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.770 2296.000 1752.050 2300.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 481.480 2100.000 482.080 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1383.770 0.000 1384.050 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2083.560 2100.000 2084.160 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1150.600 2100.000 1151.200 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1502.840 2100.000 1503.440 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.810 2296.000 751.090 2300.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.760 4.000 1465.360 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 463.800 2100.000 464.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.010 2296.000 668.290 2300.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1641.560 4.000 1642.160 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2136.600 2100.000 2137.200 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 939.800 2100.000 940.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1713.640 2100.000 1714.240 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.570 2296.000 1489.850 2300.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1923.080 4.000 1923.680 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2222.280 4.000 2222.880 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1872.760 2100.000 1873.360 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1608.920 2100.000 1609.520 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1976.120 4.000 1976.720 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1323.050 2296.000 1323.330 2300.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2186.920 4.000 2187.520 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 410.760 2100.000 411.360 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.970 2296.000 1347.250 2300.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 2296.000 48.210 2300.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1681.850 0.000 1682.130 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1513.490 2296.000 1513.770 2300.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1660.600 2100.000 1661.200 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 919.400 4.000 920.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1115.240 2100.000 1115.840 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1573.290 2296.000 1573.570 2300.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2013.970 2296.000 2014.250 2300.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2030.520 2100.000 2031.120 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2101.240 2100.000 2101.840 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1813.410 0.000 1813.690 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2003.850 0.000 2004.130 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1515.330 0.000 1515.610 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1621.130 2296.000 1621.410 2300.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 76.200 2100.000 76.800 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1561.330 2296.000 1561.610 2300.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.810 0.000 1349.090 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 886.760 2100.000 887.360 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2239.960 4.000 2240.560 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1817.000 4.000 1817.600 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2189.640 2100.000 2190.240 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.010 2296.000 1335.290 2300.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.410 2296.000 203.690 2300.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 453.650 2296.000 453.930 2300.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 745.320 2100.000 745.920 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 199.960 2100.000 200.560 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1872.290 0.000 1872.570 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1326.040 2100.000 1326.640 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1669.890 0.000 1670.170 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2051.690 0.000 2051.970 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2048.200 2100.000 2048.800 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.050 2296.000 1001.330 2300.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2080.840 4.000 2081.440 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1645.970 0.000 1646.250 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.370 2296.000 560.650 2300.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1979.930 0.000 1980.210 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.570 2296.000 822.850 2300.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1811.570 2296.000 1811.850 2300.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.000 4.000 1307.600 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.690 2296.000 441.970 2300.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 446.120 2100.000 446.720 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1905.400 4.000 1906.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1379.080 2100.000 1379.680 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1908.170 0.000 1908.450 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 40.840 2100.000 41.440 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1062.200 2100.000 1062.800 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2098.520 4.000 2099.120 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2027.800 4.000 2028.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1954.170 2296.000 1954.450 2300.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 2296.000 96.050 2300.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.090 0.000 1265.370 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1500.120 4.000 1500.720 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1859.410 2296.000 1859.690 2300.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2171.960 2100.000 2172.560 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1443.570 0.000 1443.850 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 763.000 2100.000 763.600 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1044.520 2100.000 1045.120 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.490 2296.000 846.770 2300.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.010 2296.000 346.290 2300.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1465.650 2296.000 1465.930 2300.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 428.440 2100.000 429.040 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.770 0.000 1039.050 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1239.330 2296.000 1239.610 2300.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1417.810 2296.000 1418.090 2300.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1944.050 0.000 1944.330 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.210 2296.000 608.490 2300.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1527.290 0.000 1527.570 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1695.960 2100.000 1696.560 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.770 2296.000 1085.050 2300.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1908.120 2100.000 1908.720 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 632.130 2296.000 632.410 2300.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1588.520 4.000 1589.120 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 674.600 2100.000 675.200 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1995.160 2100.000 1995.760 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1290.680 2100.000 1291.280 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1606.200 4.000 1606.800 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 851.400 2100.000 852.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 833.720 2100.000 834.320 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1623.880 4.000 1624.480 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1597.210 2296.000 1597.490 2300.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 534.520 2100.000 535.120 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 287.000 2100.000 287.600 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1573.560 2100.000 1574.160 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 2296.000 286.490 2300.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 2296.000 37.170 2300.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1668.050 2296.000 1668.330 2300.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1537.410 2296.000 1537.690 2300.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1308.360 2100.000 1308.960 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 774.730 2296.000 775.010 2300.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.730 2296.000 1097.010 2300.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2073.770 2296.000 2074.050 2300.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.930 2296.000 370.210 2300.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2151.560 4.000 2152.160 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1855.080 2100.000 1855.680 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1775.690 2296.000 1775.970 2300.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1382.850 2296.000 1383.130 2300.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 709.960 2100.000 710.560 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1731.320 2100.000 1731.920 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1967.970 0.000 1968.250 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1287.170 2296.000 1287.450 2300.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1097.560 2100.000 1098.160 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1633.090 2296.000 1633.370 2300.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1622.050 0.000 1622.330 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1048.890 2296.000 1049.170 2300.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1132.920 2100.000 1133.520 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1825.370 0.000 1825.650 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 93.880 2100.000 94.480 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 738.850 2296.000 739.130 2300.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2025.930 2296.000 2026.210 2300.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1705.770 0.000 1706.050 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 569.880 2100.000 570.480 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.930 0.000 1313.210 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1703.930 2296.000 1704.210 2300.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1185.960 2100.000 1186.560 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2204.600 4.000 2205.200 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 2296.000 13.250 2300.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1026.840 2100.000 1027.440 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 2296.000 786.970 2300.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 991.480 2100.000 992.080 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1991.890 0.000 1992.170 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.970 2296.000 358.250 2300.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1966.130 2296.000 1966.410 2300.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1894.370 2296.000 1894.650 2300.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 2296.000 108.010 2300.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1834.680 4.000 1835.280 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1678.280 2100.000 1678.880 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.810 2296.000 1073.090 2300.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1239.000 2100.000 1239.600 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 904.440 2100.000 905.040 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1784.360 2100.000 1784.960 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.170 2296.000 965.450 2300.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1432.120 2100.000 1432.720 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.130 2296.000 977.410 2300.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.530 2296.000 1501.810 2300.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.010 0.000 967.290 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2169.240 4.000 2169.840 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 715.850 2296.000 716.130 2300.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.490 2296.000 1168.770 2300.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 587.560 2100.000 588.160 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.250 2296.000 596.530 2300.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1441.730 2296.000 1442.010 2300.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 129.240 2100.000 129.840 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2027.770 0.000 2028.050 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2207.320 2100.000 2207.920 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 304.680 2100.000 305.280 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1727.850 2296.000 1728.130 2300.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 605.240 2100.000 605.840 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 692.280 2100.000 692.880 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1642.920 2100.000 1643.520 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.290 2296.000 1251.570 2300.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.720 4.000 1412.320 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1168.280 2100.000 1168.880 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.410 2296.000 1215.690 2300.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 375.400 2100.000 376.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1799.320 4.000 1799.920 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1555.880 2100.000 1556.480 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 58.520 2100.000 59.120 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 253.000 2100.000 253.600 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.530 0.000 1110.810 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1836.410 0.000 1836.690 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2074.690 0.000 2074.970 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.490 2296.000 501.770 2300.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 2296.000 334.330 2300.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 2296.000 119.970 2300.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.920 4.000 1711.520 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1591.240 2100.000 1591.840 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1925.800 2100.000 1926.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1847.450 2296.000 1847.730 2300.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1625.240 2100.000 1625.840 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2293.000 4.000 2293.600 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 164.600 2100.000 165.200 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1787.650 2296.000 1787.930 2300.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1485.160 2100.000 1485.760 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 727.640 2100.000 728.240 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.610 2296.000 1132.890 2300.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.210 2296.000 1275.490 2300.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.650 2296.000 798.930 2300.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.810 2296.000 1740.090 2300.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.930 0.000 991.210 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1361.400 2100.000 1362.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 2296.000 430.010 2300.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2049.850 2296.000 2050.130 2300.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 2296.000 394.130 2300.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1549.370 2296.000 1549.650 2300.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1993.800 4.000 1994.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1837.400 2100.000 1838.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 2296.000 465.890 2300.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2011.480 4.000 2012.080 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.930 2296.000 1037.210 2300.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 816.040 2100.000 816.640 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1882.410 2296.000 1882.690 2300.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1517.800 4.000 1518.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1376.360 4.000 1376.960 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1959.800 2100.000 1960.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2045.480 4.000 2046.080 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1477.610 2296.000 1477.890 2300.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1823.530 2296.000 1823.810 2300.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2133.880 4.000 2134.480 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 621.560 2100.000 622.160 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.170 0.000 896.450 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.490 2296.000 524.770 2300.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1120.650 2296.000 1120.930 2300.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1467.480 2100.000 1468.080 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.890 2296.000 382.170 2300.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2116.200 4.000 2116.800 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 2296.000 155.850 2300.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 357.720 2100.000 358.320 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 2296.000 1299.410 2300.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 656.920 2100.000 657.520 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1802.040 2100.000 1802.640 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2061.810 2296.000 2062.090 2300.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 182.280 2100.000 182.880 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1676.920 4.000 1677.520 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 111.560 2100.000 112.160 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.370 2296.000 882.650 2300.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 270.680 2100.000 271.280 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.200 4.000 1130.800 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1680.010 2296.000 1680.290 2300.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1801.450 0.000 1801.730 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.770 2296.000 1407.050 2300.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1753.610 0.000 1753.890 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 23.160 2100.000 23.760 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.160 4.000 1553.760 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1419.650 0.000 1419.930 4.000 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 2296.000 25.210 2300.000 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 894.330 2296.000 894.610 2300.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 4.000 1219.200 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1943.480 2100.000 1944.080 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 4.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1289.010 0.000 1289.290 4.000 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 2296.000 263.490 2300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 2296.000 84.090 2300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.530 2296.000 1156.810 2300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 2296.000 191.730 2300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.290 2296.000 1918.570 2300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.690 2296.000 1453.970 2300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 552.200 2100.000 552.800 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 4.000 1113.120 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.680 4.000 1359.280 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.850 2296.000 1061.130 2300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1978.090 2296.000 1978.370 2300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1447.080 4.000 1447.680 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 146.920 2100.000 147.520 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1538.200 2100.000 1538.800 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.970 2296.000 1025.250 2300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.050 2296.000 656.330 2300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1520.520 2100.000 1521.120 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1503.370 0.000 1503.650 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.690 2296.000 1108.970 2300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1717.730 0.000 1718.010 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 798.360 2100.000 798.960 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.890 0.000 1325.170 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.130 2296.000 954.410 2300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.490 0.000 1122.770 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.970 0.000 1301.250 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1575.130 0.000 1575.410 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.090 2296.000 322.370 2300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 943.090 0.000 943.370 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1289.320 4.000 1289.920 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1942.210 2296.000 1942.490 2300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1930.250 2296.000 1930.530 2300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 2242.680 2100.000 2243.280 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1691.970 2296.000 1692.250 2300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 2296.000 274.530 2300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1887.720 4.000 1888.320 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1191.490 2296.000 1191.770 2300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1414.440 2100.000 1415.040 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1449.800 2100.000 1450.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 2296.000 215.650 2300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 235.320 2100.000 235.920 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 322.360 2100.000 322.960 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1634.010 0.000 1634.290 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1221.320 2100.000 1221.920 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1763.960 4.000 1764.560 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1789.490 0.000 1789.770 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.450 2296.000 1203.730 2300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.530 2296.000 834.810 2300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1799.610 2296.000 1799.890 2300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.170 2296.000 942.450 2300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1848.370 0.000 1848.650 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.960 4.000 1254.560 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.330 2296.000 227.610 2300.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2085.730 2296.000 2086.010 2300.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1835.490 2296.000 1835.770 2300.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.530 2296.000 489.810 2300.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.770 2296.000 763.050 2300.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1563.170 0.000 1563.450 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.090 2296.000 644.370 2300.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1746.280 4.000 1746.880 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1890.440 2100.000 1891.040 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 810.610 2296.000 810.890 2300.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 2296.000 167.810 2300.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.970 2296.000 680.250 2300.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1656.090 2296.000 1656.370 2300.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.890 2296.000 1371.170 2300.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 405.810 2296.000 406.090 2300.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2257.640 4.000 2258.240 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1079.880 2100.000 1080.480 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.570 2296.000 1144.850 2300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2096.000 956.120 2100.000 956.720 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2287.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2287.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2094.380 2287.605 ;
      LAYER met1 ;
        RECT 5.520 4.460 2097.070 2295.640 ;
      LAYER met2 ;
        RECT 9.290 2295.720 12.690 2296.000 ;
        RECT 13.530 2295.720 24.650 2296.000 ;
        RECT 25.490 2295.720 36.610 2296.000 ;
        RECT 37.450 2295.720 47.650 2296.000 ;
        RECT 48.490 2295.720 59.610 2296.000 ;
        RECT 60.450 2295.720 71.570 2296.000 ;
        RECT 72.410 2295.720 83.530 2296.000 ;
        RECT 84.370 2295.720 95.490 2296.000 ;
        RECT 96.330 2295.720 107.450 2296.000 ;
        RECT 108.290 2295.720 119.410 2296.000 ;
        RECT 120.250 2295.720 131.370 2296.000 ;
        RECT 132.210 2295.720 143.330 2296.000 ;
        RECT 144.170 2295.720 155.290 2296.000 ;
        RECT 156.130 2295.720 167.250 2296.000 ;
        RECT 168.090 2295.720 179.210 2296.000 ;
        RECT 180.050 2295.720 191.170 2296.000 ;
        RECT 192.010 2295.720 203.130 2296.000 ;
        RECT 203.970 2295.720 215.090 2296.000 ;
        RECT 215.930 2295.720 227.050 2296.000 ;
        RECT 227.890 2295.720 239.010 2296.000 ;
        RECT 239.850 2295.720 250.970 2296.000 ;
        RECT 251.810 2295.720 262.930 2296.000 ;
        RECT 263.770 2295.720 273.970 2296.000 ;
        RECT 274.810 2295.720 285.930 2296.000 ;
        RECT 286.770 2295.720 297.890 2296.000 ;
        RECT 298.730 2295.720 309.850 2296.000 ;
        RECT 310.690 2295.720 321.810 2296.000 ;
        RECT 322.650 2295.720 333.770 2296.000 ;
        RECT 334.610 2295.720 345.730 2296.000 ;
        RECT 346.570 2295.720 357.690 2296.000 ;
        RECT 358.530 2295.720 369.650 2296.000 ;
        RECT 370.490 2295.720 381.610 2296.000 ;
        RECT 382.450 2295.720 393.570 2296.000 ;
        RECT 394.410 2295.720 405.530 2296.000 ;
        RECT 406.370 2295.720 417.490 2296.000 ;
        RECT 418.330 2295.720 429.450 2296.000 ;
        RECT 430.290 2295.720 441.410 2296.000 ;
        RECT 442.250 2295.720 453.370 2296.000 ;
        RECT 454.210 2295.720 465.330 2296.000 ;
        RECT 466.170 2295.720 477.290 2296.000 ;
        RECT 478.130 2295.720 489.250 2296.000 ;
        RECT 490.090 2295.720 501.210 2296.000 ;
        RECT 502.050 2295.720 512.250 2296.000 ;
        RECT 513.090 2295.720 524.210 2296.000 ;
        RECT 525.050 2295.720 536.170 2296.000 ;
        RECT 537.010 2295.720 548.130 2296.000 ;
        RECT 548.970 2295.720 560.090 2296.000 ;
        RECT 560.930 2295.720 572.050 2296.000 ;
        RECT 572.890 2295.720 584.010 2296.000 ;
        RECT 584.850 2295.720 595.970 2296.000 ;
        RECT 596.810 2295.720 607.930 2296.000 ;
        RECT 608.770 2295.720 619.890 2296.000 ;
        RECT 620.730 2295.720 631.850 2296.000 ;
        RECT 632.690 2295.720 643.810 2296.000 ;
        RECT 644.650 2295.720 655.770 2296.000 ;
        RECT 656.610 2295.720 667.730 2296.000 ;
        RECT 668.570 2295.720 679.690 2296.000 ;
        RECT 680.530 2295.720 691.650 2296.000 ;
        RECT 692.490 2295.720 703.610 2296.000 ;
        RECT 704.450 2295.720 715.570 2296.000 ;
        RECT 716.410 2295.720 727.530 2296.000 ;
        RECT 728.370 2295.720 738.570 2296.000 ;
        RECT 739.410 2295.720 750.530 2296.000 ;
        RECT 751.370 2295.720 762.490 2296.000 ;
        RECT 763.330 2295.720 774.450 2296.000 ;
        RECT 775.290 2295.720 786.410 2296.000 ;
        RECT 787.250 2295.720 798.370 2296.000 ;
        RECT 799.210 2295.720 810.330 2296.000 ;
        RECT 811.170 2295.720 822.290 2296.000 ;
        RECT 823.130 2295.720 834.250 2296.000 ;
        RECT 835.090 2295.720 846.210 2296.000 ;
        RECT 847.050 2295.720 858.170 2296.000 ;
        RECT 859.010 2295.720 870.130 2296.000 ;
        RECT 870.970 2295.720 882.090 2296.000 ;
        RECT 882.930 2295.720 894.050 2296.000 ;
        RECT 894.890 2295.720 906.010 2296.000 ;
        RECT 906.850 2295.720 917.970 2296.000 ;
        RECT 918.810 2295.720 929.930 2296.000 ;
        RECT 930.770 2295.720 941.890 2296.000 ;
        RECT 942.730 2295.720 953.850 2296.000 ;
        RECT 954.690 2295.720 964.890 2296.000 ;
        RECT 965.730 2295.720 976.850 2296.000 ;
        RECT 977.690 2295.720 988.810 2296.000 ;
        RECT 989.650 2295.720 1000.770 2296.000 ;
        RECT 1001.610 2295.720 1012.730 2296.000 ;
        RECT 1013.570 2295.720 1024.690 2296.000 ;
        RECT 1025.530 2295.720 1036.650 2296.000 ;
        RECT 1037.490 2295.720 1048.610 2296.000 ;
        RECT 1049.450 2295.720 1060.570 2296.000 ;
        RECT 1061.410 2295.720 1072.530 2296.000 ;
        RECT 1073.370 2295.720 1084.490 2296.000 ;
        RECT 1085.330 2295.720 1096.450 2296.000 ;
        RECT 1097.290 2295.720 1108.410 2296.000 ;
        RECT 1109.250 2295.720 1120.370 2296.000 ;
        RECT 1121.210 2295.720 1132.330 2296.000 ;
        RECT 1133.170 2295.720 1144.290 2296.000 ;
        RECT 1145.130 2295.720 1156.250 2296.000 ;
        RECT 1157.090 2295.720 1168.210 2296.000 ;
        RECT 1169.050 2295.720 1180.170 2296.000 ;
        RECT 1181.010 2295.720 1191.210 2296.000 ;
        RECT 1192.050 2295.720 1203.170 2296.000 ;
        RECT 1204.010 2295.720 1215.130 2296.000 ;
        RECT 1215.970 2295.720 1227.090 2296.000 ;
        RECT 1227.930 2295.720 1239.050 2296.000 ;
        RECT 1239.890 2295.720 1251.010 2296.000 ;
        RECT 1251.850 2295.720 1262.970 2296.000 ;
        RECT 1263.810 2295.720 1274.930 2296.000 ;
        RECT 1275.770 2295.720 1286.890 2296.000 ;
        RECT 1287.730 2295.720 1298.850 2296.000 ;
        RECT 1299.690 2295.720 1310.810 2296.000 ;
        RECT 1311.650 2295.720 1322.770 2296.000 ;
        RECT 1323.610 2295.720 1334.730 2296.000 ;
        RECT 1335.570 2295.720 1346.690 2296.000 ;
        RECT 1347.530 2295.720 1358.650 2296.000 ;
        RECT 1359.490 2295.720 1370.610 2296.000 ;
        RECT 1371.450 2295.720 1382.570 2296.000 ;
        RECT 1383.410 2295.720 1394.530 2296.000 ;
        RECT 1395.370 2295.720 1406.490 2296.000 ;
        RECT 1407.330 2295.720 1417.530 2296.000 ;
        RECT 1418.370 2295.720 1429.490 2296.000 ;
        RECT 1430.330 2295.720 1441.450 2296.000 ;
        RECT 1442.290 2295.720 1453.410 2296.000 ;
        RECT 1454.250 2295.720 1465.370 2296.000 ;
        RECT 1466.210 2295.720 1477.330 2296.000 ;
        RECT 1478.170 2295.720 1489.290 2296.000 ;
        RECT 1490.130 2295.720 1501.250 2296.000 ;
        RECT 1502.090 2295.720 1513.210 2296.000 ;
        RECT 1514.050 2295.720 1525.170 2296.000 ;
        RECT 1526.010 2295.720 1537.130 2296.000 ;
        RECT 1537.970 2295.720 1549.090 2296.000 ;
        RECT 1549.930 2295.720 1561.050 2296.000 ;
        RECT 1561.890 2295.720 1573.010 2296.000 ;
        RECT 1573.850 2295.720 1584.970 2296.000 ;
        RECT 1585.810 2295.720 1596.930 2296.000 ;
        RECT 1597.770 2295.720 1608.890 2296.000 ;
        RECT 1609.730 2295.720 1620.850 2296.000 ;
        RECT 1621.690 2295.720 1632.810 2296.000 ;
        RECT 1633.650 2295.720 1643.850 2296.000 ;
        RECT 1644.690 2295.720 1655.810 2296.000 ;
        RECT 1656.650 2295.720 1667.770 2296.000 ;
        RECT 1668.610 2295.720 1679.730 2296.000 ;
        RECT 1680.570 2295.720 1691.690 2296.000 ;
        RECT 1692.530 2295.720 1703.650 2296.000 ;
        RECT 1704.490 2295.720 1715.610 2296.000 ;
        RECT 1716.450 2295.720 1727.570 2296.000 ;
        RECT 1728.410 2295.720 1739.530 2296.000 ;
        RECT 1740.370 2295.720 1751.490 2296.000 ;
        RECT 1752.330 2295.720 1763.450 2296.000 ;
        RECT 1764.290 2295.720 1775.410 2296.000 ;
        RECT 1776.250 2295.720 1787.370 2296.000 ;
        RECT 1788.210 2295.720 1799.330 2296.000 ;
        RECT 1800.170 2295.720 1811.290 2296.000 ;
        RECT 1812.130 2295.720 1823.250 2296.000 ;
        RECT 1824.090 2295.720 1835.210 2296.000 ;
        RECT 1836.050 2295.720 1847.170 2296.000 ;
        RECT 1848.010 2295.720 1859.130 2296.000 ;
        RECT 1859.970 2295.720 1870.170 2296.000 ;
        RECT 1871.010 2295.720 1882.130 2296.000 ;
        RECT 1882.970 2295.720 1894.090 2296.000 ;
        RECT 1894.930 2295.720 1906.050 2296.000 ;
        RECT 1906.890 2295.720 1918.010 2296.000 ;
        RECT 1918.850 2295.720 1929.970 2296.000 ;
        RECT 1930.810 2295.720 1941.930 2296.000 ;
        RECT 1942.770 2295.720 1953.890 2296.000 ;
        RECT 1954.730 2295.720 1965.850 2296.000 ;
        RECT 1966.690 2295.720 1977.810 2296.000 ;
        RECT 1978.650 2295.720 1989.770 2296.000 ;
        RECT 1990.610 2295.720 2001.730 2296.000 ;
        RECT 2002.570 2295.720 2013.690 2296.000 ;
        RECT 2014.530 2295.720 2025.650 2296.000 ;
        RECT 2026.490 2295.720 2037.610 2296.000 ;
        RECT 2038.450 2295.720 2049.570 2296.000 ;
        RECT 2050.410 2295.720 2061.530 2296.000 ;
        RECT 2062.370 2295.720 2073.490 2296.000 ;
        RECT 2074.330 2295.720 2085.450 2296.000 ;
        RECT 2086.290 2295.720 2096.490 2296.000 ;
        RECT 9.290 4.280 2097.040 2295.720 ;
        RECT 9.290 4.000 13.610 4.280 ;
        RECT 14.450 4.000 25.570 4.280 ;
        RECT 26.410 4.000 37.530 4.280 ;
        RECT 38.370 4.000 49.490 4.280 ;
        RECT 50.330 4.000 61.450 4.280 ;
        RECT 62.290 4.000 73.410 4.280 ;
        RECT 74.250 4.000 85.370 4.280 ;
        RECT 86.210 4.000 97.330 4.280 ;
        RECT 98.170 4.000 109.290 4.280 ;
        RECT 110.130 4.000 121.250 4.280 ;
        RECT 122.090 4.000 133.210 4.280 ;
        RECT 134.050 4.000 145.170 4.280 ;
        RECT 146.010 4.000 157.130 4.280 ;
        RECT 157.970 4.000 169.090 4.280 ;
        RECT 169.930 4.000 181.050 4.280 ;
        RECT 181.890 4.000 193.010 4.280 ;
        RECT 193.850 4.000 204.970 4.280 ;
        RECT 205.810 4.000 216.930 4.280 ;
        RECT 217.770 4.000 228.890 4.280 ;
        RECT 229.730 4.000 239.930 4.280 ;
        RECT 240.770 4.000 251.890 4.280 ;
        RECT 252.730 4.000 263.850 4.280 ;
        RECT 264.690 4.000 275.810 4.280 ;
        RECT 276.650 4.000 287.770 4.280 ;
        RECT 288.610 4.000 299.730 4.280 ;
        RECT 300.570 4.000 311.690 4.280 ;
        RECT 312.530 4.000 323.650 4.280 ;
        RECT 324.490 4.000 335.610 4.280 ;
        RECT 336.450 4.000 347.570 4.280 ;
        RECT 348.410 4.000 359.530 4.280 ;
        RECT 360.370 4.000 371.490 4.280 ;
        RECT 372.330 4.000 383.450 4.280 ;
        RECT 384.290 4.000 395.410 4.280 ;
        RECT 396.250 4.000 407.370 4.280 ;
        RECT 408.210 4.000 419.330 4.280 ;
        RECT 420.170 4.000 431.290 4.280 ;
        RECT 432.130 4.000 443.250 4.280 ;
        RECT 444.090 4.000 455.210 4.280 ;
        RECT 456.050 4.000 466.250 4.280 ;
        RECT 467.090 4.000 478.210 4.280 ;
        RECT 479.050 4.000 490.170 4.280 ;
        RECT 491.010 4.000 502.130 4.280 ;
        RECT 502.970 4.000 514.090 4.280 ;
        RECT 514.930 4.000 526.050 4.280 ;
        RECT 526.890 4.000 538.010 4.280 ;
        RECT 538.850 4.000 549.970 4.280 ;
        RECT 550.810 4.000 561.930 4.280 ;
        RECT 562.770 4.000 573.890 4.280 ;
        RECT 574.730 4.000 585.850 4.280 ;
        RECT 586.690 4.000 597.810 4.280 ;
        RECT 598.650 4.000 609.770 4.280 ;
        RECT 610.610 4.000 621.730 4.280 ;
        RECT 622.570 4.000 633.690 4.280 ;
        RECT 634.530 4.000 645.650 4.280 ;
        RECT 646.490 4.000 657.610 4.280 ;
        RECT 658.450 4.000 669.570 4.280 ;
        RECT 670.410 4.000 681.530 4.280 ;
        RECT 682.370 4.000 692.570 4.280 ;
        RECT 693.410 4.000 704.530 4.280 ;
        RECT 705.370 4.000 716.490 4.280 ;
        RECT 717.330 4.000 728.450 4.280 ;
        RECT 729.290 4.000 740.410 4.280 ;
        RECT 741.250 4.000 752.370 4.280 ;
        RECT 753.210 4.000 764.330 4.280 ;
        RECT 765.170 4.000 776.290 4.280 ;
        RECT 777.130 4.000 788.250 4.280 ;
        RECT 789.090 4.000 800.210 4.280 ;
        RECT 801.050 4.000 812.170 4.280 ;
        RECT 813.010 4.000 824.130 4.280 ;
        RECT 824.970 4.000 836.090 4.280 ;
        RECT 836.930 4.000 848.050 4.280 ;
        RECT 848.890 4.000 860.010 4.280 ;
        RECT 860.850 4.000 871.970 4.280 ;
        RECT 872.810 4.000 883.930 4.280 ;
        RECT 884.770 4.000 895.890 4.280 ;
        RECT 896.730 4.000 907.850 4.280 ;
        RECT 908.690 4.000 918.890 4.280 ;
        RECT 919.730 4.000 930.850 4.280 ;
        RECT 931.690 4.000 942.810 4.280 ;
        RECT 943.650 4.000 954.770 4.280 ;
        RECT 955.610 4.000 966.730 4.280 ;
        RECT 967.570 4.000 978.690 4.280 ;
        RECT 979.530 4.000 990.650 4.280 ;
        RECT 991.490 4.000 1002.610 4.280 ;
        RECT 1003.450 4.000 1014.570 4.280 ;
        RECT 1015.410 4.000 1026.530 4.280 ;
        RECT 1027.370 4.000 1038.490 4.280 ;
        RECT 1039.330 4.000 1050.450 4.280 ;
        RECT 1051.290 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1074.370 4.280 ;
        RECT 1075.210 4.000 1086.330 4.280 ;
        RECT 1087.170 4.000 1098.290 4.280 ;
        RECT 1099.130 4.000 1110.250 4.280 ;
        RECT 1111.090 4.000 1122.210 4.280 ;
        RECT 1123.050 4.000 1134.170 4.280 ;
        RECT 1135.010 4.000 1145.210 4.280 ;
        RECT 1146.050 4.000 1157.170 4.280 ;
        RECT 1158.010 4.000 1169.130 4.280 ;
        RECT 1169.970 4.000 1181.090 4.280 ;
        RECT 1181.930 4.000 1193.050 4.280 ;
        RECT 1193.890 4.000 1205.010 4.280 ;
        RECT 1205.850 4.000 1216.970 4.280 ;
        RECT 1217.810 4.000 1228.930 4.280 ;
        RECT 1229.770 4.000 1240.890 4.280 ;
        RECT 1241.730 4.000 1252.850 4.280 ;
        RECT 1253.690 4.000 1264.810 4.280 ;
        RECT 1265.650 4.000 1276.770 4.280 ;
        RECT 1277.610 4.000 1288.730 4.280 ;
        RECT 1289.570 4.000 1300.690 4.280 ;
        RECT 1301.530 4.000 1312.650 4.280 ;
        RECT 1313.490 4.000 1324.610 4.280 ;
        RECT 1325.450 4.000 1336.570 4.280 ;
        RECT 1337.410 4.000 1348.530 4.280 ;
        RECT 1349.370 4.000 1360.490 4.280 ;
        RECT 1361.330 4.000 1371.530 4.280 ;
        RECT 1372.370 4.000 1383.490 4.280 ;
        RECT 1384.330 4.000 1395.450 4.280 ;
        RECT 1396.290 4.000 1407.410 4.280 ;
        RECT 1408.250 4.000 1419.370 4.280 ;
        RECT 1420.210 4.000 1431.330 4.280 ;
        RECT 1432.170 4.000 1443.290 4.280 ;
        RECT 1444.130 4.000 1455.250 4.280 ;
        RECT 1456.090 4.000 1467.210 4.280 ;
        RECT 1468.050 4.000 1479.170 4.280 ;
        RECT 1480.010 4.000 1491.130 4.280 ;
        RECT 1491.970 4.000 1503.090 4.280 ;
        RECT 1503.930 4.000 1515.050 4.280 ;
        RECT 1515.890 4.000 1527.010 4.280 ;
        RECT 1527.850 4.000 1538.970 4.280 ;
        RECT 1539.810 4.000 1550.930 4.280 ;
        RECT 1551.770 4.000 1562.890 4.280 ;
        RECT 1563.730 4.000 1574.850 4.280 ;
        RECT 1575.690 4.000 1586.810 4.280 ;
        RECT 1587.650 4.000 1597.850 4.280 ;
        RECT 1598.690 4.000 1609.810 4.280 ;
        RECT 1610.650 4.000 1621.770 4.280 ;
        RECT 1622.610 4.000 1633.730 4.280 ;
        RECT 1634.570 4.000 1645.690 4.280 ;
        RECT 1646.530 4.000 1657.650 4.280 ;
        RECT 1658.490 4.000 1669.610 4.280 ;
        RECT 1670.450 4.000 1681.570 4.280 ;
        RECT 1682.410 4.000 1693.530 4.280 ;
        RECT 1694.370 4.000 1705.490 4.280 ;
        RECT 1706.330 4.000 1717.450 4.280 ;
        RECT 1718.290 4.000 1729.410 4.280 ;
        RECT 1730.250 4.000 1741.370 4.280 ;
        RECT 1742.210 4.000 1753.330 4.280 ;
        RECT 1754.170 4.000 1765.290 4.280 ;
        RECT 1766.130 4.000 1777.250 4.280 ;
        RECT 1778.090 4.000 1789.210 4.280 ;
        RECT 1790.050 4.000 1801.170 4.280 ;
        RECT 1802.010 4.000 1813.130 4.280 ;
        RECT 1813.970 4.000 1825.090 4.280 ;
        RECT 1825.930 4.000 1836.130 4.280 ;
        RECT 1836.970 4.000 1848.090 4.280 ;
        RECT 1848.930 4.000 1860.050 4.280 ;
        RECT 1860.890 4.000 1872.010 4.280 ;
        RECT 1872.850 4.000 1883.970 4.280 ;
        RECT 1884.810 4.000 1895.930 4.280 ;
        RECT 1896.770 4.000 1907.890 4.280 ;
        RECT 1908.730 4.000 1919.850 4.280 ;
        RECT 1920.690 4.000 1931.810 4.280 ;
        RECT 1932.650 4.000 1943.770 4.280 ;
        RECT 1944.610 4.000 1955.730 4.280 ;
        RECT 1956.570 4.000 1967.690 4.280 ;
        RECT 1968.530 4.000 1979.650 4.280 ;
        RECT 1980.490 4.000 1991.610 4.280 ;
        RECT 1992.450 4.000 2003.570 4.280 ;
        RECT 2004.410 4.000 2015.530 4.280 ;
        RECT 2016.370 4.000 2027.490 4.280 ;
        RECT 2028.330 4.000 2039.450 4.280 ;
        RECT 2040.290 4.000 2051.410 4.280 ;
        RECT 2052.250 4.000 2062.450 4.280 ;
        RECT 2063.290 4.000 2074.410 4.280 ;
        RECT 2075.250 4.000 2086.370 4.280 ;
        RECT 2087.210 4.000 2097.040 4.280 ;
      LAYER met3 ;
        RECT 3.990 2279.040 2096.000 2287.685 ;
        RECT 3.990 2277.640 2095.600 2279.040 ;
        RECT 3.990 2276.320 2096.000 2277.640 ;
        RECT 4.400 2274.920 2096.000 2276.320 ;
        RECT 3.990 2261.360 2096.000 2274.920 ;
        RECT 3.990 2259.960 2095.600 2261.360 ;
        RECT 3.990 2258.640 2096.000 2259.960 ;
        RECT 4.400 2257.240 2096.000 2258.640 ;
        RECT 3.990 2243.680 2096.000 2257.240 ;
        RECT 3.990 2242.280 2095.600 2243.680 ;
        RECT 3.990 2240.960 2096.000 2242.280 ;
        RECT 4.400 2239.560 2096.000 2240.960 ;
        RECT 3.990 2226.000 2096.000 2239.560 ;
        RECT 3.990 2224.600 2095.600 2226.000 ;
        RECT 3.990 2223.280 2096.000 2224.600 ;
        RECT 4.400 2221.880 2096.000 2223.280 ;
        RECT 3.990 2208.320 2096.000 2221.880 ;
        RECT 3.990 2206.920 2095.600 2208.320 ;
        RECT 3.990 2205.600 2096.000 2206.920 ;
        RECT 4.400 2204.200 2096.000 2205.600 ;
        RECT 3.990 2190.640 2096.000 2204.200 ;
        RECT 3.990 2189.240 2095.600 2190.640 ;
        RECT 3.990 2187.920 2096.000 2189.240 ;
        RECT 4.400 2186.520 2096.000 2187.920 ;
        RECT 3.990 2172.960 2096.000 2186.520 ;
        RECT 3.990 2171.560 2095.600 2172.960 ;
        RECT 3.990 2170.240 2096.000 2171.560 ;
        RECT 4.400 2168.840 2096.000 2170.240 ;
        RECT 3.990 2155.280 2096.000 2168.840 ;
        RECT 3.990 2153.880 2095.600 2155.280 ;
        RECT 3.990 2152.560 2096.000 2153.880 ;
        RECT 4.400 2151.160 2096.000 2152.560 ;
        RECT 3.990 2137.600 2096.000 2151.160 ;
        RECT 3.990 2136.200 2095.600 2137.600 ;
        RECT 3.990 2134.880 2096.000 2136.200 ;
        RECT 4.400 2133.480 2096.000 2134.880 ;
        RECT 3.990 2119.920 2096.000 2133.480 ;
        RECT 3.990 2118.520 2095.600 2119.920 ;
        RECT 3.990 2117.200 2096.000 2118.520 ;
        RECT 4.400 2115.800 2096.000 2117.200 ;
        RECT 3.990 2102.240 2096.000 2115.800 ;
        RECT 3.990 2100.840 2095.600 2102.240 ;
        RECT 3.990 2099.520 2096.000 2100.840 ;
        RECT 4.400 2098.120 2096.000 2099.520 ;
        RECT 3.990 2084.560 2096.000 2098.120 ;
        RECT 3.990 2083.160 2095.600 2084.560 ;
        RECT 3.990 2081.840 2096.000 2083.160 ;
        RECT 4.400 2080.440 2096.000 2081.840 ;
        RECT 3.990 2066.880 2096.000 2080.440 ;
        RECT 3.990 2065.480 2095.600 2066.880 ;
        RECT 3.990 2064.160 2096.000 2065.480 ;
        RECT 4.400 2062.760 2096.000 2064.160 ;
        RECT 3.990 2049.200 2096.000 2062.760 ;
        RECT 3.990 2047.800 2095.600 2049.200 ;
        RECT 3.990 2046.480 2096.000 2047.800 ;
        RECT 4.400 2045.080 2096.000 2046.480 ;
        RECT 3.990 2031.520 2096.000 2045.080 ;
        RECT 3.990 2030.120 2095.600 2031.520 ;
        RECT 3.990 2028.800 2096.000 2030.120 ;
        RECT 4.400 2027.400 2096.000 2028.800 ;
        RECT 3.990 2013.840 2096.000 2027.400 ;
        RECT 3.990 2012.480 2095.600 2013.840 ;
        RECT 4.400 2012.440 2095.600 2012.480 ;
        RECT 4.400 2011.080 2096.000 2012.440 ;
        RECT 3.990 1996.160 2096.000 2011.080 ;
        RECT 3.990 1994.800 2095.600 1996.160 ;
        RECT 4.400 1994.760 2095.600 1994.800 ;
        RECT 4.400 1993.400 2096.000 1994.760 ;
        RECT 3.990 1978.480 2096.000 1993.400 ;
        RECT 3.990 1977.120 2095.600 1978.480 ;
        RECT 4.400 1977.080 2095.600 1977.120 ;
        RECT 4.400 1975.720 2096.000 1977.080 ;
        RECT 3.990 1960.800 2096.000 1975.720 ;
        RECT 3.990 1959.440 2095.600 1960.800 ;
        RECT 4.400 1959.400 2095.600 1959.440 ;
        RECT 4.400 1958.040 2096.000 1959.400 ;
        RECT 3.990 1944.480 2096.000 1958.040 ;
        RECT 3.990 1943.080 2095.600 1944.480 ;
        RECT 3.990 1941.760 2096.000 1943.080 ;
        RECT 4.400 1940.360 2096.000 1941.760 ;
        RECT 3.990 1926.800 2096.000 1940.360 ;
        RECT 3.990 1925.400 2095.600 1926.800 ;
        RECT 3.990 1924.080 2096.000 1925.400 ;
        RECT 4.400 1922.680 2096.000 1924.080 ;
        RECT 3.990 1909.120 2096.000 1922.680 ;
        RECT 3.990 1907.720 2095.600 1909.120 ;
        RECT 3.990 1906.400 2096.000 1907.720 ;
        RECT 4.400 1905.000 2096.000 1906.400 ;
        RECT 3.990 1891.440 2096.000 1905.000 ;
        RECT 3.990 1890.040 2095.600 1891.440 ;
        RECT 3.990 1888.720 2096.000 1890.040 ;
        RECT 4.400 1887.320 2096.000 1888.720 ;
        RECT 3.990 1873.760 2096.000 1887.320 ;
        RECT 3.990 1872.360 2095.600 1873.760 ;
        RECT 3.990 1871.040 2096.000 1872.360 ;
        RECT 4.400 1869.640 2096.000 1871.040 ;
        RECT 3.990 1856.080 2096.000 1869.640 ;
        RECT 3.990 1854.680 2095.600 1856.080 ;
        RECT 3.990 1853.360 2096.000 1854.680 ;
        RECT 4.400 1851.960 2096.000 1853.360 ;
        RECT 3.990 1838.400 2096.000 1851.960 ;
        RECT 3.990 1837.000 2095.600 1838.400 ;
        RECT 3.990 1835.680 2096.000 1837.000 ;
        RECT 4.400 1834.280 2096.000 1835.680 ;
        RECT 3.990 1820.720 2096.000 1834.280 ;
        RECT 3.990 1819.320 2095.600 1820.720 ;
        RECT 3.990 1818.000 2096.000 1819.320 ;
        RECT 4.400 1816.600 2096.000 1818.000 ;
        RECT 3.990 1803.040 2096.000 1816.600 ;
        RECT 3.990 1801.640 2095.600 1803.040 ;
        RECT 3.990 1800.320 2096.000 1801.640 ;
        RECT 4.400 1798.920 2096.000 1800.320 ;
        RECT 3.990 1785.360 2096.000 1798.920 ;
        RECT 3.990 1783.960 2095.600 1785.360 ;
        RECT 3.990 1782.640 2096.000 1783.960 ;
        RECT 4.400 1781.240 2096.000 1782.640 ;
        RECT 3.990 1767.680 2096.000 1781.240 ;
        RECT 3.990 1766.280 2095.600 1767.680 ;
        RECT 3.990 1764.960 2096.000 1766.280 ;
        RECT 4.400 1763.560 2096.000 1764.960 ;
        RECT 3.990 1750.000 2096.000 1763.560 ;
        RECT 3.990 1748.600 2095.600 1750.000 ;
        RECT 3.990 1747.280 2096.000 1748.600 ;
        RECT 4.400 1745.880 2096.000 1747.280 ;
        RECT 3.990 1732.320 2096.000 1745.880 ;
        RECT 3.990 1730.920 2095.600 1732.320 ;
        RECT 3.990 1729.600 2096.000 1730.920 ;
        RECT 4.400 1728.200 2096.000 1729.600 ;
        RECT 3.990 1714.640 2096.000 1728.200 ;
        RECT 3.990 1713.240 2095.600 1714.640 ;
        RECT 3.990 1711.920 2096.000 1713.240 ;
        RECT 4.400 1710.520 2096.000 1711.920 ;
        RECT 3.990 1696.960 2096.000 1710.520 ;
        RECT 3.990 1695.560 2095.600 1696.960 ;
        RECT 3.990 1694.240 2096.000 1695.560 ;
        RECT 4.400 1692.840 2096.000 1694.240 ;
        RECT 3.990 1679.280 2096.000 1692.840 ;
        RECT 3.990 1677.920 2095.600 1679.280 ;
        RECT 4.400 1677.880 2095.600 1677.920 ;
        RECT 4.400 1676.520 2096.000 1677.880 ;
        RECT 3.990 1661.600 2096.000 1676.520 ;
        RECT 3.990 1660.240 2095.600 1661.600 ;
        RECT 4.400 1660.200 2095.600 1660.240 ;
        RECT 4.400 1658.840 2096.000 1660.200 ;
        RECT 3.990 1643.920 2096.000 1658.840 ;
        RECT 3.990 1642.560 2095.600 1643.920 ;
        RECT 4.400 1642.520 2095.600 1642.560 ;
        RECT 4.400 1641.160 2096.000 1642.520 ;
        RECT 3.990 1626.240 2096.000 1641.160 ;
        RECT 3.990 1624.880 2095.600 1626.240 ;
        RECT 4.400 1624.840 2095.600 1624.880 ;
        RECT 4.400 1623.480 2096.000 1624.840 ;
        RECT 3.990 1609.920 2096.000 1623.480 ;
        RECT 3.990 1608.520 2095.600 1609.920 ;
        RECT 3.990 1607.200 2096.000 1608.520 ;
        RECT 4.400 1605.800 2096.000 1607.200 ;
        RECT 3.990 1592.240 2096.000 1605.800 ;
        RECT 3.990 1590.840 2095.600 1592.240 ;
        RECT 3.990 1589.520 2096.000 1590.840 ;
        RECT 4.400 1588.120 2096.000 1589.520 ;
        RECT 3.990 1574.560 2096.000 1588.120 ;
        RECT 3.990 1573.160 2095.600 1574.560 ;
        RECT 3.990 1571.840 2096.000 1573.160 ;
        RECT 4.400 1570.440 2096.000 1571.840 ;
        RECT 3.990 1556.880 2096.000 1570.440 ;
        RECT 3.990 1555.480 2095.600 1556.880 ;
        RECT 3.990 1554.160 2096.000 1555.480 ;
        RECT 4.400 1552.760 2096.000 1554.160 ;
        RECT 3.990 1539.200 2096.000 1552.760 ;
        RECT 3.990 1537.800 2095.600 1539.200 ;
        RECT 3.990 1536.480 2096.000 1537.800 ;
        RECT 4.400 1535.080 2096.000 1536.480 ;
        RECT 3.990 1521.520 2096.000 1535.080 ;
        RECT 3.990 1520.120 2095.600 1521.520 ;
        RECT 3.990 1518.800 2096.000 1520.120 ;
        RECT 4.400 1517.400 2096.000 1518.800 ;
        RECT 3.990 1503.840 2096.000 1517.400 ;
        RECT 3.990 1502.440 2095.600 1503.840 ;
        RECT 3.990 1501.120 2096.000 1502.440 ;
        RECT 4.400 1499.720 2096.000 1501.120 ;
        RECT 3.990 1486.160 2096.000 1499.720 ;
        RECT 3.990 1484.760 2095.600 1486.160 ;
        RECT 3.990 1483.440 2096.000 1484.760 ;
        RECT 4.400 1482.040 2096.000 1483.440 ;
        RECT 3.990 1468.480 2096.000 1482.040 ;
        RECT 3.990 1467.080 2095.600 1468.480 ;
        RECT 3.990 1465.760 2096.000 1467.080 ;
        RECT 4.400 1464.360 2096.000 1465.760 ;
        RECT 3.990 1450.800 2096.000 1464.360 ;
        RECT 3.990 1449.400 2095.600 1450.800 ;
        RECT 3.990 1448.080 2096.000 1449.400 ;
        RECT 4.400 1446.680 2096.000 1448.080 ;
        RECT 3.990 1433.120 2096.000 1446.680 ;
        RECT 3.990 1431.720 2095.600 1433.120 ;
        RECT 3.990 1430.400 2096.000 1431.720 ;
        RECT 4.400 1429.000 2096.000 1430.400 ;
        RECT 3.990 1415.440 2096.000 1429.000 ;
        RECT 3.990 1414.040 2095.600 1415.440 ;
        RECT 3.990 1412.720 2096.000 1414.040 ;
        RECT 4.400 1411.320 2096.000 1412.720 ;
        RECT 3.990 1397.760 2096.000 1411.320 ;
        RECT 3.990 1396.360 2095.600 1397.760 ;
        RECT 3.990 1395.040 2096.000 1396.360 ;
        RECT 4.400 1393.640 2096.000 1395.040 ;
        RECT 3.990 1380.080 2096.000 1393.640 ;
        RECT 3.990 1378.680 2095.600 1380.080 ;
        RECT 3.990 1377.360 2096.000 1378.680 ;
        RECT 4.400 1375.960 2096.000 1377.360 ;
        RECT 3.990 1362.400 2096.000 1375.960 ;
        RECT 3.990 1361.000 2095.600 1362.400 ;
        RECT 3.990 1359.680 2096.000 1361.000 ;
        RECT 4.400 1358.280 2096.000 1359.680 ;
        RECT 3.990 1344.720 2096.000 1358.280 ;
        RECT 3.990 1343.360 2095.600 1344.720 ;
        RECT 4.400 1343.320 2095.600 1343.360 ;
        RECT 4.400 1341.960 2096.000 1343.320 ;
        RECT 3.990 1327.040 2096.000 1341.960 ;
        RECT 3.990 1325.680 2095.600 1327.040 ;
        RECT 4.400 1325.640 2095.600 1325.680 ;
        RECT 4.400 1324.280 2096.000 1325.640 ;
        RECT 3.990 1309.360 2096.000 1324.280 ;
        RECT 3.990 1308.000 2095.600 1309.360 ;
        RECT 4.400 1307.960 2095.600 1308.000 ;
        RECT 4.400 1306.600 2096.000 1307.960 ;
        RECT 3.990 1291.680 2096.000 1306.600 ;
        RECT 3.990 1290.320 2095.600 1291.680 ;
        RECT 4.400 1290.280 2095.600 1290.320 ;
        RECT 4.400 1288.920 2096.000 1290.280 ;
        RECT 3.990 1275.360 2096.000 1288.920 ;
        RECT 3.990 1273.960 2095.600 1275.360 ;
        RECT 3.990 1272.640 2096.000 1273.960 ;
        RECT 4.400 1271.240 2096.000 1272.640 ;
        RECT 3.990 1257.680 2096.000 1271.240 ;
        RECT 3.990 1256.280 2095.600 1257.680 ;
        RECT 3.990 1254.960 2096.000 1256.280 ;
        RECT 4.400 1253.560 2096.000 1254.960 ;
        RECT 3.990 1240.000 2096.000 1253.560 ;
        RECT 3.990 1238.600 2095.600 1240.000 ;
        RECT 3.990 1237.280 2096.000 1238.600 ;
        RECT 4.400 1235.880 2096.000 1237.280 ;
        RECT 3.990 1222.320 2096.000 1235.880 ;
        RECT 3.990 1220.920 2095.600 1222.320 ;
        RECT 3.990 1219.600 2096.000 1220.920 ;
        RECT 4.400 1218.200 2096.000 1219.600 ;
        RECT 3.990 1204.640 2096.000 1218.200 ;
        RECT 3.990 1203.240 2095.600 1204.640 ;
        RECT 3.990 1201.920 2096.000 1203.240 ;
        RECT 4.400 1200.520 2096.000 1201.920 ;
        RECT 3.990 1186.960 2096.000 1200.520 ;
        RECT 3.990 1185.560 2095.600 1186.960 ;
        RECT 3.990 1184.240 2096.000 1185.560 ;
        RECT 4.400 1182.840 2096.000 1184.240 ;
        RECT 3.990 1169.280 2096.000 1182.840 ;
        RECT 3.990 1167.880 2095.600 1169.280 ;
        RECT 3.990 1166.560 2096.000 1167.880 ;
        RECT 4.400 1165.160 2096.000 1166.560 ;
        RECT 3.990 1151.600 2096.000 1165.160 ;
        RECT 3.990 1150.200 2095.600 1151.600 ;
        RECT 3.990 1148.880 2096.000 1150.200 ;
        RECT 4.400 1147.480 2096.000 1148.880 ;
        RECT 3.990 1133.920 2096.000 1147.480 ;
        RECT 3.990 1132.520 2095.600 1133.920 ;
        RECT 3.990 1131.200 2096.000 1132.520 ;
        RECT 4.400 1129.800 2096.000 1131.200 ;
        RECT 3.990 1116.240 2096.000 1129.800 ;
        RECT 3.990 1114.840 2095.600 1116.240 ;
        RECT 3.990 1113.520 2096.000 1114.840 ;
        RECT 4.400 1112.120 2096.000 1113.520 ;
        RECT 3.990 1098.560 2096.000 1112.120 ;
        RECT 3.990 1097.160 2095.600 1098.560 ;
        RECT 3.990 1095.840 2096.000 1097.160 ;
        RECT 4.400 1094.440 2096.000 1095.840 ;
        RECT 3.990 1080.880 2096.000 1094.440 ;
        RECT 3.990 1079.480 2095.600 1080.880 ;
        RECT 3.990 1078.160 2096.000 1079.480 ;
        RECT 4.400 1076.760 2096.000 1078.160 ;
        RECT 3.990 1063.200 2096.000 1076.760 ;
        RECT 3.990 1061.800 2095.600 1063.200 ;
        RECT 3.990 1060.480 2096.000 1061.800 ;
        RECT 4.400 1059.080 2096.000 1060.480 ;
        RECT 3.990 1045.520 2096.000 1059.080 ;
        RECT 3.990 1044.120 2095.600 1045.520 ;
        RECT 3.990 1042.800 2096.000 1044.120 ;
        RECT 4.400 1041.400 2096.000 1042.800 ;
        RECT 3.990 1027.840 2096.000 1041.400 ;
        RECT 3.990 1026.440 2095.600 1027.840 ;
        RECT 3.990 1025.120 2096.000 1026.440 ;
        RECT 4.400 1023.720 2096.000 1025.120 ;
        RECT 3.990 1010.160 2096.000 1023.720 ;
        RECT 3.990 1008.800 2095.600 1010.160 ;
        RECT 4.400 1008.760 2095.600 1008.800 ;
        RECT 4.400 1007.400 2096.000 1008.760 ;
        RECT 3.990 992.480 2096.000 1007.400 ;
        RECT 3.990 991.120 2095.600 992.480 ;
        RECT 4.400 991.080 2095.600 991.120 ;
        RECT 4.400 989.720 2096.000 991.080 ;
        RECT 3.990 974.800 2096.000 989.720 ;
        RECT 3.990 973.440 2095.600 974.800 ;
        RECT 4.400 973.400 2095.600 973.440 ;
        RECT 4.400 972.040 2096.000 973.400 ;
        RECT 3.990 957.120 2096.000 972.040 ;
        RECT 3.990 955.760 2095.600 957.120 ;
        RECT 4.400 955.720 2095.600 955.760 ;
        RECT 4.400 954.360 2096.000 955.720 ;
        RECT 3.990 940.800 2096.000 954.360 ;
        RECT 3.990 939.400 2095.600 940.800 ;
        RECT 3.990 938.080 2096.000 939.400 ;
        RECT 4.400 936.680 2096.000 938.080 ;
        RECT 3.990 923.120 2096.000 936.680 ;
        RECT 3.990 921.720 2095.600 923.120 ;
        RECT 3.990 920.400 2096.000 921.720 ;
        RECT 4.400 919.000 2096.000 920.400 ;
        RECT 3.990 905.440 2096.000 919.000 ;
        RECT 3.990 904.040 2095.600 905.440 ;
        RECT 3.990 902.720 2096.000 904.040 ;
        RECT 4.400 901.320 2096.000 902.720 ;
        RECT 3.990 887.760 2096.000 901.320 ;
        RECT 3.990 886.360 2095.600 887.760 ;
        RECT 3.990 885.040 2096.000 886.360 ;
        RECT 4.400 883.640 2096.000 885.040 ;
        RECT 3.990 870.080 2096.000 883.640 ;
        RECT 3.990 868.680 2095.600 870.080 ;
        RECT 3.990 867.360 2096.000 868.680 ;
        RECT 4.400 865.960 2096.000 867.360 ;
        RECT 3.990 852.400 2096.000 865.960 ;
        RECT 3.990 851.000 2095.600 852.400 ;
        RECT 3.990 849.680 2096.000 851.000 ;
        RECT 4.400 848.280 2096.000 849.680 ;
        RECT 3.990 834.720 2096.000 848.280 ;
        RECT 3.990 833.320 2095.600 834.720 ;
        RECT 3.990 832.000 2096.000 833.320 ;
        RECT 4.400 830.600 2096.000 832.000 ;
        RECT 3.990 817.040 2096.000 830.600 ;
        RECT 3.990 815.640 2095.600 817.040 ;
        RECT 3.990 814.320 2096.000 815.640 ;
        RECT 4.400 812.920 2096.000 814.320 ;
        RECT 3.990 799.360 2096.000 812.920 ;
        RECT 3.990 797.960 2095.600 799.360 ;
        RECT 3.990 796.640 2096.000 797.960 ;
        RECT 4.400 795.240 2096.000 796.640 ;
        RECT 3.990 781.680 2096.000 795.240 ;
        RECT 3.990 780.280 2095.600 781.680 ;
        RECT 3.990 778.960 2096.000 780.280 ;
        RECT 4.400 777.560 2096.000 778.960 ;
        RECT 3.990 764.000 2096.000 777.560 ;
        RECT 3.990 762.600 2095.600 764.000 ;
        RECT 3.990 761.280 2096.000 762.600 ;
        RECT 4.400 759.880 2096.000 761.280 ;
        RECT 3.990 746.320 2096.000 759.880 ;
        RECT 3.990 744.920 2095.600 746.320 ;
        RECT 3.990 743.600 2096.000 744.920 ;
        RECT 4.400 742.200 2096.000 743.600 ;
        RECT 3.990 728.640 2096.000 742.200 ;
        RECT 3.990 727.240 2095.600 728.640 ;
        RECT 3.990 725.920 2096.000 727.240 ;
        RECT 4.400 724.520 2096.000 725.920 ;
        RECT 3.990 710.960 2096.000 724.520 ;
        RECT 3.990 709.560 2095.600 710.960 ;
        RECT 3.990 708.240 2096.000 709.560 ;
        RECT 4.400 706.840 2096.000 708.240 ;
        RECT 3.990 693.280 2096.000 706.840 ;
        RECT 3.990 691.880 2095.600 693.280 ;
        RECT 3.990 690.560 2096.000 691.880 ;
        RECT 4.400 689.160 2096.000 690.560 ;
        RECT 3.990 675.600 2096.000 689.160 ;
        RECT 3.990 674.240 2095.600 675.600 ;
        RECT 4.400 674.200 2095.600 674.240 ;
        RECT 4.400 672.840 2096.000 674.200 ;
        RECT 3.990 657.920 2096.000 672.840 ;
        RECT 3.990 656.560 2095.600 657.920 ;
        RECT 4.400 656.520 2095.600 656.560 ;
        RECT 4.400 655.160 2096.000 656.520 ;
        RECT 3.990 640.240 2096.000 655.160 ;
        RECT 3.990 638.880 2095.600 640.240 ;
        RECT 4.400 638.840 2095.600 638.880 ;
        RECT 4.400 637.480 2096.000 638.840 ;
        RECT 3.990 622.560 2096.000 637.480 ;
        RECT 3.990 621.200 2095.600 622.560 ;
        RECT 4.400 621.160 2095.600 621.200 ;
        RECT 4.400 619.800 2096.000 621.160 ;
        RECT 3.990 606.240 2096.000 619.800 ;
        RECT 3.990 604.840 2095.600 606.240 ;
        RECT 3.990 603.520 2096.000 604.840 ;
        RECT 4.400 602.120 2096.000 603.520 ;
        RECT 3.990 588.560 2096.000 602.120 ;
        RECT 3.990 587.160 2095.600 588.560 ;
        RECT 3.990 585.840 2096.000 587.160 ;
        RECT 4.400 584.440 2096.000 585.840 ;
        RECT 3.990 570.880 2096.000 584.440 ;
        RECT 3.990 569.480 2095.600 570.880 ;
        RECT 3.990 568.160 2096.000 569.480 ;
        RECT 4.400 566.760 2096.000 568.160 ;
        RECT 3.990 553.200 2096.000 566.760 ;
        RECT 3.990 551.800 2095.600 553.200 ;
        RECT 3.990 550.480 2096.000 551.800 ;
        RECT 4.400 549.080 2096.000 550.480 ;
        RECT 3.990 535.520 2096.000 549.080 ;
        RECT 3.990 534.120 2095.600 535.520 ;
        RECT 3.990 532.800 2096.000 534.120 ;
        RECT 4.400 531.400 2096.000 532.800 ;
        RECT 3.990 517.840 2096.000 531.400 ;
        RECT 3.990 516.440 2095.600 517.840 ;
        RECT 3.990 515.120 2096.000 516.440 ;
        RECT 4.400 513.720 2096.000 515.120 ;
        RECT 3.990 500.160 2096.000 513.720 ;
        RECT 3.990 498.760 2095.600 500.160 ;
        RECT 3.990 497.440 2096.000 498.760 ;
        RECT 4.400 496.040 2096.000 497.440 ;
        RECT 3.990 482.480 2096.000 496.040 ;
        RECT 3.990 481.080 2095.600 482.480 ;
        RECT 3.990 479.760 2096.000 481.080 ;
        RECT 4.400 478.360 2096.000 479.760 ;
        RECT 3.990 464.800 2096.000 478.360 ;
        RECT 3.990 463.400 2095.600 464.800 ;
        RECT 3.990 462.080 2096.000 463.400 ;
        RECT 4.400 460.680 2096.000 462.080 ;
        RECT 3.990 447.120 2096.000 460.680 ;
        RECT 3.990 445.720 2095.600 447.120 ;
        RECT 3.990 444.400 2096.000 445.720 ;
        RECT 4.400 443.000 2096.000 444.400 ;
        RECT 3.990 429.440 2096.000 443.000 ;
        RECT 3.990 428.040 2095.600 429.440 ;
        RECT 3.990 426.720 2096.000 428.040 ;
        RECT 4.400 425.320 2096.000 426.720 ;
        RECT 3.990 411.760 2096.000 425.320 ;
        RECT 3.990 410.360 2095.600 411.760 ;
        RECT 3.990 409.040 2096.000 410.360 ;
        RECT 4.400 407.640 2096.000 409.040 ;
        RECT 3.990 394.080 2096.000 407.640 ;
        RECT 3.990 392.680 2095.600 394.080 ;
        RECT 3.990 391.360 2096.000 392.680 ;
        RECT 4.400 389.960 2096.000 391.360 ;
        RECT 3.990 376.400 2096.000 389.960 ;
        RECT 3.990 375.000 2095.600 376.400 ;
        RECT 3.990 373.680 2096.000 375.000 ;
        RECT 4.400 372.280 2096.000 373.680 ;
        RECT 3.990 358.720 2096.000 372.280 ;
        RECT 3.990 357.320 2095.600 358.720 ;
        RECT 3.990 356.000 2096.000 357.320 ;
        RECT 4.400 354.600 2096.000 356.000 ;
        RECT 3.990 341.040 2096.000 354.600 ;
        RECT 3.990 339.680 2095.600 341.040 ;
        RECT 4.400 339.640 2095.600 339.680 ;
        RECT 4.400 338.280 2096.000 339.640 ;
        RECT 3.990 323.360 2096.000 338.280 ;
        RECT 3.990 322.000 2095.600 323.360 ;
        RECT 4.400 321.960 2095.600 322.000 ;
        RECT 4.400 320.600 2096.000 321.960 ;
        RECT 3.990 305.680 2096.000 320.600 ;
        RECT 3.990 304.320 2095.600 305.680 ;
        RECT 4.400 304.280 2095.600 304.320 ;
        RECT 4.400 302.920 2096.000 304.280 ;
        RECT 3.990 288.000 2096.000 302.920 ;
        RECT 3.990 286.640 2095.600 288.000 ;
        RECT 4.400 286.600 2095.600 286.640 ;
        RECT 4.400 285.240 2096.000 286.600 ;
        RECT 3.990 271.680 2096.000 285.240 ;
        RECT 3.990 270.280 2095.600 271.680 ;
        RECT 3.990 268.960 2096.000 270.280 ;
        RECT 4.400 267.560 2096.000 268.960 ;
        RECT 3.990 254.000 2096.000 267.560 ;
        RECT 3.990 252.600 2095.600 254.000 ;
        RECT 3.990 251.280 2096.000 252.600 ;
        RECT 4.400 249.880 2096.000 251.280 ;
        RECT 3.990 236.320 2096.000 249.880 ;
        RECT 3.990 234.920 2095.600 236.320 ;
        RECT 3.990 233.600 2096.000 234.920 ;
        RECT 4.400 232.200 2096.000 233.600 ;
        RECT 3.990 218.640 2096.000 232.200 ;
        RECT 3.990 217.240 2095.600 218.640 ;
        RECT 3.990 215.920 2096.000 217.240 ;
        RECT 4.400 214.520 2096.000 215.920 ;
        RECT 3.990 200.960 2096.000 214.520 ;
        RECT 3.990 199.560 2095.600 200.960 ;
        RECT 3.990 198.240 2096.000 199.560 ;
        RECT 4.400 196.840 2096.000 198.240 ;
        RECT 3.990 183.280 2096.000 196.840 ;
        RECT 3.990 181.880 2095.600 183.280 ;
        RECT 3.990 180.560 2096.000 181.880 ;
        RECT 4.400 179.160 2096.000 180.560 ;
        RECT 3.990 165.600 2096.000 179.160 ;
        RECT 3.990 164.200 2095.600 165.600 ;
        RECT 3.990 162.880 2096.000 164.200 ;
        RECT 4.400 161.480 2096.000 162.880 ;
        RECT 3.990 147.920 2096.000 161.480 ;
        RECT 3.990 146.520 2095.600 147.920 ;
        RECT 3.990 145.200 2096.000 146.520 ;
        RECT 4.400 143.800 2096.000 145.200 ;
        RECT 3.990 130.240 2096.000 143.800 ;
        RECT 3.990 128.840 2095.600 130.240 ;
        RECT 3.990 127.520 2096.000 128.840 ;
        RECT 4.400 126.120 2096.000 127.520 ;
        RECT 3.990 112.560 2096.000 126.120 ;
        RECT 3.990 111.160 2095.600 112.560 ;
        RECT 3.990 109.840 2096.000 111.160 ;
        RECT 4.400 108.440 2096.000 109.840 ;
        RECT 3.990 94.880 2096.000 108.440 ;
        RECT 3.990 93.480 2095.600 94.880 ;
        RECT 3.990 92.160 2096.000 93.480 ;
        RECT 4.400 90.760 2096.000 92.160 ;
        RECT 3.990 77.200 2096.000 90.760 ;
        RECT 3.990 75.800 2095.600 77.200 ;
        RECT 3.990 74.480 2096.000 75.800 ;
        RECT 4.400 73.080 2096.000 74.480 ;
        RECT 3.990 59.520 2096.000 73.080 ;
        RECT 3.990 58.120 2095.600 59.520 ;
        RECT 3.990 56.800 2096.000 58.120 ;
        RECT 4.400 55.400 2096.000 56.800 ;
        RECT 3.990 41.840 2096.000 55.400 ;
        RECT 3.990 40.440 2095.600 41.840 ;
        RECT 3.990 39.120 2096.000 40.440 ;
        RECT 4.400 37.720 2096.000 39.120 ;
        RECT 3.990 24.160 2096.000 37.720 ;
        RECT 3.990 22.760 2095.600 24.160 ;
        RECT 3.990 21.440 2096.000 22.760 ;
        RECT 4.400 20.040 2096.000 21.440 ;
        RECT 3.990 10.715 2096.000 20.040 ;
      LAYER met4 ;
        RECT 59.175 10.640 97.440 2287.760 ;
        RECT 99.840 10.640 2077.065 2287.760 ;
  END
END Ibtida_top_dffram_cv
END LIBRARY

